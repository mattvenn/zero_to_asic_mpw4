magic
tech sky130A
magscale 1 2
timestamp 1640163700
<< metal1 >>
rect 75822 703604 75828 703656
rect 75880 703644 75886 703656
rect 202598 703644 202604 703656
rect 75880 703616 202604 703644
rect 75880 703604 75886 703616
rect 202598 703604 202604 703616
rect 202656 703604 202662 703656
rect 86862 703536 86868 703588
rect 86920 703576 86926 703588
rect 234982 703576 234988 703588
rect 86920 703548 234988 703576
rect 86920 703536 86926 703548
rect 234982 703536 234988 703548
rect 235040 703536 235046 703588
rect 67634 703468 67640 703520
rect 67692 703508 67698 703520
rect 267458 703508 267464 703520
rect 67692 703480 267464 703508
rect 67692 703468 67698 703480
rect 267458 703468 267464 703480
rect 267516 703468 267522 703520
rect 93762 703400 93768 703452
rect 93820 703440 93826 703452
rect 300118 703440 300124 703452
rect 93820 703412 300124 703440
rect 93820 703400 93826 703412
rect 300118 703400 300124 703412
rect 300176 703400 300182 703452
rect 59262 703332 59268 703384
rect 59320 703372 59326 703384
rect 283834 703372 283840 703384
rect 59320 703344 283840 703372
rect 59320 703332 59326 703344
rect 283834 703332 283840 703344
rect 283892 703332 283898 703384
rect 73062 703264 73068 703316
rect 73120 703304 73126 703316
rect 332502 703304 332508 703316
rect 73120 703276 332508 703304
rect 73120 703264 73126 703276
rect 332502 703264 332508 703276
rect 332560 703264 332566 703316
rect 130378 703196 130384 703248
rect 130436 703236 130442 703248
rect 413646 703236 413652 703248
rect 130436 703208 413652 703236
rect 130436 703196 130442 703208
rect 413646 703196 413652 703208
rect 413704 703196 413710 703248
rect 62022 703128 62028 703180
rect 62080 703168 62086 703180
rect 348786 703168 348792 703180
rect 62080 703140 348792 703168
rect 62080 703128 62086 703140
rect 348786 703128 348792 703140
rect 348844 703128 348850 703180
rect 98730 703060 98736 703112
rect 98788 703100 98794 703112
rect 397454 703100 397460 703112
rect 98788 703072 397460 703100
rect 98788 703060 98794 703072
rect 397454 703060 397460 703072
rect 397512 703060 397518 703112
rect 124858 702992 124864 703044
rect 124916 703032 124922 703044
rect 429838 703032 429844 703044
rect 124916 703004 429844 703032
rect 124916 702992 124922 703004
rect 429838 702992 429844 703004
rect 429896 702992 429902 703044
rect 57882 702924 57888 702976
rect 57940 702964 57946 702976
rect 364978 702964 364984 702976
rect 57940 702936 364984 702964
rect 57940 702924 57946 702936
rect 364978 702924 364984 702936
rect 365036 702924 365042 702976
rect 126238 702856 126244 702908
rect 126296 702896 126302 702908
rect 462314 702896 462320 702908
rect 126296 702868 462320 702896
rect 126296 702856 126302 702868
rect 462314 702856 462320 702868
rect 462372 702856 462378 702908
rect 71038 702788 71044 702840
rect 71096 702828 71102 702840
rect 494790 702828 494796 702840
rect 71096 702800 494796 702828
rect 71096 702788 71102 702800
rect 494790 702788 494796 702800
rect 494848 702788 494854 702840
rect 97902 702720 97908 702772
rect 97960 702760 97966 702772
rect 478506 702760 478512 702772
rect 97960 702732 478512 702760
rect 97960 702720 97966 702732
rect 478506 702720 478512 702732
rect 478564 702720 478570 702772
rect 128998 702652 129004 702704
rect 129056 702692 129062 702704
rect 543458 702692 543464 702704
rect 129056 702664 543464 702692
rect 129056 702652 129062 702664
rect 543458 702652 543464 702664
rect 543516 702652 543522 702704
rect 8110 702584 8116 702636
rect 8168 702624 8174 702636
rect 89806 702624 89812 702636
rect 8168 702596 89812 702624
rect 8168 702584 8174 702596
rect 89806 702584 89812 702596
rect 89864 702584 89870 702636
rect 94498 702584 94504 702636
rect 94556 702624 94562 702636
rect 527174 702624 527180 702636
rect 94556 702596 527180 702624
rect 94556 702584 94562 702596
rect 527174 702584 527180 702596
rect 527232 702584 527238 702636
rect 55122 702516 55128 702568
rect 55180 702556 55186 702568
rect 580258 702556 580264 702568
rect 55180 702528 580264 702556
rect 55180 702516 55186 702528
rect 580258 702516 580264 702528
rect 580316 702516 580322 702568
rect 66162 702448 66168 702500
rect 66220 702488 66226 702500
rect 559650 702488 559656 702500
rect 66220 702460 559656 702488
rect 66220 702448 66226 702460
rect 559650 702448 559656 702460
rect 559708 702448 559714 702500
rect 83458 700272 83464 700324
rect 83516 700312 83522 700324
rect 89162 700312 89168 700324
rect 83516 700284 89168 700312
rect 83516 700272 83522 700284
rect 89162 700272 89168 700284
rect 89220 700272 89226 700324
rect 105446 700312 105452 700324
rect 93826 700284 105452 700312
rect 88978 700204 88984 700256
rect 89036 700244 89042 700256
rect 93826 700244 93854 700284
rect 105446 700272 105452 700284
rect 105504 700272 105510 700324
rect 133138 700272 133144 700324
rect 133196 700312 133202 700324
rect 218974 700312 218980 700324
rect 133196 700284 218980 700312
rect 133196 700272 133202 700284
rect 218974 700272 218980 700284
rect 219032 700272 219038 700324
rect 89036 700216 93854 700244
rect 89036 700204 89042 700216
rect 24302 698912 24308 698964
rect 24360 698952 24366 698964
rect 79318 698952 79324 698964
rect 24360 698924 79324 698952
rect 24360 698912 24366 698924
rect 79318 698912 79324 698924
rect 79376 698912 79382 698964
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 22738 670732 22744 670744
rect 3568 670704 22744 670732
rect 3568 670692 3574 670704
rect 22738 670692 22744 670704
rect 22796 670692 22802 670744
rect 2774 656956 2780 657008
rect 2832 656996 2838 657008
rect 4798 656996 4804 657008
rect 2832 656968 4804 656996
rect 2832 656956 2838 656968
rect 4798 656956 4804 656968
rect 4856 656956 4862 657008
rect 3510 632068 3516 632120
rect 3568 632108 3574 632120
rect 25498 632108 25504 632120
rect 3568 632080 25504 632108
rect 3568 632068 3574 632080
rect 25498 632068 25504 632080
rect 25556 632068 25562 632120
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 36538 618304 36544 618316
rect 3568 618276 36544 618304
rect 3568 618264 3574 618276
rect 36538 618264 36544 618276
rect 36596 618264 36602 618316
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 87598 605860 87604 605872
rect 3568 605832 87604 605860
rect 3568 605820 3574 605832
rect 87598 605820 87604 605832
rect 87656 605820 87662 605872
rect 79318 600244 79324 600296
rect 79376 600284 79382 600296
rect 79962 600284 79968 600296
rect 79376 600256 79968 600284
rect 79376 600244 79382 600256
rect 79962 600244 79968 600256
rect 80020 600244 80026 600296
rect 67450 599564 67456 599616
rect 67508 599604 67514 599616
rect 88978 599604 88984 599616
rect 67508 599576 88984 599604
rect 67508 599564 67514 599576
rect 88978 599564 88984 599576
rect 89036 599564 89042 599616
rect 79962 598952 79968 599004
rect 80020 598992 80026 599004
rect 114554 598992 114560 599004
rect 80020 598964 114560 598992
rect 80020 598952 80026 598964
rect 114554 598952 114560 598964
rect 114612 598952 114618 599004
rect 40034 598204 40040 598256
rect 40092 598244 40098 598256
rect 88886 598244 88892 598256
rect 40092 598216 88892 598244
rect 40092 598204 40098 598216
rect 88886 598204 88892 598216
rect 88944 598204 88950 598256
rect 67542 596776 67548 596828
rect 67600 596816 67606 596828
rect 169754 596816 169760 596828
rect 67600 596788 169760 596816
rect 67600 596776 67606 596788
rect 169754 596776 169760 596788
rect 169812 596776 169818 596828
rect 88978 595416 88984 595468
rect 89036 595456 89042 595468
rect 108298 595456 108304 595468
rect 89036 595428 108304 595456
rect 89036 595416 89042 595428
rect 108298 595416 108304 595428
rect 108356 595456 108362 595468
rect 582742 595456 582748 595468
rect 108356 595428 582748 595456
rect 108356 595416 108362 595428
rect 582742 595416 582748 595428
rect 582800 595416 582806 595468
rect 79778 594804 79784 594856
rect 79836 594844 79842 594856
rect 105538 594844 105544 594856
rect 79836 594816 105544 594844
rect 79836 594804 79842 594816
rect 105538 594804 105544 594816
rect 105596 594804 105602 594856
rect 87598 594396 87604 594448
rect 87656 594436 87662 594448
rect 91186 594436 91192 594448
rect 87656 594408 91192 594436
rect 87656 594396 87662 594408
rect 91186 594396 91192 594408
rect 91244 594396 91250 594448
rect 86218 593376 86224 593428
rect 86276 593416 86282 593428
rect 128538 593416 128544 593428
rect 86276 593388 128544 593416
rect 86276 593376 86282 593388
rect 128538 593376 128544 593388
rect 128596 593416 128602 593428
rect 582742 593416 582748 593428
rect 128596 593388 582748 593416
rect 128596 593376 128602 593388
rect 582742 593376 582748 593388
rect 582800 593376 582806 593428
rect 4798 592628 4804 592680
rect 4856 592668 4862 592680
rect 69014 592668 69020 592680
rect 4856 592640 69020 592668
rect 4856 592628 4862 592640
rect 69014 592628 69020 592640
rect 69072 592628 69078 592680
rect 75638 592084 75644 592136
rect 75696 592124 75702 592136
rect 96614 592124 96620 592136
rect 75696 592096 96620 592124
rect 75696 592084 75702 592096
rect 96614 592084 96620 592096
rect 96672 592084 96678 592136
rect 77938 592016 77944 592068
rect 77996 592056 78002 592068
rect 102134 592056 102140 592068
rect 77996 592028 102140 592056
rect 77996 592016 78002 592028
rect 102134 592016 102140 592028
rect 102192 592016 102198 592068
rect 70302 590724 70308 590776
rect 70360 590764 70366 590776
rect 75178 590764 75184 590776
rect 70360 590736 75184 590764
rect 70360 590724 70366 590736
rect 75178 590724 75184 590736
rect 75236 590724 75242 590776
rect 84102 590724 84108 590776
rect 84160 590764 84166 590776
rect 95878 590764 95884 590776
rect 84160 590736 95884 590764
rect 84160 590724 84166 590736
rect 95878 590724 95884 590736
rect 95936 590724 95942 590776
rect 78398 590656 78404 590708
rect 78456 590696 78462 590708
rect 100754 590696 100760 590708
rect 78456 590668 100760 590696
rect 78456 590656 78462 590668
rect 100754 590656 100760 590668
rect 100812 590656 100818 590708
rect 75178 589908 75184 589960
rect 75236 589948 75242 589960
rect 89714 589948 89720 589960
rect 75236 589920 89720 589948
rect 75236 589908 75242 589920
rect 89714 589908 89720 589920
rect 89772 589908 89778 589960
rect 72878 589364 72884 589416
rect 72936 589404 72942 589416
rect 93854 589404 93860 589416
rect 72936 589376 93860 589404
rect 72936 589364 72942 589376
rect 93854 589364 93860 589376
rect 93912 589364 93918 589416
rect 4798 589296 4804 589348
rect 4856 589336 4862 589348
rect 74856 589336 74862 589348
rect 4856 589308 74862 589336
rect 4856 589296 4862 589308
rect 74856 589296 74862 589308
rect 74914 589336 74920 589348
rect 75638 589336 75644 589348
rect 74914 589308 75644 589336
rect 74914 589296 74920 589308
rect 75638 589296 75644 589308
rect 75696 589296 75702 589348
rect 82630 589228 82636 589280
rect 82688 589268 82694 589280
rect 86954 589268 86960 589280
rect 82688 589240 86960 589268
rect 82688 589228 82694 589240
rect 86954 589228 86960 589240
rect 87012 589228 87018 589280
rect 69474 588616 69480 588668
rect 69532 588656 69538 588668
rect 69532 588628 80054 588656
rect 69532 588616 69538 588628
rect 80026 588520 80054 588628
rect 85298 588548 85304 588600
rect 85356 588588 85362 588600
rect 87046 588588 87052 588600
rect 85356 588560 87052 588588
rect 85356 588548 85362 588560
rect 87046 588548 87052 588560
rect 87104 588588 87110 588600
rect 113174 588588 113180 588600
rect 87104 588560 113180 588588
rect 87104 588548 87110 588560
rect 113174 588548 113180 588560
rect 113232 588548 113238 588600
rect 80026 588492 88932 588520
rect 83734 588412 83740 588464
rect 83792 588412 83798 588464
rect 52362 587868 52368 587920
rect 52420 587908 52426 587920
rect 66806 587908 66812 587920
rect 52420 587880 66812 587908
rect 52420 587868 52426 587880
rect 66806 587868 66812 587880
rect 66864 587868 66870 587920
rect 83752 587840 83780 588412
rect 88904 588328 88932 588492
rect 88886 588276 88892 588328
rect 88944 588276 88950 588328
rect 100754 588140 100760 588192
rect 100812 588180 100818 588192
rect 103514 588180 103520 588192
rect 100812 588152 103520 588180
rect 100812 588140 100818 588152
rect 103514 588140 103520 588152
rect 103572 588140 103578 588192
rect 92474 587840 92480 587852
rect 83752 587812 92480 587840
rect 92474 587800 92480 587812
rect 92532 587800 92538 587852
rect 59170 586508 59176 586560
rect 59228 586548 59234 586560
rect 66254 586548 66260 586560
rect 59228 586520 66260 586548
rect 59228 586508 59234 586520
rect 66254 586508 66260 586520
rect 66312 586508 66318 586560
rect 48222 585148 48228 585200
rect 48280 585188 48286 585200
rect 67726 585188 67732 585200
rect 48280 585160 67732 585188
rect 48280 585148 48286 585160
rect 67726 585148 67732 585160
rect 67784 585148 67790 585200
rect 91922 584400 91928 584452
rect 91980 584440 91986 584452
rect 93762 584440 93768 584452
rect 91980 584412 93768 584440
rect 91980 584400 91986 584412
rect 93762 584400 93768 584412
rect 93820 584440 93826 584452
rect 124214 584440 124220 584452
rect 93820 584412 124220 584440
rect 93820 584400 93826 584412
rect 124214 584400 124220 584412
rect 124272 584400 124278 584452
rect 91830 583652 91836 583704
rect 91888 583692 91894 583704
rect 93762 583692 93768 583704
rect 91888 583664 93768 583692
rect 91888 583652 91894 583664
rect 93762 583652 93768 583664
rect 93820 583692 93826 583704
rect 94498 583692 94504 583704
rect 93820 583664 94504 583692
rect 93820 583652 93826 583664
rect 94498 583652 94504 583664
rect 94556 583652 94562 583704
rect 50890 582360 50896 582412
rect 50948 582400 50954 582412
rect 66806 582400 66812 582412
rect 50948 582372 66812 582400
rect 50948 582360 50954 582372
rect 66806 582360 66812 582372
rect 66864 582360 66870 582412
rect 91094 581000 91100 581052
rect 91152 581040 91158 581052
rect 104158 581040 104164 581052
rect 91152 581012 104164 581040
rect 91152 581000 91158 581012
rect 104158 581000 104164 581012
rect 104216 581000 104222 581052
rect 2774 580456 2780 580508
rect 2832 580496 2838 580508
rect 4798 580496 4804 580508
rect 2832 580468 4804 580496
rect 2832 580456 2838 580468
rect 4798 580456 4804 580468
rect 4856 580456 4862 580508
rect 64782 579640 64788 579692
rect 64840 579680 64846 579692
rect 66806 579680 66812 579692
rect 64840 579652 66812 579680
rect 64840 579640 64846 579652
rect 66806 579640 66812 579652
rect 66864 579640 66870 579692
rect 91094 578212 91100 578264
rect 91152 578252 91158 578264
rect 121638 578252 121644 578264
rect 91152 578224 121644 578252
rect 91152 578212 91158 578224
rect 121638 578212 121644 578224
rect 121696 578212 121702 578264
rect 143442 577464 143448 577516
rect 143500 577504 143506 577516
rect 582466 577504 582472 577516
rect 143500 577476 582472 577504
rect 143500 577464 143506 577476
rect 582466 577464 582472 577476
rect 582524 577464 582530 577516
rect 91094 576852 91100 576904
rect 91152 576892 91158 576904
rect 142154 576892 142160 576904
rect 91152 576864 142160 576892
rect 91152 576852 91158 576864
rect 142154 576852 142160 576864
rect 142212 576892 142218 576904
rect 143442 576892 143448 576904
rect 142212 576864 143448 576892
rect 142212 576852 142218 576864
rect 143442 576852 143448 576864
rect 143500 576852 143506 576904
rect 25498 576104 25504 576156
rect 25556 576144 25562 576156
rect 47854 576144 47860 576156
rect 25556 576116 47860 576144
rect 25556 576104 25562 576116
rect 47854 576104 47860 576116
rect 47912 576104 47918 576156
rect 91186 576104 91192 576156
rect 91244 576144 91250 576156
rect 105630 576144 105636 576156
rect 91244 576116 105636 576144
rect 91244 576104 91250 576116
rect 105630 576104 105636 576116
rect 105688 576104 105694 576156
rect 47854 575492 47860 575544
rect 47912 575532 47918 575544
rect 48130 575532 48136 575544
rect 47912 575504 48136 575532
rect 47912 575492 47918 575504
rect 48130 575492 48136 575504
rect 48188 575532 48194 575544
rect 66898 575532 66904 575544
rect 48188 575504 66904 575532
rect 48188 575492 48194 575504
rect 66898 575492 66904 575504
rect 66956 575492 66962 575544
rect 55030 574744 55036 574796
rect 55088 574784 55094 574796
rect 67450 574784 67456 574796
rect 55088 574756 67456 574784
rect 55088 574744 55094 574756
rect 67450 574744 67456 574756
rect 67508 574744 67514 574796
rect 91094 574744 91100 574796
rect 91152 574784 91158 574796
rect 95142 574784 95148 574796
rect 91152 574756 95148 574784
rect 91152 574744 91158 574756
rect 95142 574744 95148 574756
rect 95200 574784 95206 574796
rect 98730 574784 98736 574796
rect 95200 574756 98736 574784
rect 95200 574744 95206 574756
rect 98730 574744 98736 574756
rect 98788 574744 98794 574796
rect 91094 572704 91100 572756
rect 91152 572744 91158 572756
rect 120626 572744 120632 572756
rect 91152 572716 120632 572744
rect 91152 572704 91158 572716
rect 120626 572704 120632 572716
rect 120684 572704 120690 572756
rect 91186 571412 91192 571464
rect 91244 571452 91250 571464
rect 108390 571452 108396 571464
rect 91244 571424 108396 571452
rect 91244 571412 91250 571424
rect 108390 571412 108396 571424
rect 108448 571412 108454 571464
rect 63310 571344 63316 571396
rect 63368 571384 63374 571396
rect 66438 571384 66444 571396
rect 63368 571356 66444 571384
rect 63368 571344 63374 571356
rect 66438 571344 66444 571356
rect 66496 571344 66502 571396
rect 91094 571344 91100 571396
rect 91152 571384 91158 571396
rect 129734 571384 129740 571396
rect 91152 571356 129740 571384
rect 91152 571344 91158 571356
rect 129734 571344 129740 571356
rect 129792 571344 129798 571396
rect 91094 569916 91100 569968
rect 91152 569956 91158 569968
rect 116578 569956 116584 569968
rect 91152 569928 116584 569956
rect 91152 569916 91158 569928
rect 116578 569916 116584 569928
rect 116636 569916 116642 569968
rect 60550 568556 60556 568608
rect 60608 568596 60614 568608
rect 66898 568596 66904 568608
rect 60608 568568 66904 568596
rect 60608 568556 60614 568568
rect 66898 568556 66904 568568
rect 66956 568556 66962 568608
rect 57790 567196 57796 567248
rect 57848 567236 57854 567248
rect 66898 567236 66904 567248
rect 57848 567208 66904 567236
rect 57848 567196 57854 567208
rect 66898 567196 66904 567208
rect 66956 567196 66962 567248
rect 88886 567196 88892 567248
rect 88944 567236 88950 567248
rect 133874 567236 133880 567248
rect 88944 567208 133880 567236
rect 88944 567196 88950 567208
rect 133874 567196 133880 567208
rect 133932 567196 133938 567248
rect 53742 566448 53748 566500
rect 53800 566488 53806 566500
rect 67542 566488 67548 566500
rect 53800 566460 67548 566488
rect 53800 566448 53806 566460
rect 67542 566448 67548 566460
rect 67600 566448 67606 566500
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 43438 565876 43444 565888
rect 3292 565848 43444 565876
rect 3292 565836 3298 565848
rect 43438 565836 43444 565848
rect 43496 565836 43502 565888
rect 91094 565836 91100 565888
rect 91152 565876 91158 565888
rect 126974 565876 126980 565888
rect 91152 565848 126980 565876
rect 91152 565836 91158 565848
rect 126974 565836 126980 565848
rect 127032 565836 127038 565888
rect 95878 565088 95884 565140
rect 95936 565128 95942 565140
rect 111794 565128 111800 565140
rect 95936 565100 111800 565128
rect 95936 565088 95942 565100
rect 111794 565088 111800 565100
rect 111852 565088 111858 565140
rect 51718 564340 51724 564392
rect 51776 564380 51782 564392
rect 55122 564380 55128 564392
rect 51776 564352 55128 564380
rect 51776 564340 51782 564352
rect 55122 564340 55128 564352
rect 55180 564380 55186 564392
rect 66806 564380 66812 564392
rect 55180 564352 66812 564380
rect 55180 564340 55186 564352
rect 66806 564340 66812 564352
rect 66864 564340 66870 564392
rect 91094 563048 91100 563100
rect 91152 563088 91158 563100
rect 133230 563088 133236 563100
rect 91152 563060 133236 563088
rect 91152 563048 91158 563060
rect 133230 563048 133236 563060
rect 133288 563048 133294 563100
rect 92198 562300 92204 562352
rect 92256 562340 92262 562352
rect 120718 562340 120724 562352
rect 92256 562312 120724 562340
rect 92256 562300 92262 562312
rect 120718 562300 120724 562312
rect 120776 562300 120782 562352
rect 35802 561688 35808 561740
rect 35860 561728 35866 561740
rect 66806 561728 66812 561740
rect 35860 561700 66812 561728
rect 35860 561688 35866 561700
rect 66806 561688 66812 561700
rect 66864 561688 66870 561740
rect 39942 560260 39948 560312
rect 40000 560300 40006 560312
rect 66530 560300 66536 560312
rect 40000 560272 66536 560300
rect 40000 560260 40006 560272
rect 66530 560260 66536 560272
rect 66588 560260 66594 560312
rect 56502 558900 56508 558952
rect 56560 558940 56566 558952
rect 66530 558940 66536 558952
rect 56560 558912 66536 558940
rect 56560 558900 56566 558912
rect 66530 558900 66536 558912
rect 66588 558900 66594 558952
rect 95142 558152 95148 558204
rect 95200 558192 95206 558204
rect 123202 558192 123208 558204
rect 95200 558164 123208 558192
rect 95200 558152 95206 558164
rect 123202 558152 123208 558164
rect 123260 558152 123266 558204
rect 50982 557540 50988 557592
rect 51040 557580 51046 557592
rect 67634 557580 67640 557592
rect 51040 557552 67640 557580
rect 51040 557540 51046 557552
rect 67634 557540 67640 557552
rect 67692 557540 67698 557592
rect 91186 557540 91192 557592
rect 91244 557580 91250 557592
rect 125594 557580 125600 557592
rect 91244 557552 125600 557580
rect 91244 557540 91250 557552
rect 125594 557540 125600 557552
rect 125652 557540 125658 557592
rect 91186 556180 91192 556232
rect 91244 556220 91250 556232
rect 121454 556220 121460 556232
rect 91244 556192 121460 556220
rect 91244 556180 91250 556192
rect 121454 556180 121460 556192
rect 121512 556180 121518 556232
rect 58894 554752 58900 554804
rect 58952 554792 58958 554804
rect 66622 554792 66628 554804
rect 58952 554764 66628 554792
rect 58952 554752 58958 554764
rect 66622 554752 66628 554764
rect 66680 554752 66686 554804
rect 91186 554752 91192 554804
rect 91244 554792 91250 554804
rect 100662 554792 100668 554804
rect 91244 554764 100668 554792
rect 91244 554752 91250 554764
rect 100662 554752 100668 554764
rect 100720 554792 100726 554804
rect 582466 554792 582472 554804
rect 100720 554764 582472 554792
rect 100720 554752 100726 554764
rect 582466 554752 582472 554764
rect 582524 554752 582530 554804
rect 3510 553800 3516 553852
rect 3568 553840 3574 553852
rect 7558 553840 7564 553852
rect 3568 553812 7564 553840
rect 3568 553800 3574 553812
rect 7558 553800 7564 553812
rect 7616 553800 7622 553852
rect 59262 553460 59268 553512
rect 59320 553500 59326 553512
rect 64138 553500 64144 553512
rect 59320 553472 64144 553500
rect 59320 553460 59326 553472
rect 64138 553460 64144 553472
rect 64196 553500 64202 553512
rect 66530 553500 66536 553512
rect 64196 553472 66536 553500
rect 64196 553460 64202 553472
rect 66530 553460 66536 553472
rect 66588 553460 66594 553512
rect 107010 553052 107016 553104
rect 107068 553092 107074 553104
rect 109034 553092 109040 553104
rect 107068 553064 109040 553092
rect 107068 553052 107074 553064
rect 109034 553052 109040 553064
rect 109092 553052 109098 553104
rect 91186 552304 91192 552356
rect 91244 552344 91250 552356
rect 95234 552344 95240 552356
rect 91244 552316 95240 552344
rect 91244 552304 91250 552316
rect 95234 552304 95240 552316
rect 95292 552304 95298 552356
rect 91186 552032 91192 552084
rect 91244 552072 91250 552084
rect 106918 552072 106924 552084
rect 91244 552044 106924 552072
rect 91244 552032 91250 552044
rect 106918 552032 106924 552044
rect 106976 552032 106982 552084
rect 60642 549244 60648 549296
rect 60700 549284 60706 549296
rect 66438 549284 66444 549296
rect 60700 549256 66444 549284
rect 60700 549244 60706 549256
rect 66438 549244 66444 549256
rect 66496 549244 66502 549296
rect 91186 549244 91192 549296
rect 91244 549284 91250 549296
rect 98730 549284 98736 549296
rect 91244 549256 98736 549284
rect 91244 549244 91250 549256
rect 98730 549244 98736 549256
rect 98788 549244 98794 549296
rect 91830 548496 91836 548548
rect 91888 548536 91894 548548
rect 121546 548536 121552 548548
rect 91888 548508 121552 548536
rect 91888 548496 91894 548508
rect 121546 548496 121552 548508
rect 121604 548496 121610 548548
rect 63402 547884 63408 547936
rect 63460 547924 63466 547936
rect 66530 547924 66536 547936
rect 63460 547896 66536 547924
rect 63460 547884 63466 547896
rect 66530 547884 66536 547896
rect 66588 547884 66594 547936
rect 62022 547748 62028 547800
rect 62080 547788 62086 547800
rect 66622 547788 66628 547800
rect 62080 547760 66628 547788
rect 62080 547748 62086 547760
rect 66622 547748 66628 547760
rect 66680 547748 66686 547800
rect 3418 547136 3424 547188
rect 3476 547176 3482 547188
rect 41230 547176 41236 547188
rect 3476 547148 41236 547176
rect 3476 547136 3482 547148
rect 41230 547136 41236 547148
rect 41288 547136 41294 547188
rect 41322 547136 41328 547188
rect 41380 547176 41386 547188
rect 62022 547176 62028 547188
rect 41380 547148 62028 547176
rect 41380 547136 41386 547148
rect 62022 547136 62028 547148
rect 62080 547136 62086 547188
rect 89990 546388 89996 546440
rect 90048 546428 90054 546440
rect 91002 546428 91008 546440
rect 90048 546400 91008 546428
rect 90048 546388 90054 546400
rect 91002 546388 91008 546400
rect 91060 546428 91066 546440
rect 126238 546428 126244 546440
rect 91060 546400 126244 546428
rect 91060 546388 91066 546400
rect 126238 546388 126244 546400
rect 126296 546388 126302 546440
rect 57514 545708 57520 545760
rect 57572 545748 57578 545760
rect 66162 545748 66168 545760
rect 57572 545720 66168 545748
rect 57572 545708 57578 545720
rect 66162 545708 66168 545720
rect 66220 545708 66226 545760
rect 91186 544348 91192 544400
rect 91244 544388 91250 544400
rect 95142 544388 95148 544400
rect 91244 544360 95148 544388
rect 91244 544348 91250 544360
rect 95142 544348 95148 544360
rect 95200 544388 95206 544400
rect 128998 544388 129004 544400
rect 95200 544360 129004 544388
rect 95200 544348 95206 544360
rect 128998 544348 129004 544360
rect 129056 544348 129062 544400
rect 57882 543736 57888 543788
rect 57940 543776 57946 543788
rect 62022 543776 62028 543788
rect 57940 543748 62028 543776
rect 57940 543736 57946 543748
rect 62022 543736 62028 543748
rect 62080 543776 62086 543788
rect 66806 543776 66812 543788
rect 62080 543748 66812 543776
rect 62080 543736 62086 543748
rect 66806 543736 66812 543748
rect 66864 543736 66870 543788
rect 41230 542376 41236 542428
rect 41288 542416 41294 542428
rect 44082 542416 44088 542428
rect 41288 542388 44088 542416
rect 41288 542376 41294 542388
rect 44082 542376 44088 542388
rect 44140 542416 44146 542428
rect 66806 542416 66812 542428
rect 44140 542388 66812 542416
rect 44140 542376 44146 542388
rect 66806 542376 66812 542388
rect 66864 542376 66870 542428
rect 91186 542376 91192 542428
rect 91244 542416 91250 542428
rect 104250 542416 104256 542428
rect 91244 542388 104256 542416
rect 91244 542376 91250 542388
rect 104250 542376 104256 542388
rect 104308 542376 104314 542428
rect 22738 541628 22744 541680
rect 22796 541668 22802 541680
rect 67082 541668 67088 541680
rect 22796 541640 67088 541668
rect 22796 541628 22802 541640
rect 67082 541628 67088 541640
rect 67140 541628 67146 541680
rect 91186 541628 91192 541680
rect 91244 541668 91250 541680
rect 136634 541668 136640 541680
rect 91244 541640 136640 541668
rect 91244 541628 91250 541640
rect 136634 541628 136640 541640
rect 136692 541628 136698 541680
rect 67542 540880 67548 540932
rect 67600 540920 67606 540932
rect 68646 540920 68652 540932
rect 67600 540892 68652 540920
rect 67600 540880 67606 540892
rect 68646 540880 68652 540892
rect 68704 540920 68710 540932
rect 582650 540920 582656 540932
rect 68704 540892 582656 540920
rect 68704 540880 68710 540892
rect 582650 540880 582656 540892
rect 582708 540880 582714 540932
rect 65978 539656 65984 539708
rect 66036 539696 66042 539708
rect 66036 539668 69888 539696
rect 66036 539656 66042 539668
rect 69860 539640 69888 539668
rect 91186 539656 91192 539708
rect 91244 539696 91250 539708
rect 93118 539696 93124 539708
rect 91244 539668 93124 539696
rect 91244 539656 91250 539668
rect 93118 539656 93124 539668
rect 93176 539656 93182 539708
rect 55122 539588 55128 539640
rect 55180 539628 55186 539640
rect 67542 539628 67548 539640
rect 55180 539600 67548 539628
rect 55180 539588 55186 539600
rect 67542 539588 67548 539600
rect 67600 539588 67606 539640
rect 69842 539588 69848 539640
rect 69900 539588 69906 539640
rect 89530 539520 89536 539572
rect 89588 539560 89594 539572
rect 89898 539560 89904 539572
rect 89588 539532 89904 539560
rect 89588 539520 89594 539532
rect 89898 539520 89904 539532
rect 89956 539520 89962 539572
rect 67082 539452 67088 539504
rect 67140 539492 67146 539504
rect 67542 539492 67548 539504
rect 67140 539464 67548 539492
rect 67140 539452 67146 539464
rect 67542 539452 67548 539464
rect 67600 539452 67606 539504
rect 67818 538908 67824 538960
rect 67876 538948 67882 538960
rect 74718 538948 74724 538960
rect 67876 538920 74724 538948
rect 67876 538908 67882 538920
rect 74718 538908 74724 538920
rect 74776 538908 74782 538960
rect 3418 538296 3424 538348
rect 3476 538336 3482 538348
rect 89530 538336 89536 538348
rect 3476 538308 89536 538336
rect 3476 538296 3482 538308
rect 89530 538296 89536 538308
rect 89588 538296 89594 538348
rect 80330 538228 80336 538280
rect 80388 538268 80394 538280
rect 80790 538268 80796 538280
rect 80388 538240 80796 538268
rect 80388 538228 80394 538240
rect 80790 538228 80796 538240
rect 80848 538268 80854 538280
rect 582558 538268 582564 538280
rect 80848 538240 582564 538268
rect 80848 538228 80854 538240
rect 582558 538228 582564 538240
rect 582616 538228 582622 538280
rect 7558 538160 7564 538212
rect 7616 538200 7622 538212
rect 70670 538200 70676 538212
rect 7616 538172 70676 538200
rect 7616 538160 7622 538172
rect 70670 538160 70676 538172
rect 70728 538160 70734 538212
rect 86862 538160 86868 538212
rect 86920 538200 86926 538212
rect 133138 538200 133144 538212
rect 86920 538172 133144 538200
rect 86920 538160 86926 538172
rect 133138 538160 133144 538172
rect 133196 538160 133202 538212
rect 72418 537480 72424 537532
rect 72476 537520 72482 537532
rect 579798 537520 579804 537532
rect 72476 537492 579804 537520
rect 72476 537480 72482 537492
rect 579798 537480 579804 537492
rect 579856 537480 579862 537532
rect 43438 536732 43444 536784
rect 43496 536772 43502 536784
rect 69658 536772 69664 536784
rect 43496 536744 69664 536772
rect 43496 536732 43502 536744
rect 69658 536732 69664 536744
rect 69716 536732 69722 536784
rect 82722 536732 82728 536784
rect 82780 536772 82786 536784
rect 130378 536772 130384 536784
rect 82780 536744 130384 536772
rect 82780 536732 82786 536744
rect 130378 536732 130384 536744
rect 130436 536732 130442 536784
rect 85482 536188 85488 536240
rect 85540 536228 85546 536240
rect 86218 536228 86224 536240
rect 85540 536200 86224 536228
rect 85540 536188 85546 536200
rect 86218 536188 86224 536200
rect 86276 536188 86282 536240
rect 36538 536052 36544 536104
rect 36596 536092 36602 536104
rect 49602 536092 49608 536104
rect 36596 536064 49608 536092
rect 36596 536052 36602 536064
rect 49602 536052 49608 536064
rect 49660 536092 49666 536104
rect 73154 536092 73160 536104
rect 49660 536064 73160 536092
rect 49660 536052 49666 536064
rect 73154 536052 73160 536064
rect 73212 536052 73218 536104
rect 73154 535440 73160 535492
rect 73212 535480 73218 535492
rect 73982 535480 73988 535492
rect 73212 535452 73988 535480
rect 73212 535440 73218 535452
rect 73982 535440 73988 535452
rect 74040 535440 74046 535492
rect 88610 535440 88616 535492
rect 88668 535480 88674 535492
rect 89622 535480 89628 535492
rect 88668 535452 89628 535480
rect 88668 535440 88674 535452
rect 89622 535440 89628 535452
rect 89680 535440 89686 535492
rect 8202 534692 8208 534744
rect 8260 534732 8266 534744
rect 91278 534732 91284 534744
rect 8260 534704 91284 534732
rect 8260 534692 8266 534704
rect 91278 534692 91284 534704
rect 91336 534692 91342 534744
rect 56502 534012 56508 534064
rect 56560 534052 56566 534064
rect 580258 534052 580264 534064
rect 56560 534024 580264 534052
rect 56560 534012 56566 534024
rect 580258 534012 580264 534024
rect 580316 534012 580322 534064
rect 67634 533400 67640 533452
rect 67692 533440 67698 533452
rect 68462 533440 68468 533452
rect 67692 533412 68468 533440
rect 67692 533400 67698 533412
rect 68462 533400 68468 533412
rect 68520 533400 68526 533452
rect 78674 533400 78680 533452
rect 78732 533440 78738 533452
rect 79502 533440 79508 533452
rect 78732 533412 79508 533440
rect 78732 533400 78738 533412
rect 79502 533400 79508 533412
rect 79560 533400 79566 533452
rect 4798 533332 4804 533384
rect 4856 533372 4862 533384
rect 91370 533372 91376 533384
rect 4856 533344 91376 533372
rect 4856 533332 4862 533344
rect 91370 533332 91376 533344
rect 91428 533332 91434 533384
rect 64782 531972 64788 532024
rect 64840 532012 64846 532024
rect 77938 532012 77944 532024
rect 64840 531984 77944 532012
rect 64840 531972 64846 531984
rect 77938 531972 77944 531984
rect 77996 531972 78002 532024
rect 23382 530544 23388 530596
rect 23440 530584 23446 530596
rect 91094 530584 91100 530596
rect 23440 530556 91100 530584
rect 23440 530544 23446 530556
rect 91094 530544 91100 530556
rect 91152 530544 91158 530596
rect 66162 529184 66168 529236
rect 66220 529224 66226 529236
rect 76466 529224 76472 529236
rect 66220 529196 76472 529224
rect 66220 529184 66226 529196
rect 76466 529184 76472 529196
rect 76524 529184 76530 529236
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 11698 514808 11704 514820
rect 3476 514780 11704 514808
rect 3476 514768 3482 514780
rect 11698 514768 11704 514780
rect 11756 514768 11762 514820
rect 39942 511232 39948 511284
rect 40000 511272 40006 511284
rect 580166 511272 580172 511284
rect 40000 511244 580172 511272
rect 40000 511232 40006 511244
rect 580166 511232 580172 511244
rect 580224 511232 580230 511284
rect 2774 501848 2780 501900
rect 2832 501888 2838 501900
rect 4798 501888 4804 501900
rect 2832 501860 4804 501888
rect 2832 501848 2838 501860
rect 4798 501848 4804 501860
rect 4856 501848 4862 501900
rect 67726 476008 67732 476060
rect 67784 476048 67790 476060
rect 76558 476048 76564 476060
rect 67784 476020 76564 476048
rect 67784 476008 67790 476020
rect 76558 476008 76564 476020
rect 76616 476008 76622 476060
rect 63310 475464 63316 475516
rect 63368 475504 63374 475516
rect 67818 475504 67824 475516
rect 63368 475476 67824 475504
rect 63368 475464 63374 475476
rect 67818 475464 67824 475476
rect 67876 475464 67882 475516
rect 3326 475328 3332 475380
rect 3384 475368 3390 475380
rect 8202 475368 8208 475380
rect 3384 475340 8208 475368
rect 3384 475328 3390 475340
rect 8202 475328 8208 475340
rect 8260 475368 8266 475380
rect 17218 475368 17224 475380
rect 8260 475340 17224 475368
rect 8260 475328 8266 475340
rect 17218 475328 17224 475340
rect 17276 475328 17282 475380
rect 57606 471248 57612 471300
rect 57664 471288 57670 471300
rect 78674 471288 78680 471300
rect 57664 471260 78680 471288
rect 57664 471248 57670 471260
rect 78674 471248 78680 471260
rect 78732 471248 78738 471300
rect 59078 468460 59084 468512
rect 59136 468500 59142 468512
rect 75914 468500 75920 468512
rect 59136 468472 75920 468500
rect 59136 468460 59142 468472
rect 75914 468460 75920 468472
rect 75972 468460 75978 468512
rect 89530 465740 89536 465792
rect 89588 465780 89594 465792
rect 125686 465780 125692 465792
rect 89588 465752 125692 465780
rect 89588 465740 89594 465752
rect 125686 465740 125692 465752
rect 125744 465740 125750 465792
rect 53650 465672 53656 465724
rect 53708 465712 53714 465724
rect 95878 465712 95884 465724
rect 53708 465684 95884 465712
rect 53708 465672 53714 465684
rect 95878 465672 95884 465684
rect 95936 465672 95942 465724
rect 66070 464312 66076 464364
rect 66128 464352 66134 464364
rect 78674 464352 78680 464364
rect 66128 464324 78680 464352
rect 66128 464312 66134 464324
rect 78674 464312 78680 464324
rect 78732 464312 78738 464364
rect 59170 462952 59176 463004
rect 59228 462992 59234 463004
rect 85574 462992 85580 463004
rect 59228 462964 85580 462992
rect 59228 462952 59234 462964
rect 85574 462952 85580 462964
rect 85632 462952 85638 463004
rect 2774 462544 2780 462596
rect 2832 462584 2838 462596
rect 4798 462584 4804 462596
rect 2832 462556 4804 462584
rect 2832 462544 2838 462556
rect 4798 462544 4804 462556
rect 4856 462544 4862 462596
rect 69014 462272 69020 462324
rect 69072 462312 69078 462324
rect 69842 462312 69848 462324
rect 69072 462284 69848 462312
rect 69072 462272 69078 462284
rect 69842 462272 69848 462284
rect 69900 462272 69906 462324
rect 52270 461592 52276 461644
rect 52328 461632 52334 461644
rect 73154 461632 73160 461644
rect 52328 461604 73160 461632
rect 52328 461592 52334 461604
rect 73154 461592 73160 461604
rect 73212 461592 73218 461644
rect 69014 460912 69020 460964
rect 69072 460952 69078 460964
rect 178034 460952 178040 460964
rect 69072 460924 178040 460952
rect 69072 460912 69078 460924
rect 178034 460912 178040 460924
rect 178092 460912 178098 460964
rect 48222 460164 48228 460216
rect 48280 460204 48286 460216
rect 82814 460204 82820 460216
rect 48280 460176 82820 460204
rect 48280 460164 48286 460176
rect 82814 460164 82820 460176
rect 82872 460164 82878 460216
rect 112438 458872 112444 458924
rect 112496 458912 112502 458924
rect 117314 458912 117320 458924
rect 112496 458884 117320 458912
rect 112496 458872 112502 458884
rect 117314 458872 117320 458884
rect 117372 458872 117378 458924
rect 106274 458804 106280 458856
rect 106332 458844 106338 458856
rect 114554 458844 114560 458856
rect 106332 458816 114560 458844
rect 106332 458804 106338 458816
rect 114554 458804 114560 458816
rect 114612 458844 114618 458856
rect 152458 458844 152464 458856
rect 114612 458816 152464 458844
rect 114612 458804 114618 458816
rect 152458 458804 152464 458816
rect 152516 458804 152522 458856
rect 52362 458192 52368 458244
rect 52420 458232 52426 458244
rect 53558 458232 53564 458244
rect 52420 458204 53564 458232
rect 52420 458192 52426 458204
rect 53558 458192 53564 458204
rect 53616 458232 53622 458244
rect 86954 458232 86960 458244
rect 53616 458204 86960 458232
rect 53616 458192 53622 458204
rect 86954 458192 86960 458204
rect 87012 458192 87018 458244
rect 63310 457444 63316 457496
rect 63368 457484 63374 457496
rect 80054 457484 80060 457496
rect 63368 457456 80060 457484
rect 63368 457444 63374 457456
rect 80054 457444 80060 457456
rect 80112 457444 80118 457496
rect 61838 456016 61844 456068
rect 61896 456056 61902 456068
rect 70486 456056 70492 456068
rect 61896 456028 70492 456056
rect 61896 456016 61902 456028
rect 70486 456016 70492 456028
rect 70544 456016 70550 456068
rect 77386 455336 77392 455388
rect 77444 455376 77450 455388
rect 77938 455376 77944 455388
rect 77444 455348 77944 455376
rect 77444 455336 77450 455348
rect 77938 455336 77944 455348
rect 77996 455336 78002 455388
rect 48130 454656 48136 454708
rect 48188 454696 48194 454708
rect 73154 454696 73160 454708
rect 48188 454668 73160 454696
rect 48188 454656 48194 454668
rect 73154 454656 73160 454668
rect 73212 454656 73218 454708
rect 77386 454112 77392 454164
rect 77444 454152 77450 454164
rect 128446 454152 128452 454164
rect 77444 454124 128452 454152
rect 77444 454112 77450 454124
rect 128446 454112 128452 454124
rect 128504 454112 128510 454164
rect 73154 454044 73160 454096
rect 73212 454084 73218 454096
rect 144178 454084 144184 454096
rect 73212 454056 144184 454084
rect 73212 454044 73218 454056
rect 144178 454044 144184 454056
rect 144236 454044 144242 454096
rect 22738 453976 22744 454028
rect 22796 454016 22802 454028
rect 23382 454016 23388 454028
rect 22796 453988 23388 454016
rect 22796 453976 22802 453988
rect 23382 453976 23388 453988
rect 23440 453976 23446 454028
rect 61746 453296 61752 453348
rect 61804 453336 61810 453348
rect 78766 453336 78772 453348
rect 61804 453308 78772 453336
rect 61804 453296 61810 453308
rect 78766 453296 78772 453308
rect 78824 453296 78830 453348
rect 82814 452684 82820 452736
rect 82872 452724 82878 452736
rect 83458 452724 83464 452736
rect 82872 452696 83464 452724
rect 82872 452684 82878 452696
rect 83458 452684 83464 452696
rect 83516 452724 83522 452736
rect 161474 452724 161480 452736
rect 83516 452696 161480 452724
rect 83516 452684 83522 452696
rect 161474 452684 161480 452696
rect 161532 452684 161538 452736
rect 22738 452616 22744 452668
rect 22796 452656 22802 452668
rect 124950 452656 124956 452668
rect 22796 452628 124956 452656
rect 22796 452616 22802 452628
rect 124950 452616 124956 452628
rect 125008 452616 125014 452668
rect 61930 451868 61936 451920
rect 61988 451908 61994 451920
rect 91554 451908 91560 451920
rect 61988 451880 91560 451908
rect 61988 451868 61994 451880
rect 91554 451868 91560 451880
rect 91612 451868 91618 451920
rect 50798 451256 50804 451308
rect 50856 451296 50862 451308
rect 74718 451296 74724 451308
rect 50856 451268 74724 451296
rect 50856 451256 50862 451268
rect 74718 451256 74724 451268
rect 74776 451256 74782 451308
rect 98638 451256 98644 451308
rect 98696 451296 98702 451308
rect 179414 451296 179420 451308
rect 98696 451268 179420 451296
rect 98696 451256 98702 451268
rect 179414 451256 179420 451268
rect 179472 451256 179478 451308
rect 4798 451188 4804 451240
rect 4856 451228 4862 451240
rect 103514 451228 103520 451240
rect 4856 451200 103520 451228
rect 4856 451188 4862 451200
rect 103514 451188 103520 451200
rect 103572 451228 103578 451240
rect 104618 451228 104624 451240
rect 103572 451200 104624 451228
rect 103572 451188 103578 451200
rect 104618 451188 104624 451200
rect 104676 451188 104682 451240
rect 173802 451188 173808 451240
rect 173860 451228 173866 451240
rect 582466 451228 582472 451240
rect 173860 451200 582472 451228
rect 173860 451188 173866 451200
rect 582466 451188 582472 451200
rect 582524 451188 582530 451240
rect 55030 450508 55036 450560
rect 55088 450548 55094 450560
rect 71774 450548 71780 450560
rect 55088 450520 71780 450548
rect 55088 450508 55094 450520
rect 71774 450508 71780 450520
rect 71832 450508 71838 450560
rect 104066 449964 104072 450016
rect 104124 450004 104130 450016
rect 104618 450004 104624 450016
rect 104124 449976 104624 450004
rect 104124 449964 104130 449976
rect 104618 449964 104624 449976
rect 104676 450004 104682 450016
rect 166994 450004 167000 450016
rect 104676 449976 167000 450004
rect 104676 449964 104682 449976
rect 166994 449964 167000 449976
rect 167052 449964 167058 450016
rect 172514 449936 172520 449948
rect 81084 449908 172520 449936
rect 50890 449828 50896 449880
rect 50948 449868 50954 449880
rect 80882 449868 80888 449880
rect 50948 449840 80888 449868
rect 50948 449828 50954 449840
rect 80882 449828 80888 449840
rect 80940 449868 80946 449880
rect 81084 449868 81112 449908
rect 172514 449896 172520 449908
rect 172572 449936 172578 449948
rect 173802 449936 173808 449948
rect 172572 449908 173808 449936
rect 172572 449896 172578 449908
rect 173802 449896 173808 449908
rect 173860 449896 173866 449948
rect 80940 449840 81112 449868
rect 80940 449828 80946 449840
rect 64690 449148 64696 449200
rect 64748 449188 64754 449200
rect 74626 449188 74632 449200
rect 64748 449160 74632 449188
rect 64748 449148 64754 449160
rect 74626 449148 74632 449160
rect 74684 449148 74690 449200
rect 116578 449148 116584 449200
rect 116636 449188 116642 449200
rect 128354 449188 128360 449200
rect 116636 449160 128360 449188
rect 116636 449148 116642 449160
rect 128354 449148 128360 449160
rect 128412 449148 128418 449200
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 40678 448576 40684 448588
rect 3200 448548 40684 448576
rect 3200 448536 3206 448548
rect 40678 448536 40684 448548
rect 40736 448536 40742 448588
rect 108298 448536 108304 448588
rect 108356 448576 108362 448588
rect 130378 448576 130384 448588
rect 108356 448548 130384 448576
rect 108356 448536 108362 448548
rect 130378 448536 130384 448548
rect 130436 448536 130442 448588
rect 11698 448468 11704 448520
rect 11756 448508 11762 448520
rect 111794 448508 111800 448520
rect 11756 448480 111800 448508
rect 11756 448468 11762 448480
rect 111794 448468 111800 448480
rect 111852 448468 111858 448520
rect 105630 447788 105636 447840
rect 105688 447828 105694 447840
rect 122926 447828 122932 447840
rect 105688 447800 122932 447828
rect 105688 447788 105694 447800
rect 122926 447788 122932 447800
rect 122984 447788 122990 447840
rect 68370 447108 68376 447160
rect 68428 447148 68434 447160
rect 88794 447148 88800 447160
rect 68428 447120 88800 447148
rect 68428 447108 68434 447120
rect 88794 447108 88800 447120
rect 88852 447108 88858 447160
rect 60458 446360 60464 446412
rect 60516 446400 60522 446412
rect 77294 446400 77300 446412
rect 60516 446372 77300 446400
rect 60516 446360 60522 446372
rect 77294 446360 77300 446372
rect 77352 446360 77358 446412
rect 111794 445816 111800 445868
rect 111852 445856 111858 445868
rect 112990 445856 112996 445868
rect 111852 445828 112996 445856
rect 111852 445816 111858 445828
rect 112990 445816 112996 445828
rect 113048 445856 113054 445868
rect 142798 445856 142804 445868
rect 113048 445828 142804 445856
rect 113048 445816 113054 445828
rect 142798 445816 142804 445828
rect 142856 445816 142862 445868
rect 76558 445748 76564 445800
rect 76616 445788 76622 445800
rect 124858 445788 124864 445800
rect 76616 445760 124864 445788
rect 76616 445748 76622 445760
rect 124858 445748 124864 445760
rect 124916 445748 124922 445800
rect 59170 444456 59176 444508
rect 59228 444496 59234 444508
rect 92474 444496 92480 444508
rect 59228 444468 92480 444496
rect 59228 444456 59234 444468
rect 92474 444456 92480 444468
rect 92532 444496 92538 444508
rect 93072 444496 93078 444508
rect 92532 444468 93078 444496
rect 92532 444456 92538 444468
rect 93072 444456 93078 444468
rect 93130 444456 93136 444508
rect 101398 444456 101404 444508
rect 101456 444496 101462 444508
rect 126238 444496 126244 444508
rect 101456 444468 126244 444496
rect 101456 444456 101462 444468
rect 126238 444456 126244 444468
rect 126296 444456 126302 444508
rect 4798 444388 4804 444440
rect 4856 444428 4862 444440
rect 118694 444428 118700 444440
rect 4856 444400 118700 444428
rect 4856 444388 4862 444400
rect 118694 444388 118700 444400
rect 118752 444388 118758 444440
rect 67358 442892 67364 442944
rect 67416 442932 67422 442944
rect 67726 442932 67732 442944
rect 67416 442904 67732 442932
rect 67416 442892 67422 442904
rect 67726 442892 67732 442904
rect 67784 442892 67790 442944
rect 60366 442212 60372 442264
rect 60424 442252 60430 442264
rect 68370 442252 68376 442264
rect 60424 442224 68376 442252
rect 60424 442212 60430 442224
rect 68370 442212 68376 442224
rect 68428 442212 68434 442264
rect 124122 439492 124128 439544
rect 124180 439532 124186 439544
rect 125686 439532 125692 439544
rect 124180 439504 125692 439532
rect 124180 439492 124186 439504
rect 125686 439492 125692 439504
rect 125744 439532 125750 439544
rect 157334 439532 157340 439544
rect 125744 439504 157340 439532
rect 125744 439492 125750 439504
rect 157334 439492 157340 439504
rect 157392 439492 157398 439544
rect 60550 439016 60556 439068
rect 60608 439056 60614 439068
rect 66990 439056 66996 439068
rect 60608 439028 66996 439056
rect 60608 439016 60614 439028
rect 66990 439016 66996 439028
rect 67048 439056 67054 439068
rect 67358 439056 67364 439068
rect 67048 439028 67364 439056
rect 67048 439016 67054 439028
rect 67358 439016 67364 439028
rect 67416 439016 67422 439068
rect 57790 438132 57796 438184
rect 57848 438172 57854 438184
rect 66070 438172 66076 438184
rect 57848 438144 66076 438172
rect 57848 438132 57854 438144
rect 66070 438132 66076 438144
rect 66128 438172 66134 438184
rect 66530 438172 66536 438184
rect 66128 438144 66536 438172
rect 66128 438132 66134 438144
rect 66530 438132 66536 438144
rect 66588 438132 66594 438184
rect 123662 438132 123668 438184
rect 123720 438172 123726 438184
rect 124214 438172 124220 438184
rect 123720 438144 124220 438172
rect 123720 438132 123726 438144
rect 124214 438132 124220 438144
rect 124272 438172 124278 438184
rect 157978 438172 157984 438184
rect 124272 438144 157984 438172
rect 124272 438132 124278 438144
rect 157978 438132 157984 438144
rect 158036 438132 158042 438184
rect 52454 436024 52460 436076
rect 52512 436064 52518 436076
rect 53742 436064 53748 436076
rect 52512 436036 53748 436064
rect 52512 436024 52518 436036
rect 53742 436024 53748 436036
rect 53800 436064 53806 436076
rect 66806 436064 66812 436076
rect 53800 436036 66812 436064
rect 53800 436024 53806 436036
rect 66806 436024 66812 436036
rect 66864 436024 66870 436076
rect 39850 435344 39856 435396
rect 39908 435384 39914 435396
rect 52454 435384 52460 435396
rect 39908 435356 52460 435384
rect 39908 435344 39914 435356
rect 52454 435344 52460 435356
rect 52512 435344 52518 435396
rect 52178 433304 52184 433356
rect 52236 433344 52242 433356
rect 65518 433344 65524 433356
rect 52236 433316 65524 433344
rect 52236 433304 52242 433316
rect 65518 433304 65524 433316
rect 65576 433304 65582 433356
rect 65536 433276 65564 433304
rect 66438 433276 66444 433288
rect 65536 433248 66444 433276
rect 66438 433236 66444 433248
rect 66496 433236 66502 433288
rect 123846 432556 123852 432608
rect 123904 432596 123910 432608
rect 171134 432596 171140 432608
rect 123904 432568 171140 432596
rect 123904 432556 123910 432568
rect 171134 432556 171140 432568
rect 171192 432596 171198 432608
rect 582374 432596 582380 432608
rect 171192 432568 582380 432596
rect 171192 432556 171198 432568
rect 582374 432556 582380 432568
rect 582432 432556 582438 432608
rect 48130 431944 48136 431996
rect 48188 431984 48194 431996
rect 48188 431956 51764 431984
rect 48188 431944 48194 431956
rect 51736 431928 51764 431956
rect 51718 431916 51724 431928
rect 51631 431888 51724 431916
rect 51718 431876 51724 431888
rect 51776 431916 51782 431928
rect 66806 431916 66812 431928
rect 51776 431888 66812 431916
rect 51776 431876 51782 431888
rect 66806 431876 66812 431888
rect 66864 431876 66870 431928
rect 34514 429088 34520 429140
rect 34572 429128 34578 429140
rect 35802 429128 35808 429140
rect 34572 429100 35808 429128
rect 34572 429088 34578 429100
rect 35802 429088 35808 429100
rect 35860 429128 35866 429140
rect 66806 429128 66812 429140
rect 35860 429100 66812 429128
rect 35860 429088 35866 429100
rect 66806 429088 66812 429100
rect 66864 429088 66870 429140
rect 15838 428408 15844 428460
rect 15896 428448 15902 428460
rect 34514 428448 34520 428460
rect 15896 428420 34520 428448
rect 15896 428408 15902 428420
rect 34514 428408 34520 428420
rect 34572 428408 34578 428460
rect 39942 425688 39948 425740
rect 40000 425728 40006 425740
rect 58986 425728 58992 425740
rect 40000 425700 58992 425728
rect 40000 425688 40006 425700
rect 58986 425688 58992 425700
rect 59044 425688 59050 425740
rect 58986 425076 58992 425128
rect 59044 425116 59050 425128
rect 66806 425116 66812 425128
rect 59044 425088 66812 425116
rect 59044 425076 59050 425088
rect 66806 425076 66812 425088
rect 66864 425076 66870 425128
rect 56502 424328 56508 424380
rect 56560 424368 56566 424380
rect 63218 424368 63224 424380
rect 56560 424340 63224 424368
rect 56560 424328 56566 424340
rect 63218 424328 63224 424340
rect 63276 424368 63282 424380
rect 66806 424368 66812 424380
rect 63276 424340 66812 424368
rect 63276 424328 63282 424340
rect 66806 424328 66812 424340
rect 66864 424328 66870 424380
rect 3418 423580 3424 423632
rect 3476 423620 3482 423632
rect 22738 423620 22744 423632
rect 3476 423592 22744 423620
rect 3476 423580 3482 423592
rect 22738 423580 22744 423592
rect 22796 423580 22802 423632
rect 50982 421540 50988 421592
rect 51040 421580 51046 421592
rect 64782 421580 64788 421592
rect 51040 421552 64788 421580
rect 51040 421540 51046 421552
rect 64782 421540 64788 421552
rect 64840 421580 64846 421592
rect 66806 421580 66812 421592
rect 64840 421552 66812 421580
rect 64840 421540 64846 421552
rect 66806 421540 66812 421552
rect 66864 421540 66870 421592
rect 123202 421540 123208 421592
rect 123260 421580 123266 421592
rect 134518 421580 134524 421592
rect 123260 421552 134524 421580
rect 123260 421540 123266 421552
rect 134518 421540 134524 421552
rect 134576 421540 134582 421592
rect 56502 419500 56508 419552
rect 56560 419540 56566 419552
rect 66898 419540 66904 419552
rect 56560 419512 66904 419540
rect 56560 419500 56566 419512
rect 66898 419500 66904 419512
rect 66956 419500 66962 419552
rect 58894 418072 58900 418124
rect 58952 418112 58958 418124
rect 65518 418112 65524 418124
rect 58952 418084 65524 418112
rect 58952 418072 58958 418084
rect 65518 418072 65524 418084
rect 65576 418112 65582 418124
rect 66438 418112 66444 418124
rect 65576 418084 66444 418112
rect 65576 418072 65582 418084
rect 66438 418072 66444 418084
rect 66496 418072 66502 418124
rect 124122 415148 124128 415200
rect 124180 415188 124186 415200
rect 129734 415188 129740 415200
rect 124180 415160 129740 415188
rect 124180 415148 124186 415160
rect 129734 415148 129740 415160
rect 129792 415148 129798 415200
rect 57790 414672 57796 414724
rect 57848 414712 57854 414724
rect 64138 414712 64144 414724
rect 57848 414684 64144 414712
rect 57848 414672 57854 414684
rect 64138 414672 64144 414684
rect 64196 414712 64202 414724
rect 66806 414712 66812 414724
rect 64196 414684 66812 414712
rect 64196 414672 64202 414684
rect 66806 414672 66812 414684
rect 66864 414672 66870 414724
rect 129734 414672 129740 414724
rect 129792 414712 129798 414724
rect 131114 414712 131120 414724
rect 129792 414684 131120 414712
rect 129792 414672 129798 414684
rect 131114 414672 131120 414684
rect 131172 414672 131178 414724
rect 123018 412564 123024 412616
rect 123076 412604 123082 412616
rect 128354 412604 128360 412616
rect 123076 412576 128360 412604
rect 123076 412564 123082 412576
rect 128354 412564 128360 412576
rect 128412 412564 128418 412616
rect 123018 411272 123024 411324
rect 123076 411312 123082 411324
rect 123478 411312 123484 411324
rect 123076 411284 123484 411312
rect 123076 411272 123082 411284
rect 123478 411272 123484 411284
rect 123536 411272 123542 411324
rect 121178 409844 121184 409896
rect 121236 409884 121242 409896
rect 135898 409884 135904 409896
rect 121236 409856 135904 409884
rect 121236 409844 121242 409856
rect 135898 409844 135904 409856
rect 135956 409844 135962 409896
rect 60642 408416 60648 408468
rect 60700 408456 60706 408468
rect 68370 408456 68376 408468
rect 60700 408428 68376 408456
rect 60700 408416 60706 408428
rect 68370 408416 68376 408428
rect 68428 408416 68434 408468
rect 124122 407736 124128 407788
rect 124180 407776 124186 407788
rect 133874 407776 133880 407788
rect 124180 407748 133880 407776
rect 124180 407736 124186 407748
rect 133874 407736 133880 407748
rect 133932 407776 133938 407788
rect 134610 407776 134616 407788
rect 133932 407748 134616 407776
rect 133932 407736 133938 407748
rect 134610 407736 134616 407748
rect 134668 407736 134674 407788
rect 63402 406580 63408 406632
rect 63460 406620 63466 406632
rect 64598 406620 64604 406632
rect 63460 406592 64604 406620
rect 63460 406580 63466 406592
rect 64598 406580 64604 406592
rect 64656 406580 64662 406632
rect 64598 406104 64604 406156
rect 64656 406144 64662 406156
rect 66254 406144 66260 406156
rect 64656 406116 66260 406144
rect 64656 406104 64662 406116
rect 66254 406104 66260 406116
rect 66312 406104 66318 406156
rect 124122 406104 124128 406156
rect 124180 406144 124186 406156
rect 126882 406144 126888 406156
rect 124180 406116 126888 406144
rect 124180 406104 124186 406116
rect 126882 406104 126888 406116
rect 126940 406104 126946 406156
rect 41322 404948 41328 405000
rect 41380 404988 41386 405000
rect 57698 404988 57704 405000
rect 41380 404960 57704 404988
rect 41380 404948 41386 404960
rect 57698 404948 57704 404960
rect 57756 404948 57762 405000
rect 57698 403588 57704 403640
rect 57756 403628 57762 403640
rect 66254 403628 66260 403640
rect 57756 403600 66260 403628
rect 57756 403588 57762 403600
rect 66254 403588 66260 403600
rect 66312 403588 66318 403640
rect 163498 403588 163504 403640
rect 163556 403628 163562 403640
rect 582374 403628 582380 403640
rect 163556 403600 582380 403628
rect 163556 403588 163562 403600
rect 582374 403588 582380 403600
rect 582432 403588 582438 403640
rect 124030 402976 124036 403028
rect 124088 403016 124094 403028
rect 163498 403016 163504 403028
rect 124088 402988 163504 403016
rect 124088 402976 124094 402988
rect 163498 402976 163504 402988
rect 163556 402976 163562 403028
rect 50890 401548 50896 401600
rect 50948 401588 50954 401600
rect 57514 401588 57520 401600
rect 50948 401560 57520 401588
rect 50948 401548 50954 401560
rect 57514 401548 57520 401560
rect 57572 401588 57578 401600
rect 66254 401588 66260 401600
rect 57572 401560 66260 401588
rect 57572 401548 57578 401560
rect 66254 401548 66260 401560
rect 66312 401548 66318 401600
rect 124122 401548 124128 401600
rect 124180 401588 124186 401600
rect 133230 401588 133236 401600
rect 124180 401560 133236 401588
rect 124180 401548 124186 401560
rect 133230 401548 133236 401560
rect 133288 401588 133294 401600
rect 133782 401588 133788 401600
rect 133288 401560 133788 401588
rect 133288 401548 133294 401560
rect 133782 401548 133788 401560
rect 133840 401548 133846 401600
rect 124950 400188 124956 400240
rect 125008 400228 125014 400240
rect 169754 400228 169760 400240
rect 125008 400200 169760 400228
rect 125008 400188 125014 400200
rect 169754 400188 169760 400200
rect 169812 400188 169818 400240
rect 123662 400120 123668 400172
rect 123720 400160 123726 400172
rect 124968 400160 124996 400188
rect 123720 400132 124996 400160
rect 123720 400120 123726 400132
rect 2774 398692 2780 398744
rect 2832 398732 2838 398744
rect 4798 398732 4804 398744
rect 2832 398704 4804 398732
rect 2832 398692 2838 398704
rect 4798 398692 4804 398704
rect 4856 398692 4862 398744
rect 43990 398080 43996 398132
rect 44048 398120 44054 398132
rect 62022 398120 62028 398132
rect 44048 398092 62028 398120
rect 44048 398080 44054 398092
rect 62022 398080 62028 398092
rect 62080 398120 62086 398132
rect 66438 398120 66444 398132
rect 62080 398092 66444 398120
rect 62080 398080 62086 398092
rect 66438 398080 66444 398092
rect 66496 398080 66502 398132
rect 44082 396720 44088 396772
rect 44140 396760 44146 396772
rect 66990 396760 66996 396772
rect 44140 396732 66996 396760
rect 44140 396720 44146 396732
rect 66990 396720 66996 396732
rect 67048 396760 67054 396772
rect 67266 396760 67272 396772
rect 67048 396732 67272 396760
rect 67048 396720 67054 396732
rect 67266 396720 67272 396732
rect 67324 396720 67330 396772
rect 121546 396040 121552 396092
rect 121604 396080 121610 396092
rect 171226 396080 171232 396092
rect 121604 396052 171232 396080
rect 121604 396040 121610 396052
rect 171226 396040 171232 396052
rect 171284 396040 171290 396092
rect 123662 395972 123668 396024
rect 123720 396012 123726 396024
rect 125594 396012 125600 396024
rect 123720 395984 125600 396012
rect 123720 395972 123726 395984
rect 125594 395972 125600 395984
rect 125652 395972 125658 396024
rect 55122 393252 55128 393304
rect 55180 393292 55186 393304
rect 61930 393292 61936 393304
rect 55180 393264 61936 393292
rect 55180 393252 55186 393264
rect 61930 393252 61936 393264
rect 61988 393292 61994 393304
rect 66806 393292 66812 393304
rect 61988 393264 66812 393292
rect 61988 393252 61994 393264
rect 66806 393252 66812 393264
rect 66864 393252 66870 393304
rect 59078 391212 59084 391264
rect 59136 391252 59142 391264
rect 59136 391224 64874 391252
rect 59136 391212 59142 391224
rect 64846 390980 64874 391224
rect 81434 390980 81440 390992
rect 64846 390952 81440 390980
rect 81434 390940 81440 390952
rect 81492 390980 81498 390992
rect 82078 390980 82084 390992
rect 81492 390952 82084 390980
rect 81492 390940 81498 390952
rect 82078 390940 82084 390952
rect 82136 390940 82142 390992
rect 115842 390532 115848 390584
rect 115900 390572 115906 390584
rect 120810 390572 120816 390584
rect 115900 390544 120816 390572
rect 115900 390532 115906 390544
rect 120810 390532 120816 390544
rect 120868 390532 120874 390584
rect 3418 389784 3424 389836
rect 3476 389824 3482 389836
rect 85482 389824 85488 389836
rect 3476 389796 85488 389824
rect 3476 389784 3482 389796
rect 85482 389784 85488 389796
rect 85540 389784 85546 389836
rect 57606 389172 57612 389224
rect 57664 389212 57670 389224
rect 86954 389212 86960 389224
rect 57664 389184 86960 389212
rect 57664 389172 57670 389184
rect 86954 389172 86960 389184
rect 87012 389172 87018 389224
rect 117774 389172 117780 389224
rect 117832 389212 117838 389224
rect 165614 389212 165620 389224
rect 117832 389184 165620 389212
rect 117832 389172 117838 389184
rect 165614 389172 165620 389184
rect 165672 389172 165678 389224
rect 49602 389104 49608 389156
rect 49660 389144 49666 389156
rect 76650 389144 76656 389156
rect 49660 389116 76656 389144
rect 49660 389104 49666 389116
rect 76650 389104 76656 389116
rect 76708 389104 76714 389156
rect 104066 389104 104072 389156
rect 104124 389144 104130 389156
rect 136634 389144 136640 389156
rect 104124 389116 136640 389144
rect 104124 389104 104130 389116
rect 136634 389104 136640 389116
rect 136692 389104 136698 389156
rect 61838 389036 61844 389088
rect 61896 389076 61902 389088
rect 61896 389048 64874 389076
rect 61896 389036 61902 389048
rect 64846 389008 64874 389048
rect 67634 389036 67640 389088
rect 67692 389076 67698 389088
rect 68462 389076 68468 389088
rect 67692 389048 68468 389076
rect 67692 389036 67698 389048
rect 68462 389036 68468 389048
rect 68520 389036 68526 389088
rect 119430 389036 119436 389088
rect 119488 389076 119494 389088
rect 120166 389076 120172 389088
rect 119488 389048 120172 389076
rect 119488 389036 119494 389048
rect 120166 389036 120172 389048
rect 120224 389036 120230 389088
rect 73154 389008 73160 389020
rect 64846 388980 73160 389008
rect 73154 388968 73160 388980
rect 73212 389008 73218 389020
rect 73338 389008 73344 389020
rect 73212 388980 73344 389008
rect 73212 388968 73218 388980
rect 73338 388968 73344 388980
rect 73396 388968 73402 389020
rect 93394 388424 93400 388476
rect 93452 388464 93458 388476
rect 112438 388464 112444 388476
rect 93452 388436 112444 388464
rect 93452 388424 93458 388436
rect 112438 388424 112444 388436
rect 112496 388424 112502 388476
rect 93670 388016 93676 388068
rect 93728 388056 93734 388068
rect 94222 388056 94228 388068
rect 93728 388028 94228 388056
rect 93728 388016 93734 388028
rect 94222 388016 94228 388028
rect 94280 388016 94286 388068
rect 79962 387812 79968 387864
rect 80020 387852 80026 387864
rect 80606 387852 80612 387864
rect 80020 387824 80612 387852
rect 80020 387812 80026 387824
rect 80606 387812 80612 387824
rect 80664 387812 80670 387864
rect 64690 387744 64696 387796
rect 64748 387784 64754 387796
rect 79318 387784 79324 387796
rect 64748 387756 79324 387784
rect 64748 387744 64754 387756
rect 79318 387744 79324 387756
rect 79376 387744 79382 387796
rect 111702 387064 111708 387116
rect 111760 387104 111766 387116
rect 120626 387104 120632 387116
rect 111760 387076 120632 387104
rect 111760 387064 111766 387076
rect 120626 387064 120632 387076
rect 120684 387064 120690 387116
rect 52270 386316 52276 386368
rect 52328 386356 52334 386368
rect 77938 386356 77944 386368
rect 52328 386328 77944 386356
rect 52328 386316 52334 386328
rect 77938 386316 77944 386328
rect 77996 386316 78002 386368
rect 61746 386248 61752 386300
rect 61804 386288 61810 386300
rect 85574 386288 85580 386300
rect 61804 386260 85580 386288
rect 61804 386248 61810 386260
rect 85574 386248 85580 386260
rect 85632 386248 85638 386300
rect 63310 384956 63316 385008
rect 63368 384996 63374 385008
rect 88978 384996 88984 385008
rect 63368 384968 88984 384996
rect 63368 384956 63374 384968
rect 88978 384956 88984 384968
rect 89036 384956 89042 385008
rect 52270 384276 52276 384328
rect 52328 384316 52334 384328
rect 122926 384316 122932 384328
rect 52328 384288 122932 384316
rect 52328 384276 52334 384288
rect 122926 384276 122932 384288
rect 122984 384276 122990 384328
rect 60458 383596 60464 383648
rect 60516 383636 60522 383648
rect 82814 383636 82820 383648
rect 60516 383608 82820 383636
rect 60516 383596 60522 383608
rect 82814 383596 82820 383608
rect 82872 383596 82878 383648
rect 108758 382916 108764 382968
rect 108816 382956 108822 382968
rect 160094 382956 160100 382968
rect 108816 382928 160100 382956
rect 108816 382916 108822 382928
rect 160094 382916 160100 382928
rect 160152 382916 160158 382968
rect 4798 381488 4804 381540
rect 4856 381528 4862 381540
rect 123478 381528 123484 381540
rect 4856 381500 123484 381528
rect 4856 381488 4862 381500
rect 123478 381488 123484 381500
rect 123536 381488 123542 381540
rect 110414 380196 110420 380248
rect 110472 380236 110478 380248
rect 158714 380236 158720 380248
rect 110472 380208 158720 380236
rect 110472 380196 110478 380208
rect 158714 380196 158720 380208
rect 158772 380196 158778 380248
rect 67726 380128 67732 380180
rect 67784 380168 67790 380180
rect 124950 380168 124956 380180
rect 67784 380140 124956 380168
rect 67784 380128 67790 380140
rect 124950 380128 124956 380140
rect 125008 380128 125014 380180
rect 53558 378768 53564 378820
rect 53616 378808 53622 378820
rect 75914 378808 75920 378820
rect 53616 378780 75920 378808
rect 53616 378768 53622 378780
rect 75914 378768 75920 378780
rect 75972 378768 75978 378820
rect 104894 376728 104900 376780
rect 104952 376768 104958 376780
rect 228358 376768 228364 376780
rect 104952 376740 228364 376768
rect 104952 376728 104958 376740
rect 228358 376728 228364 376740
rect 228416 376728 228422 376780
rect 52178 375980 52184 376032
rect 52236 376020 52242 376032
rect 163590 376020 163596 376032
rect 52236 375992 163596 376020
rect 52236 375980 52242 375992
rect 163590 375980 163596 375992
rect 163648 375980 163654 376032
rect 39850 375368 39856 375420
rect 39908 375408 39914 375420
rect 188338 375408 188344 375420
rect 39908 375380 188344 375408
rect 39908 375368 39914 375380
rect 188338 375368 188344 375380
rect 188396 375368 188402 375420
rect 118694 374688 118700 374740
rect 118752 374728 118758 374740
rect 165706 374728 165712 374740
rect 118752 374700 165712 374728
rect 118752 374688 118758 374700
rect 165706 374688 165712 374700
rect 165764 374688 165770 374740
rect 70302 374620 70308 374672
rect 70360 374660 70366 374672
rect 164326 374660 164332 374672
rect 70360 374632 164332 374660
rect 70360 374620 70366 374632
rect 164326 374620 164332 374632
rect 164384 374620 164390 374672
rect 71682 374212 71688 374264
rect 71740 374252 71746 374264
rect 73154 374252 73160 374264
rect 71740 374224 73160 374252
rect 71740 374212 71746 374224
rect 73154 374212 73160 374224
rect 73212 374212 73218 374264
rect 3418 373260 3424 373312
rect 3476 373300 3482 373312
rect 118602 373300 118608 373312
rect 3476 373272 118608 373300
rect 3476 373260 3482 373272
rect 118602 373260 118608 373272
rect 118660 373260 118666 373312
rect 67542 372648 67548 372700
rect 67600 372688 67606 372700
rect 201494 372688 201500 372700
rect 67600 372660 201500 372688
rect 67600 372648 67606 372660
rect 201494 372648 201500 372660
rect 201552 372648 201558 372700
rect 142062 372580 142068 372632
rect 142120 372620 142126 372632
rect 331214 372620 331220 372632
rect 142120 372592 331220 372620
rect 142120 372580 142126 372592
rect 331214 372580 331220 372592
rect 331272 372580 331278 372632
rect 129734 371288 129740 371340
rect 129792 371328 129798 371340
rect 232498 371328 232504 371340
rect 129792 371300 232504 371328
rect 129792 371288 129798 371300
rect 232498 371288 232504 371300
rect 232556 371288 232562 371340
rect 81434 371220 81440 371272
rect 81492 371260 81498 371272
rect 240502 371260 240508 371272
rect 81492 371232 240508 371260
rect 81492 371220 81498 371232
rect 240502 371220 240508 371232
rect 240560 371220 240566 371272
rect 3142 370472 3148 370524
rect 3200 370512 3206 370524
rect 7558 370512 7564 370524
rect 3200 370484 7564 370512
rect 3200 370472 3206 370484
rect 7558 370472 7564 370484
rect 7616 370512 7622 370524
rect 11698 370512 11704 370524
rect 7616 370484 11704 370512
rect 7616 370472 7622 370484
rect 11698 370472 11704 370484
rect 11756 370472 11762 370524
rect 60366 370472 60372 370524
rect 60424 370512 60430 370524
rect 78674 370512 78680 370524
rect 60424 370484 78680 370512
rect 60424 370472 60430 370484
rect 78674 370472 78680 370484
rect 78732 370472 78738 370524
rect 79962 370472 79968 370524
rect 80020 370512 80026 370524
rect 161566 370512 161572 370524
rect 80020 370484 161572 370512
rect 80020 370472 80026 370484
rect 161566 370472 161572 370484
rect 161624 370472 161630 370524
rect 73154 369860 73160 369912
rect 73212 369900 73218 369912
rect 188430 369900 188436 369912
rect 73212 369872 188436 369900
rect 73212 369860 73218 369872
rect 188430 369860 188436 369872
rect 188488 369860 188494 369912
rect 107470 369180 107476 369232
rect 107528 369220 107534 369232
rect 151078 369220 151084 369232
rect 107528 369192 151084 369220
rect 107528 369180 107534 369192
rect 151078 369180 151084 369192
rect 151136 369180 151142 369232
rect 62022 369112 62028 369164
rect 62080 369152 62086 369164
rect 111794 369152 111800 369164
rect 62080 369124 111800 369152
rect 62080 369112 62086 369124
rect 111794 369112 111800 369124
rect 111852 369112 111858 369164
rect 125594 368908 125600 368960
rect 125652 368948 125658 368960
rect 126238 368948 126244 368960
rect 125652 368920 126244 368948
rect 125652 368908 125658 368920
rect 126238 368908 126244 368920
rect 126296 368908 126302 368960
rect 126238 368500 126244 368552
rect 126296 368540 126302 368552
rect 231118 368540 231124 368552
rect 126296 368512 231124 368540
rect 126296 368500 126302 368512
rect 231118 368500 231124 368512
rect 231176 368500 231182 368552
rect 99282 367752 99288 367804
rect 99340 367792 99346 367804
rect 170398 367792 170404 367804
rect 99340 367764 170404 367792
rect 99340 367752 99346 367764
rect 170398 367752 170404 367764
rect 170456 367752 170462 367804
rect 132494 367072 132500 367124
rect 132552 367112 132558 367124
rect 251266 367112 251272 367124
rect 132552 367084 251272 367112
rect 132552 367072 132558 367084
rect 251266 367072 251272 367084
rect 251324 367072 251330 367124
rect 137278 367004 137284 367056
rect 137336 367044 137342 367056
rect 137830 367044 137836 367056
rect 137336 367016 137836 367044
rect 137336 367004 137342 367016
rect 137830 367004 137836 367016
rect 137888 367004 137894 367056
rect 137830 365780 137836 365832
rect 137888 365820 137894 365832
rect 162118 365820 162124 365832
rect 137888 365792 162124 365820
rect 137888 365780 137894 365792
rect 162118 365780 162124 365792
rect 162176 365780 162182 365832
rect 78674 365712 78680 365764
rect 78732 365752 78738 365764
rect 243170 365752 243176 365764
rect 78732 365724 243176 365752
rect 78732 365712 78738 365724
rect 243170 365712 243176 365724
rect 243228 365712 243234 365764
rect 93118 365644 93124 365696
rect 93176 365684 93182 365696
rect 93670 365684 93676 365696
rect 93176 365656 93676 365684
rect 93176 365644 93182 365656
rect 93670 365644 93676 365656
rect 93728 365684 93734 365696
rect 128354 365684 128360 365696
rect 93728 365656 128360 365684
rect 93728 365644 93734 365656
rect 128354 365644 128360 365656
rect 128412 365684 128418 365696
rect 128998 365684 129004 365696
rect 128412 365656 129004 365684
rect 128412 365644 128418 365656
rect 128998 365644 129004 365656
rect 129056 365644 129062 365696
rect 79318 364964 79324 365016
rect 79376 365004 79382 365016
rect 122926 365004 122932 365016
rect 79376 364976 122932 365004
rect 79376 364964 79382 364976
rect 122926 364964 122932 364976
rect 122984 364964 122990 365016
rect 128354 364964 128360 365016
rect 128412 365004 128418 365016
rect 212902 365004 212908 365016
rect 128412 364976 212908 365004
rect 128412 364964 128418 364976
rect 212902 364964 212908 364976
rect 212960 364964 212966 365016
rect 98730 362992 98736 363044
rect 98788 363032 98794 363044
rect 181530 363032 181536 363044
rect 98788 363004 181536 363032
rect 98788 362992 98794 363004
rect 181530 362992 181536 363004
rect 181588 362992 181594 363044
rect 80054 362924 80060 362976
rect 80112 362964 80118 362976
rect 81342 362964 81348 362976
rect 80112 362936 81348 362964
rect 80112 362924 80118 362936
rect 81342 362924 81348 362936
rect 81400 362964 81406 362976
rect 251174 362964 251180 362976
rect 81400 362936 251180 362964
rect 81400 362924 81406 362936
rect 251174 362924 251180 362936
rect 251232 362924 251238 362976
rect 197998 361672 198004 361684
rect 84166 361644 198004 361672
rect 78766 361564 78772 361616
rect 78824 361604 78830 361616
rect 79962 361604 79968 361616
rect 78824 361576 79968 361604
rect 78824 361564 78830 361576
rect 79962 361564 79968 361576
rect 80020 361604 80026 361616
rect 84166 361604 84194 361644
rect 197998 361632 198004 361644
rect 198056 361632 198062 361684
rect 80020 361576 84194 361604
rect 80020 361564 80026 361576
rect 117222 361564 117228 361616
rect 117280 361604 117286 361616
rect 241514 361604 241520 361616
rect 117280 361576 241520 361604
rect 117280 361564 117286 361576
rect 241514 361564 241520 361576
rect 241572 361564 241578 361616
rect 115198 360204 115204 360256
rect 115256 360244 115262 360256
rect 115842 360244 115848 360256
rect 115256 360216 115848 360244
rect 115256 360204 115262 360216
rect 115842 360204 115848 360216
rect 115900 360244 115906 360256
rect 214558 360244 214564 360256
rect 115900 360216 214564 360244
rect 115900 360204 115906 360216
rect 214558 360204 214564 360216
rect 214616 360204 214622 360256
rect 71590 359456 71596 359508
rect 71648 359496 71654 359508
rect 123110 359496 123116 359508
rect 71648 359468 123116 359496
rect 71648 359456 71654 359468
rect 123110 359456 123116 359468
rect 123168 359456 123174 359508
rect 122926 358844 122932 358896
rect 122984 358884 122990 358896
rect 186958 358884 186964 358896
rect 122984 358856 186964 358884
rect 122984 358844 122990 358856
rect 186958 358844 186964 358856
rect 187016 358844 187022 358896
rect 124950 358776 124956 358828
rect 125008 358816 125014 358828
rect 224218 358816 224224 358828
rect 125008 358788 224224 358816
rect 125008 358776 125014 358788
rect 224218 358776 224224 358788
rect 224276 358776 224282 358828
rect 105630 358028 105636 358080
rect 105688 358068 105694 358080
rect 155310 358068 155316 358080
rect 105688 358040 155316 358068
rect 105688 358028 105694 358040
rect 155310 358028 155316 358040
rect 155368 358028 155374 358080
rect 155862 357484 155868 357536
rect 155920 357524 155926 357536
rect 176010 357524 176016 357536
rect 155920 357496 176016 357524
rect 155920 357484 155926 357496
rect 176010 357484 176016 357496
rect 176068 357484 176074 357536
rect 140682 357416 140688 357468
rect 140740 357456 140746 357468
rect 207658 357456 207664 357468
rect 140740 357428 207664 357456
rect 140740 357416 140746 357428
rect 207658 357416 207664 357428
rect 207716 357416 207722 357468
rect 70394 356736 70400 356788
rect 70452 356776 70458 356788
rect 71682 356776 71688 356788
rect 70452 356748 71688 356776
rect 70452 356736 70458 356748
rect 71682 356736 71688 356748
rect 71740 356736 71746 356788
rect 102134 356124 102140 356176
rect 102192 356164 102198 356176
rect 193858 356164 193864 356176
rect 102192 356136 193864 356164
rect 102192 356124 102198 356136
rect 193858 356124 193864 356136
rect 193916 356124 193922 356176
rect 71682 356056 71688 356108
rect 71740 356096 71746 356108
rect 238018 356096 238024 356108
rect 71740 356068 238024 356096
rect 71740 356056 71746 356068
rect 238018 356056 238024 356068
rect 238076 356056 238082 356108
rect 90358 354764 90364 354816
rect 90416 354804 90422 354816
rect 191098 354804 191104 354816
rect 90416 354776 191104 354804
rect 90416 354764 90422 354776
rect 191098 354764 191104 354776
rect 191156 354764 191162 354816
rect 128354 354696 128360 354748
rect 128412 354736 128418 354748
rect 230474 354736 230480 354748
rect 128412 354708 230480 354736
rect 128412 354696 128418 354708
rect 230474 354696 230480 354708
rect 230532 354696 230538 354748
rect 134610 353336 134616 353388
rect 134668 353376 134674 353388
rect 138014 353376 138020 353388
rect 134668 353348 138020 353376
rect 134668 353336 134674 353348
rect 138014 353336 138020 353348
rect 138072 353376 138078 353388
rect 169018 353376 169024 353388
rect 138072 353348 169024 353376
rect 138072 353336 138078 353348
rect 169018 353336 169024 353348
rect 169076 353336 169082 353388
rect 65610 353268 65616 353320
rect 65668 353308 65674 353320
rect 67634 353308 67640 353320
rect 65668 353280 67640 353308
rect 65668 353268 65674 353280
rect 67634 353268 67640 353280
rect 67692 353268 67698 353320
rect 69842 353268 69848 353320
rect 69900 353308 69906 353320
rect 184290 353308 184296 353320
rect 69900 353280 184296 353308
rect 69900 353268 69906 353280
rect 184290 353268 184296 353280
rect 184348 353268 184354 353320
rect 202138 352724 202144 352776
rect 202196 352764 202202 352776
rect 202782 352764 202788 352776
rect 202196 352736 202788 352764
rect 202196 352724 202202 352736
rect 202782 352724 202788 352736
rect 202840 352724 202846 352776
rect 97810 352520 97816 352572
rect 97868 352560 97874 352572
rect 154666 352560 154672 352572
rect 97868 352532 154672 352560
rect 97868 352520 97874 352532
rect 154666 352520 154672 352532
rect 154724 352520 154730 352572
rect 202782 352520 202788 352572
rect 202840 352560 202846 352572
rect 580166 352560 580172 352572
rect 202840 352532 580172 352560
rect 202840 352520 202846 352532
rect 580166 352520 580172 352532
rect 580224 352520 580230 352572
rect 144178 351908 144184 351960
rect 144236 351948 144242 351960
rect 146294 351948 146300 351960
rect 144236 351920 146300 351948
rect 144236 351908 144242 351920
rect 146294 351908 146300 351920
rect 146352 351948 146358 351960
rect 195422 351948 195428 351960
rect 146352 351920 195428 351948
rect 146352 351908 146358 351920
rect 195422 351908 195428 351920
rect 195480 351908 195486 351960
rect 104802 351228 104808 351280
rect 104860 351268 104866 351280
rect 120718 351268 120724 351280
rect 104860 351240 120724 351268
rect 104860 351228 104866 351240
rect 120718 351228 120724 351240
rect 120776 351228 120782 351280
rect 110322 351160 110328 351212
rect 110380 351200 110386 351212
rect 155218 351200 155224 351212
rect 110380 351172 155224 351200
rect 110380 351160 110386 351172
rect 155218 351160 155224 351172
rect 155276 351160 155282 351212
rect 85482 350548 85488 350600
rect 85540 350588 85546 350600
rect 90358 350588 90364 350600
rect 85540 350560 90364 350588
rect 85540 350548 85546 350560
rect 90358 350548 90364 350560
rect 90416 350548 90422 350600
rect 123478 350548 123484 350600
rect 123536 350588 123542 350600
rect 177390 350588 177396 350600
rect 123536 350560 177396 350588
rect 123536 350548 123542 350560
rect 177390 350548 177396 350560
rect 177448 350548 177454 350600
rect 63310 349800 63316 349852
rect 63368 349840 63374 349852
rect 71590 349840 71596 349852
rect 63368 349812 71596 349840
rect 63368 349800 63374 349812
rect 71590 349800 71596 349812
rect 71648 349840 71654 349852
rect 222838 349840 222844 349852
rect 71648 349812 222844 349840
rect 71648 349800 71654 349812
rect 222838 349800 222844 349812
rect 222896 349800 222902 349852
rect 118694 349120 118700 349172
rect 118752 349160 118758 349172
rect 119338 349160 119344 349172
rect 118752 349132 119344 349160
rect 118752 349120 118758 349132
rect 119338 349120 119344 349132
rect 119396 349160 119402 349172
rect 249794 349160 249800 349172
rect 119396 349132 249800 349160
rect 119396 349120 119402 349132
rect 249794 349120 249800 349132
rect 249852 349120 249858 349172
rect 92290 349052 92296 349104
rect 92348 349092 92354 349104
rect 118786 349092 118792 349104
rect 92348 349064 118792 349092
rect 92348 349052 92354 349064
rect 118786 349052 118792 349064
rect 118844 349092 118850 349104
rect 119430 349092 119436 349104
rect 118844 349064 119436 349092
rect 118844 349052 118850 349064
rect 119430 349052 119436 349064
rect 119488 349052 119494 349104
rect 122742 348440 122748 348492
rect 122800 348480 122806 348492
rect 130470 348480 130476 348492
rect 122800 348452 130476 348480
rect 122800 348440 122806 348452
rect 130470 348440 130476 348452
rect 130528 348440 130534 348492
rect 96522 348372 96528 348424
rect 96580 348412 96586 348424
rect 128446 348412 128452 348424
rect 96580 348384 128452 348412
rect 96580 348372 96586 348384
rect 128446 348372 128452 348384
rect 128504 348372 128510 348424
rect 142798 348372 142804 348424
rect 142856 348412 142862 348424
rect 156046 348412 156052 348424
rect 142856 348384 156052 348412
rect 142856 348372 142862 348384
rect 156046 348372 156052 348384
rect 156104 348372 156110 348424
rect 133138 347760 133144 347812
rect 133196 347800 133202 347812
rect 222930 347800 222936 347812
rect 133196 347772 222936 347800
rect 133196 347760 133202 347772
rect 222930 347760 222936 347772
rect 222988 347760 222994 347812
rect 78582 347012 78588 347064
rect 78640 347052 78646 347064
rect 93118 347052 93124 347064
rect 78640 347024 93124 347052
rect 78640 347012 78646 347024
rect 93118 347012 93124 347024
rect 93176 347012 93182 347064
rect 96430 347012 96436 347064
rect 96488 347052 96494 347064
rect 116578 347052 116584 347064
rect 96488 347024 116584 347052
rect 96488 347012 96494 347024
rect 116578 347012 116584 347024
rect 116636 347012 116642 347064
rect 135162 346468 135168 346520
rect 135220 346508 135226 346520
rect 198090 346508 198096 346520
rect 135220 346480 198096 346508
rect 135220 346468 135226 346480
rect 198090 346468 198096 346480
rect 198148 346468 198154 346520
rect 66070 346400 66076 346452
rect 66128 346440 66134 346452
rect 196710 346440 196716 346452
rect 66128 346412 196716 346440
rect 66128 346400 66134 346412
rect 196710 346400 196716 346412
rect 196768 346400 196774 346452
rect 3142 346332 3148 346384
rect 3200 346372 3206 346384
rect 33778 346372 33784 346384
rect 3200 346344 33784 346372
rect 3200 346332 3206 346344
rect 33778 346332 33784 346344
rect 33836 346332 33842 346384
rect 92382 345652 92388 345704
rect 92440 345692 92446 345704
rect 121454 345692 121460 345704
rect 92440 345664 121460 345692
rect 92440 345652 92446 345664
rect 121454 345652 121460 345664
rect 121512 345652 121518 345704
rect 143534 345108 143540 345160
rect 143592 345148 143598 345160
rect 183002 345148 183008 345160
rect 143592 345120 183008 345148
rect 143592 345108 143598 345120
rect 183002 345108 183008 345120
rect 183060 345108 183066 345160
rect 67266 345040 67272 345092
rect 67324 345080 67330 345092
rect 224310 345080 224316 345092
rect 67324 345052 224316 345080
rect 67324 345040 67330 345052
rect 224310 345040 224316 345052
rect 224368 345040 224374 345092
rect 49602 344292 49608 344344
rect 49660 344332 49666 344344
rect 82814 344332 82820 344344
rect 49660 344304 82820 344332
rect 49660 344292 49666 344304
rect 82814 344292 82820 344304
rect 82872 344292 82878 344344
rect 99374 343680 99380 343732
rect 99432 343720 99438 343732
rect 100110 343720 100116 343732
rect 99432 343692 100116 343720
rect 99432 343680 99438 343692
rect 100110 343680 100116 343692
rect 100168 343720 100174 343732
rect 167638 343720 167644 343732
rect 100168 343692 167644 343720
rect 100168 343680 100174 343692
rect 167638 343680 167644 343692
rect 167696 343680 167702 343732
rect 97258 343612 97264 343664
rect 97316 343652 97322 343664
rect 246298 343652 246304 343664
rect 97316 343624 246304 343652
rect 97316 343612 97322 343624
rect 246298 343612 246304 343624
rect 246356 343612 246362 343664
rect 134242 342320 134248 342372
rect 134300 342360 134306 342372
rect 173342 342360 173348 342372
rect 134300 342332 173348 342360
rect 134300 342320 134306 342332
rect 173342 342320 173348 342332
rect 173400 342320 173406 342372
rect 67634 342252 67640 342304
rect 67692 342292 67698 342304
rect 167730 342292 167736 342304
rect 67692 342264 167736 342292
rect 67692 342252 67698 342264
rect 167730 342252 167736 342264
rect 167788 342252 167794 342304
rect 141418 341068 141424 341080
rect 122806 341040 141424 341068
rect 61746 340960 61752 341012
rect 61804 341000 61810 341012
rect 122806 341000 122834 341040
rect 141418 341028 141424 341040
rect 141476 341028 141482 341080
rect 61804 340972 122834 341000
rect 61804 340960 61810 340972
rect 140774 340960 140780 341012
rect 140832 341000 140838 341012
rect 225598 341000 225604 341012
rect 140832 340972 225604 341000
rect 140832 340960 140838 340972
rect 225598 340960 225604 340972
rect 225656 340960 225662 341012
rect 60550 340892 60556 340944
rect 60608 340932 60614 340944
rect 145374 340932 145380 340944
rect 60608 340904 145380 340932
rect 60608 340892 60614 340904
rect 145374 340892 145380 340904
rect 145432 340892 145438 340944
rect 146202 340892 146208 340944
rect 146260 340932 146266 340944
rect 357434 340932 357440 340944
rect 146260 340904 357440 340932
rect 146260 340892 146266 340904
rect 357434 340892 357440 340904
rect 357492 340892 357498 340944
rect 74350 340144 74356 340196
rect 74408 340184 74414 340196
rect 93210 340184 93216 340196
rect 74408 340156 93216 340184
rect 74408 340144 74414 340156
rect 93210 340144 93216 340156
rect 93268 340144 93274 340196
rect 63218 339532 63224 339584
rect 63276 339572 63282 339584
rect 159450 339572 159456 339584
rect 63276 339544 159456 339572
rect 63276 339532 63282 339544
rect 159450 339532 159456 339544
rect 159508 339532 159514 339584
rect 115934 339464 115940 339516
rect 115992 339504 115998 339516
rect 244274 339504 244280 339516
rect 115992 339476 244280 339504
rect 115992 339464 115998 339476
rect 244274 339464 244280 339476
rect 244332 339464 244338 339516
rect 137002 338172 137008 338224
rect 137060 338212 137066 338224
rect 164878 338212 164884 338224
rect 137060 338184 164884 338212
rect 137060 338172 137066 338184
rect 164878 338172 164884 338184
rect 164936 338172 164942 338224
rect 71774 338104 71780 338156
rect 71832 338144 71838 338156
rect 216030 338144 216036 338156
rect 71832 338116 216036 338144
rect 71832 338104 71838 338116
rect 216030 338104 216036 338116
rect 216088 338104 216094 338156
rect 66162 337424 66168 337476
rect 66220 337464 66226 337476
rect 74534 337464 74540 337476
rect 66220 337436 74540 337464
rect 66220 337424 66226 337436
rect 74534 337424 74540 337436
rect 74592 337424 74598 337476
rect 54846 337356 54852 337408
rect 54904 337396 54910 337408
rect 86954 337396 86960 337408
rect 54904 337368 86960 337396
rect 54904 337356 54910 337368
rect 86954 337356 86960 337368
rect 87012 337356 87018 337408
rect 120074 337356 120080 337408
rect 120132 337396 120138 337408
rect 140774 337396 140780 337408
rect 120132 337368 140780 337396
rect 120132 337356 120138 337368
rect 140774 337356 140780 337368
rect 140832 337356 140838 337408
rect 92842 336812 92848 336864
rect 92900 336852 92906 336864
rect 178770 336852 178776 336864
rect 92900 336824 178776 336852
rect 92900 336812 92906 336824
rect 178770 336812 178776 336824
rect 178828 336812 178834 336864
rect 146938 336744 146944 336796
rect 146996 336784 147002 336796
rect 252646 336784 252652 336796
rect 146996 336756 252652 336784
rect 146996 336744 147002 336756
rect 252646 336744 252652 336756
rect 252704 336744 252710 336796
rect 113174 335996 113180 336048
rect 113232 336036 113238 336048
rect 139394 336036 139400 336048
rect 113232 336008 139400 336036
rect 113232 335996 113238 336008
rect 139394 335996 139400 336008
rect 139452 335996 139458 336048
rect 140774 335996 140780 336048
rect 140832 336036 140838 336048
rect 146938 336036 146944 336048
rect 140832 336008 146944 336036
rect 140832 335996 140838 336008
rect 146938 335996 146944 336008
rect 146996 335996 147002 336048
rect 61838 335384 61844 335436
rect 61896 335424 61902 335436
rect 203518 335424 203524 335436
rect 61896 335396 203524 335424
rect 61896 335384 61902 335396
rect 203518 335384 203524 335396
rect 203576 335384 203582 335436
rect 149146 335316 149152 335368
rect 149204 335356 149210 335368
rect 335354 335356 335360 335368
rect 149204 335328 335360 335356
rect 149204 335316 149210 335328
rect 335354 335316 335360 335328
rect 335412 335316 335418 335368
rect 60458 334568 60464 334620
rect 60516 334608 60522 334620
rect 113174 334608 113180 334620
rect 60516 334580 113180 334608
rect 60516 334568 60522 334580
rect 113174 334568 113180 334580
rect 113232 334568 113238 334620
rect 115658 334024 115664 334076
rect 115716 334064 115722 334076
rect 173250 334064 173256 334076
rect 115716 334036 173256 334064
rect 115716 334024 115722 334036
rect 173250 334024 173256 334036
rect 173308 334024 173314 334076
rect 59262 333956 59268 334008
rect 59320 333996 59326 334008
rect 89898 333996 89904 334008
rect 59320 333968 89904 333996
rect 59320 333956 59326 333968
rect 89898 333956 89904 333968
rect 89956 333956 89962 334008
rect 104250 333956 104256 334008
rect 104308 333996 104314 334008
rect 220170 333996 220176 334008
rect 104308 333968 220176 333996
rect 104308 333956 104314 333968
rect 220170 333956 220176 333968
rect 220228 333956 220234 334008
rect 91554 333072 91560 333124
rect 91612 333112 91618 333124
rect 94498 333112 94504 333124
rect 91612 333084 94504 333112
rect 91612 333072 91618 333084
rect 94498 333072 94504 333084
rect 94556 333072 94562 333124
rect 113634 332664 113640 332716
rect 113692 332704 113698 332716
rect 160830 332704 160836 332716
rect 113692 332676 160836 332704
rect 113692 332664 113698 332676
rect 160830 332664 160836 332676
rect 160888 332664 160894 332716
rect 71866 332596 71872 332648
rect 71924 332636 71930 332648
rect 73062 332636 73068 332648
rect 71924 332608 73068 332636
rect 71924 332596 71930 332608
rect 73062 332596 73068 332608
rect 73120 332636 73126 332648
rect 133322 332636 133328 332648
rect 73120 332608 133328 332636
rect 73120 332596 73126 332608
rect 133322 332596 133328 332608
rect 133380 332596 133386 332648
rect 133414 332596 133420 332648
rect 133472 332636 133478 332648
rect 170490 332636 170496 332648
rect 133472 332608 170496 332636
rect 133472 332596 133478 332608
rect 170490 332596 170496 332608
rect 170548 332596 170554 332648
rect 91002 332528 91008 332580
rect 91060 332568 91066 332580
rect 93854 332568 93860 332580
rect 91060 332540 93860 332568
rect 91060 332528 91066 332540
rect 93854 332528 93860 332540
rect 93912 332528 93918 332580
rect 207658 331848 207664 331900
rect 207716 331888 207722 331900
rect 239398 331888 239404 331900
rect 207716 331860 239404 331888
rect 207716 331848 207722 331860
rect 239398 331848 239404 331860
rect 239456 331848 239462 331900
rect 129734 331440 129740 331492
rect 129792 331480 129798 331492
rect 130102 331480 130108 331492
rect 129792 331452 130108 331480
rect 129792 331440 129798 331452
rect 130102 331440 130108 331452
rect 130160 331440 130166 331492
rect 53742 331304 53748 331356
rect 53800 331344 53806 331356
rect 129734 331344 129740 331356
rect 53800 331316 129740 331344
rect 53800 331304 53806 331316
rect 129734 331304 129740 331316
rect 129792 331304 129798 331356
rect 141234 331304 141240 331356
rect 141292 331344 141298 331356
rect 157426 331344 157432 331356
rect 141292 331316 157432 331344
rect 141292 331304 141298 331316
rect 157426 331304 157432 331316
rect 157484 331304 157490 331356
rect 107194 331236 107200 331288
rect 107252 331276 107258 331288
rect 189718 331276 189724 331288
rect 107252 331248 189724 331276
rect 107252 331236 107258 331248
rect 189718 331236 189724 331248
rect 189776 331236 189782 331288
rect 56502 331168 56508 331220
rect 56560 331208 56566 331220
rect 123478 331208 123484 331220
rect 56560 331180 123484 331208
rect 56560 331168 56566 331180
rect 123478 331168 123484 331180
rect 123536 331168 123542 331220
rect 78674 331100 78680 331152
rect 78732 331140 78738 331152
rect 79318 331140 79324 331152
rect 78732 331112 79324 331140
rect 78732 331100 78738 331112
rect 79318 331100 79324 331112
rect 79376 331100 79382 331152
rect 82722 331100 82728 331152
rect 82780 331140 82786 331152
rect 83458 331140 83464 331152
rect 82780 331112 83464 331140
rect 82780 331100 82786 331112
rect 83458 331100 83464 331112
rect 83516 331100 83522 331152
rect 95786 331100 95792 331152
rect 95844 331140 95850 331152
rect 96430 331140 96436 331152
rect 95844 331112 96436 331140
rect 95844 331100 95850 331112
rect 96430 331100 96436 331112
rect 96488 331100 96494 331152
rect 117774 331100 117780 331152
rect 117832 331140 117838 331152
rect 118602 331140 118608 331152
rect 117832 331112 118608 331140
rect 117832 331100 117838 331112
rect 118602 331100 118608 331112
rect 118660 331100 118666 331152
rect 118694 331100 118700 331152
rect 118752 331140 118758 331152
rect 119430 331140 119436 331152
rect 118752 331112 119436 331140
rect 118752 331100 118758 331112
rect 119430 331100 119436 331112
rect 119488 331100 119494 331152
rect 137830 331100 137836 331152
rect 137888 331140 137894 331152
rect 139394 331140 139400 331152
rect 137888 331112 139400 331140
rect 137888 331100 137894 331112
rect 139394 331100 139400 331112
rect 139452 331100 139458 331152
rect 144178 331100 144184 331152
rect 144236 331140 144242 331152
rect 144822 331140 144828 331152
rect 144236 331112 144828 331140
rect 144236 331100 144242 331112
rect 144822 331100 144828 331112
rect 144880 331100 144886 331152
rect 198090 330556 198096 330608
rect 198148 330596 198154 330608
rect 247126 330596 247132 330608
rect 198148 330568 247132 330596
rect 198148 330556 198154 330568
rect 247126 330556 247132 330568
rect 247184 330556 247190 330608
rect 25498 330488 25504 330540
rect 25556 330528 25562 330540
rect 56502 330528 56508 330540
rect 25556 330500 56508 330528
rect 25556 330488 25562 330500
rect 56502 330488 56508 330500
rect 56560 330488 56566 330540
rect 85850 330488 85856 330540
rect 85908 330528 85914 330540
rect 97258 330528 97264 330540
rect 85908 330500 97264 330528
rect 85908 330488 85914 330500
rect 97258 330488 97264 330500
rect 97316 330488 97322 330540
rect 101490 330488 101496 330540
rect 101548 330528 101554 330540
rect 132586 330528 132592 330540
rect 101548 330500 132592 330528
rect 101548 330488 101554 330500
rect 132586 330488 132592 330500
rect 132644 330488 132650 330540
rect 157426 330488 157432 330540
rect 157484 330528 157490 330540
rect 213822 330528 213828 330540
rect 157484 330500 213828 330528
rect 157484 330488 157490 330500
rect 213822 330488 213828 330500
rect 213880 330488 213886 330540
rect 107746 330352 107752 330404
rect 107804 330392 107810 330404
rect 108022 330392 108028 330404
rect 107804 330364 108028 330392
rect 107804 330352 107810 330364
rect 108022 330352 108028 330364
rect 108080 330352 108086 330404
rect 127710 330352 127716 330404
rect 127768 330392 127774 330404
rect 133414 330392 133420 330404
rect 127768 330364 133420 330392
rect 127768 330352 127774 330364
rect 133414 330352 133420 330364
rect 133472 330352 133478 330404
rect 139210 330352 139216 330404
rect 139268 330392 139274 330404
rect 143442 330392 143448 330404
rect 139268 330364 143448 330392
rect 139268 330352 139274 330364
rect 143442 330352 143448 330364
rect 143500 330352 143506 330404
rect 97258 330080 97264 330132
rect 97316 330120 97322 330132
rect 98730 330120 98736 330132
rect 97316 330092 98736 330120
rect 97316 330080 97322 330092
rect 98730 330080 98736 330092
rect 98788 330080 98794 330132
rect 100018 330080 100024 330132
rect 100076 330120 100082 330132
rect 101398 330120 101404 330132
rect 100076 330092 101404 330120
rect 100076 330080 100082 330092
rect 101398 330080 101404 330092
rect 101456 330080 101462 330132
rect 110598 330080 110604 330132
rect 110656 330120 110662 330132
rect 111702 330120 111708 330132
rect 110656 330092 111708 330120
rect 110656 330080 110662 330092
rect 111702 330080 111708 330092
rect 111760 330080 111766 330132
rect 88610 329944 88616 329996
rect 88668 329984 88674 329996
rect 89622 329984 89628 329996
rect 88668 329956 89628 329984
rect 88668 329944 88674 329956
rect 89622 329944 89628 329956
rect 89680 329944 89686 329996
rect 63402 329808 63408 329860
rect 63460 329848 63466 329860
rect 74534 329848 74540 329860
rect 63460 329820 74540 329848
rect 63460 329808 63466 329820
rect 74534 329808 74540 329820
rect 74592 329808 74598 329860
rect 136910 329808 136916 329860
rect 136968 329848 136974 329860
rect 137922 329848 137928 329860
rect 136968 329820 137928 329848
rect 136968 329808 136974 329820
rect 137922 329808 137928 329820
rect 137980 329808 137986 329860
rect 149054 329808 149060 329860
rect 149112 329848 149118 329860
rect 154298 329848 154304 329860
rect 149112 329820 154304 329848
rect 149112 329808 149118 329820
rect 154298 329808 154304 329820
rect 154356 329808 154362 329860
rect 154574 329808 154580 329860
rect 154632 329848 154638 329860
rect 159358 329848 159364 329860
rect 154632 329820 159364 329848
rect 154632 329808 154638 329820
rect 159358 329808 159364 329820
rect 159416 329808 159422 329860
rect 50522 329740 50528 329792
rect 50580 329780 50586 329792
rect 50798 329780 50804 329792
rect 50580 329752 50804 329780
rect 50580 329740 50586 329752
rect 50798 329740 50804 329752
rect 50856 329780 50862 329792
rect 135162 329780 135168 329792
rect 50856 329752 135168 329780
rect 50856 329740 50862 329752
rect 135162 329740 135168 329752
rect 135220 329740 135226 329792
rect 36538 329060 36544 329112
rect 36596 329100 36602 329112
rect 50522 329100 50528 329112
rect 36596 329072 50528 329100
rect 36596 329060 36602 329072
rect 50522 329060 50528 329072
rect 50580 329060 50586 329112
rect 133414 329060 133420 329112
rect 133472 329100 133478 329112
rect 184198 329100 184204 329112
rect 133472 329072 184204 329100
rect 133472 329060 133478 329072
rect 184198 329060 184204 329072
rect 184256 329060 184262 329112
rect 32398 328448 32404 328500
rect 32456 328488 32462 328500
rect 124950 328488 124956 328500
rect 32456 328460 124956 328488
rect 32456 328448 32462 328460
rect 124950 328448 124956 328460
rect 125008 328448 125014 328500
rect 143442 328448 143448 328500
rect 143500 328488 143506 328500
rect 147398 328488 147404 328500
rect 143500 328460 147404 328488
rect 143500 328448 143506 328460
rect 147398 328448 147404 328460
rect 147456 328448 147462 328500
rect 148962 328448 148968 328500
rect 149020 328488 149026 328500
rect 177482 328488 177488 328500
rect 149020 328460 177488 328488
rect 149020 328448 149026 328460
rect 177482 328448 177488 328460
rect 177540 328448 177546 328500
rect 67818 328380 67824 328432
rect 67876 328420 67882 328432
rect 71866 328420 71872 328432
rect 67876 328392 71872 328420
rect 67876 328380 67882 328392
rect 71866 328380 71872 328392
rect 71924 328380 71930 328432
rect 151722 327768 151728 327820
rect 151780 327808 151786 327820
rect 162210 327808 162216 327820
rect 151780 327780 162216 327808
rect 151780 327768 151786 327780
rect 162210 327768 162216 327780
rect 162268 327768 162274 327820
rect 153930 327700 153936 327752
rect 153988 327740 153994 327752
rect 164970 327740 164976 327752
rect 153988 327712 164976 327740
rect 153988 327700 153994 327712
rect 164970 327700 164976 327712
rect 165028 327700 165034 327752
rect 76466 327156 76472 327208
rect 76524 327196 76530 327208
rect 154390 327196 154396 327208
rect 76524 327168 154396 327196
rect 76524 327156 76530 327168
rect 154390 327156 154396 327168
rect 154448 327156 154454 327208
rect 22738 327088 22744 327140
rect 22796 327128 22802 327140
rect 122926 327128 122932 327140
rect 22796 327100 122932 327128
rect 22796 327088 22802 327100
rect 122926 327088 122932 327100
rect 122984 327128 122990 327140
rect 123662 327128 123668 327140
rect 122984 327100 123668 327128
rect 122984 327088 122990 327100
rect 123662 327088 123668 327100
rect 123720 327088 123726 327140
rect 154298 327088 154304 327140
rect 154356 327128 154362 327140
rect 154850 327128 154856 327140
rect 154356 327100 154856 327128
rect 154356 327088 154362 327100
rect 154850 327088 154856 327100
rect 154908 327088 154914 327140
rect 68646 327020 68652 327072
rect 68704 327060 68710 327072
rect 99374 327060 99380 327072
rect 68704 327032 99380 327060
rect 68704 327020 68710 327032
rect 99374 327020 99380 327032
rect 99432 327060 99438 327072
rect 100110 327060 100116 327072
rect 99432 327032 100116 327060
rect 99432 327020 99438 327032
rect 100110 327020 100116 327032
rect 100168 327020 100174 327072
rect 133322 327020 133328 327072
rect 133380 327060 133386 327072
rect 141234 327060 141240 327072
rect 133380 327032 141240 327060
rect 133380 327020 133386 327032
rect 141234 327020 141240 327032
rect 141292 327020 141298 327072
rect 141418 327020 141424 327072
rect 141476 327060 141482 327072
rect 141476 327032 142154 327060
rect 141476 327020 141482 327032
rect 68554 326952 68560 327004
rect 68612 326992 68618 327004
rect 69382 326992 69388 327004
rect 68612 326964 69388 326992
rect 68612 326952 68618 326964
rect 69382 326952 69388 326964
rect 69440 326952 69446 327004
rect 70026 326952 70032 327004
rect 70084 326992 70090 327004
rect 76558 326992 76564 327004
rect 70084 326964 76564 326992
rect 70084 326952 70090 326964
rect 76558 326952 76564 326964
rect 76616 326952 76622 327004
rect 67726 326884 67732 326936
rect 67784 326924 67790 326936
rect 69566 326924 69572 326936
rect 67784 326896 69572 326924
rect 67784 326884 67790 326896
rect 69566 326884 69572 326896
rect 69624 326884 69630 326936
rect 142126 326924 142154 327032
rect 152090 327020 152096 327072
rect 152148 327060 152154 327072
rect 154390 327060 154396 327072
rect 152148 327032 154396 327060
rect 152148 327020 152154 327032
rect 154390 327020 154396 327032
rect 154448 327020 154454 327072
rect 147398 326952 147404 327004
rect 147456 326992 147462 327004
rect 147456 326964 161474 326992
rect 147456 326952 147462 326964
rect 153102 326924 153108 326936
rect 142126 326896 153108 326924
rect 153102 326884 153108 326896
rect 153160 326884 153166 326936
rect 154298 326884 154304 326936
rect 154356 326924 154362 326936
rect 155862 326924 155868 326936
rect 154356 326896 155868 326924
rect 154356 326884 154362 326896
rect 155862 326884 155868 326896
rect 155920 326884 155926 326936
rect 161446 326380 161474 326964
rect 242158 326380 242164 326392
rect 161446 326352 242164 326380
rect 242158 326340 242164 326352
rect 242216 326340 242222 326392
rect 59078 325660 59084 325712
rect 59136 325700 59142 325712
rect 67174 325700 67180 325712
rect 59136 325672 67180 325700
rect 59136 325660 59142 325672
rect 67174 325660 67180 325672
rect 67232 325660 67238 325712
rect 156414 325660 156420 325712
rect 156472 325700 156478 325712
rect 360194 325700 360200 325712
rect 156472 325672 360200 325700
rect 156472 325660 156478 325672
rect 360194 325660 360200 325672
rect 360252 325660 360258 325712
rect 67358 325592 67364 325644
rect 67416 325632 67422 325644
rect 67726 325632 67732 325644
rect 67416 325604 67732 325632
rect 67416 325592 67422 325604
rect 67726 325592 67732 325604
rect 67784 325592 67790 325644
rect 157150 325320 157156 325372
rect 157208 325360 157214 325372
rect 158714 325360 158720 325372
rect 157208 325332 158720 325360
rect 157208 325320 157214 325332
rect 158714 325320 158720 325332
rect 158772 325320 158778 325372
rect 157242 324912 157248 324964
rect 157300 324952 157306 324964
rect 203610 324952 203616 324964
rect 157300 324924 203616 324952
rect 157300 324912 157306 324924
rect 203610 324912 203616 324924
rect 203668 324912 203674 324964
rect 52362 324300 52368 324352
rect 52420 324340 52426 324352
rect 66898 324340 66904 324352
rect 52420 324312 66904 324340
rect 52420 324300 52426 324312
rect 66898 324300 66904 324312
rect 66956 324300 66962 324352
rect 60642 322940 60648 322992
rect 60700 322980 60706 322992
rect 66806 322980 66812 322992
rect 60700 322952 66812 322980
rect 60700 322940 60706 322952
rect 66806 322940 66812 322952
rect 66864 322940 66870 322992
rect 156874 322940 156880 322992
rect 156932 322980 156938 322992
rect 204990 322980 204996 322992
rect 156932 322952 204996 322980
rect 156932 322940 156938 322952
rect 204990 322940 204996 322952
rect 205048 322940 205054 322992
rect 176010 322260 176016 322312
rect 176068 322300 176074 322312
rect 189810 322300 189816 322312
rect 176068 322272 189816 322300
rect 176068 322260 176074 322272
rect 189810 322260 189816 322272
rect 189868 322260 189874 322312
rect 158714 322192 158720 322244
rect 158772 322232 158778 322244
rect 248414 322232 248420 322244
rect 158772 322204 248420 322232
rect 158772 322192 158778 322204
rect 248414 322192 248420 322204
rect 248472 322192 248478 322244
rect 61930 321580 61936 321632
rect 61988 321620 61994 321632
rect 61988 321592 64874 321620
rect 61988 321580 61994 321592
rect 64846 321552 64874 321592
rect 157242 321580 157248 321632
rect 157300 321620 157306 321632
rect 163682 321620 163688 321632
rect 157300 321592 163688 321620
rect 157300 321580 157306 321592
rect 163682 321580 163688 321592
rect 163740 321580 163746 321632
rect 65610 321552 65616 321564
rect 64846 321524 65616 321552
rect 65610 321512 65616 321524
rect 65668 321552 65674 321564
rect 66438 321552 66444 321564
rect 65668 321524 66444 321552
rect 65668 321512 65674 321524
rect 66438 321512 66444 321524
rect 66496 321512 66502 321564
rect 155862 320900 155868 320952
rect 155920 320940 155926 320952
rect 196618 320940 196624 320952
rect 155920 320912 196624 320940
rect 155920 320900 155926 320912
rect 196618 320900 196624 320912
rect 196676 320900 196682 320952
rect 67358 320832 67364 320884
rect 67416 320872 67422 320884
rect 68278 320872 68284 320884
rect 67416 320844 68284 320872
rect 67416 320832 67422 320844
rect 68278 320832 68284 320844
rect 68336 320832 68342 320884
rect 178678 320832 178684 320884
rect 178736 320872 178742 320884
rect 236638 320872 236644 320884
rect 178736 320844 236644 320872
rect 178736 320832 178742 320844
rect 236638 320832 236644 320844
rect 236696 320832 236702 320884
rect 218698 320152 218704 320204
rect 218756 320192 218762 320204
rect 219342 320192 219348 320204
rect 218756 320164 219348 320192
rect 218756 320152 218762 320164
rect 219342 320152 219348 320164
rect 219400 320192 219406 320204
rect 295978 320192 295984 320204
rect 219400 320164 295984 320192
rect 219400 320152 219406 320164
rect 295978 320152 295984 320164
rect 296036 320152 296042 320204
rect 4062 320084 4068 320136
rect 4120 320124 4126 320136
rect 4798 320124 4804 320136
rect 4120 320096 4804 320124
rect 4120 320084 4126 320096
rect 4798 320084 4804 320096
rect 4856 320084 4862 320136
rect 167730 319472 167736 319524
rect 167788 319512 167794 319524
rect 206370 319512 206376 319524
rect 167788 319484 206376 319512
rect 167788 319472 167794 319484
rect 206370 319472 206376 319484
rect 206428 319472 206434 319524
rect 164878 319404 164884 319456
rect 164936 319444 164942 319456
rect 238110 319444 238116 319456
rect 164936 319416 238116 319444
rect 164936 319404 164942 319416
rect 238110 319404 238116 319416
rect 238168 319404 238174 319456
rect 64414 318792 64420 318844
rect 64472 318832 64478 318844
rect 66806 318832 66812 318844
rect 64472 318804 66812 318832
rect 64472 318792 64478 318804
rect 66806 318792 66812 318804
rect 66864 318792 66870 318844
rect 157242 318792 157248 318844
rect 157300 318832 157306 318844
rect 160922 318832 160928 318844
rect 157300 318804 160928 318832
rect 157300 318792 157306 318804
rect 160922 318792 160928 318804
rect 160980 318792 160986 318844
rect 208486 318792 208492 318844
rect 208544 318832 208550 318844
rect 209130 318832 209136 318844
rect 208544 318804 209136 318832
rect 208544 318792 208550 318804
rect 209130 318792 209136 318804
rect 209188 318832 209194 318844
rect 284938 318832 284944 318844
rect 209188 318804 284944 318832
rect 209188 318792 209194 318804
rect 284938 318792 284944 318804
rect 284996 318792 285002 318844
rect 219710 318384 219716 318436
rect 219768 318424 219774 318436
rect 220170 318424 220176 318436
rect 219768 318396 220176 318424
rect 219768 318384 219774 318396
rect 220170 318384 220176 318396
rect 220228 318384 220234 318436
rect 11698 318044 11704 318096
rect 11756 318084 11762 318096
rect 53834 318084 53840 318096
rect 11756 318056 53840 318084
rect 11756 318044 11762 318056
rect 53834 318044 53840 318056
rect 53892 318044 53898 318096
rect 164970 318044 164976 318096
rect 165028 318084 165034 318096
rect 224862 318084 224868 318096
rect 165028 318056 224868 318084
rect 165028 318044 165034 318056
rect 224862 318044 224868 318056
rect 224920 318044 224926 318096
rect 56502 317500 56508 317552
rect 56560 317540 56566 317552
rect 66806 317540 66812 317552
rect 56560 317512 66812 317540
rect 56560 317500 56566 317512
rect 66806 317500 66812 317512
rect 66864 317500 66870 317552
rect 53834 317432 53840 317484
rect 53892 317472 53898 317484
rect 54938 317472 54944 317484
rect 53892 317444 54944 317472
rect 53892 317432 53898 317444
rect 54938 317432 54944 317444
rect 54996 317472 55002 317484
rect 66898 317472 66904 317484
rect 54996 317444 66904 317472
rect 54996 317432 55002 317444
rect 66898 317432 66904 317444
rect 66956 317432 66962 317484
rect 219710 317432 219716 317484
rect 219768 317472 219774 317484
rect 304994 317472 305000 317484
rect 219768 317444 305000 317472
rect 219768 317432 219774 317444
rect 304994 317432 305000 317444
rect 305052 317432 305058 317484
rect 157242 317364 157248 317416
rect 157300 317404 157306 317416
rect 161566 317404 161572 317416
rect 157300 317376 161572 317404
rect 157300 317364 157306 317376
rect 161566 317364 161572 317376
rect 161624 317404 161630 317416
rect 162762 317404 162768 317416
rect 161624 317376 162768 317404
rect 161624 317364 161630 317376
rect 162762 317364 162768 317376
rect 162820 317364 162826 317416
rect 162762 316752 162768 316804
rect 162820 316792 162826 316804
rect 173158 316792 173164 316804
rect 162820 316764 173164 316792
rect 162820 316752 162826 316764
rect 173158 316752 173164 316764
rect 173216 316752 173222 316804
rect 178770 316752 178776 316804
rect 178828 316792 178834 316804
rect 249058 316792 249064 316804
rect 178828 316764 249064 316792
rect 178828 316752 178834 316764
rect 249058 316752 249064 316764
rect 249116 316752 249122 316804
rect 163774 316684 163780 316736
rect 163832 316724 163838 316736
rect 242250 316724 242256 316736
rect 163832 316696 242256 316724
rect 163832 316684 163838 316696
rect 242250 316684 242256 316696
rect 242308 316684 242314 316736
rect 63310 315936 63316 315988
rect 63368 315976 63374 315988
rect 66806 315976 66812 315988
rect 63368 315948 66812 315976
rect 63368 315936 63374 315948
rect 66806 315936 66812 315948
rect 66864 315936 66870 315988
rect 157242 315324 157248 315376
rect 157300 315364 157306 315376
rect 164326 315364 164332 315376
rect 157300 315336 164332 315364
rect 157300 315324 157306 315336
rect 164326 315324 164332 315336
rect 164384 315324 164390 315376
rect 35158 315256 35164 315308
rect 35216 315296 35222 315308
rect 63310 315296 63316 315308
rect 35216 315268 63316 315296
rect 35216 315256 35222 315268
rect 63310 315256 63316 315268
rect 63368 315256 63374 315308
rect 160922 315256 160928 315308
rect 160980 315296 160986 315308
rect 246022 315296 246028 315308
rect 160980 315268 246028 315296
rect 160980 315256 160986 315268
rect 246022 315256 246028 315268
rect 246080 315256 246086 315308
rect 156782 314644 156788 314696
rect 156840 314684 156846 314696
rect 160738 314684 160744 314696
rect 156840 314656 160744 314684
rect 156840 314644 156846 314656
rect 160738 314644 160744 314656
rect 160796 314644 160802 314696
rect 164326 314644 164332 314696
rect 164384 314684 164390 314696
rect 165062 314684 165068 314696
rect 164384 314656 165068 314684
rect 164384 314644 164390 314656
rect 165062 314644 165068 314656
rect 165120 314644 165126 314696
rect 224862 314644 224868 314696
rect 224920 314684 224926 314696
rect 269758 314684 269764 314696
rect 224920 314656 269764 314684
rect 224920 314644 224926 314656
rect 269758 314644 269764 314656
rect 269816 314644 269822 314696
rect 158070 313896 158076 313948
rect 158128 313936 158134 313948
rect 199470 313936 199476 313948
rect 158128 313908 199476 313936
rect 158128 313896 158134 313908
rect 199470 313896 199476 313908
rect 199528 313896 199534 313948
rect 226334 313352 226340 313404
rect 226392 313392 226398 313404
rect 288434 313392 288440 313404
rect 226392 313364 288440 313392
rect 226392 313352 226398 313364
rect 288434 313352 288440 313364
rect 288492 313352 288498 313404
rect 53558 313284 53564 313336
rect 53616 313324 53622 313336
rect 61654 313324 61660 313336
rect 53616 313296 61660 313324
rect 53616 313284 53622 313296
rect 61654 313284 61660 313296
rect 61712 313324 61718 313336
rect 66898 313324 66904 313336
rect 61712 313296 66904 313324
rect 61712 313284 61718 313296
rect 66898 313284 66904 313296
rect 66956 313284 66962 313336
rect 187050 313284 187056 313336
rect 187108 313324 187114 313336
rect 187602 313324 187608 313336
rect 187108 313296 187608 313324
rect 187108 313284 187114 313296
rect 187602 313284 187608 313296
rect 187660 313324 187666 313336
rect 268378 313324 268384 313336
rect 187660 313296 268384 313324
rect 187660 313284 187666 313296
rect 268378 313284 268384 313296
rect 268436 313284 268442 313336
rect 64782 313216 64788 313268
rect 64840 313256 64846 313268
rect 66806 313256 66812 313268
rect 64840 313228 66812 313256
rect 64840 313216 64846 313228
rect 66806 313216 66812 313228
rect 66864 313216 66870 313268
rect 189810 312536 189816 312588
rect 189868 312576 189874 312588
rect 239214 312576 239220 312588
rect 189868 312548 239220 312576
rect 189868 312536 189874 312548
rect 239214 312536 239220 312548
rect 239272 312536 239278 312588
rect 246298 312536 246304 312588
rect 246356 312576 246362 312588
rect 255406 312576 255412 312588
rect 246356 312548 255412 312576
rect 246356 312536 246362 312548
rect 255406 312536 255412 312548
rect 255464 312536 255470 312588
rect 156414 311856 156420 311908
rect 156472 311896 156478 311908
rect 218698 311896 218704 311908
rect 156472 311868 218704 311896
rect 156472 311856 156478 311868
rect 218698 311856 218704 311868
rect 218756 311856 218762 311908
rect 220078 311856 220084 311908
rect 220136 311896 220142 311908
rect 220722 311896 220728 311908
rect 220136 311868 220728 311896
rect 220136 311856 220142 311868
rect 220722 311856 220728 311868
rect 220780 311896 220786 311908
rect 304258 311896 304264 311908
rect 220780 311868 304264 311896
rect 220780 311856 220786 311868
rect 304258 311856 304264 311868
rect 304316 311856 304322 311908
rect 64598 311788 64604 311840
rect 64656 311828 64662 311840
rect 66438 311828 66444 311840
rect 64656 311800 66444 311828
rect 64656 311788 64662 311800
rect 66438 311788 66444 311800
rect 66496 311788 66502 311840
rect 184290 311176 184296 311228
rect 184348 311216 184354 311228
rect 230014 311216 230020 311228
rect 184348 311188 230020 311216
rect 184348 311176 184354 311188
rect 230014 311176 230020 311188
rect 230072 311176 230078 311228
rect 173342 311108 173348 311160
rect 173400 311148 173406 311160
rect 235994 311148 236000 311160
rect 173400 311120 236000 311148
rect 173400 311108 173406 311120
rect 235994 311108 236000 311120
rect 236052 311108 236058 311160
rect 157242 310496 157248 310548
rect 157300 310536 157306 310548
rect 180150 310536 180156 310548
rect 157300 310508 180156 310536
rect 157300 310496 157306 310508
rect 180150 310496 180156 310508
rect 180208 310496 180214 310548
rect 204990 310428 204996 310480
rect 205048 310468 205054 310480
rect 209958 310468 209964 310480
rect 205048 310440 209964 310468
rect 205048 310428 205054 310440
rect 209958 310428 209964 310440
rect 210016 310428 210022 310480
rect 170490 309748 170496 309800
rect 170548 309788 170554 309800
rect 191190 309788 191196 309800
rect 170548 309760 191196 309788
rect 170548 309748 170554 309760
rect 191190 309748 191196 309760
rect 191248 309748 191254 309800
rect 156138 309272 156144 309324
rect 156196 309312 156202 309324
rect 158070 309312 158076 309324
rect 156196 309284 158076 309312
rect 156196 309272 156202 309284
rect 158070 309272 158076 309284
rect 158128 309272 158134 309324
rect 157242 309204 157248 309256
rect 157300 309244 157306 309256
rect 199378 309244 199384 309256
rect 157300 309216 199384 309244
rect 157300 309204 157306 309216
rect 199378 309204 199384 309216
rect 199436 309204 199442 309256
rect 53650 309136 53656 309188
rect 53708 309176 53714 309188
rect 66806 309176 66812 309188
rect 53708 309148 66812 309176
rect 53708 309136 53714 309148
rect 66806 309136 66812 309148
rect 66864 309136 66870 309188
rect 191282 309136 191288 309188
rect 191340 309176 191346 309188
rect 254026 309176 254032 309188
rect 191340 309148 254032 309176
rect 191340 309136 191346 309148
rect 254026 309136 254032 309148
rect 254084 309136 254090 309188
rect 167822 309068 167828 309120
rect 167880 309108 167886 309120
rect 168282 309108 168288 309120
rect 167880 309080 168288 309108
rect 167880 309068 167886 309080
rect 168282 309068 168288 309080
rect 168340 309108 168346 309120
rect 226334 309108 226340 309120
rect 168340 309080 226340 309108
rect 168340 309068 168346 309080
rect 226334 309068 226340 309080
rect 226392 309068 226398 309120
rect 156690 308456 156696 308508
rect 156748 308496 156754 308508
rect 159542 308496 159548 308508
rect 156748 308468 159548 308496
rect 156748 308456 156754 308468
rect 159542 308456 159548 308468
rect 159600 308456 159606 308508
rect 14458 308388 14464 308440
rect 14516 308428 14522 308440
rect 67634 308428 67640 308440
rect 14516 308400 67640 308428
rect 14516 308388 14522 308400
rect 67634 308388 67640 308400
rect 67692 308388 67698 308440
rect 193122 307844 193128 307896
rect 193180 307884 193186 307896
rect 280154 307884 280160 307896
rect 193180 307856 280160 307884
rect 193180 307844 193186 307856
rect 280154 307844 280160 307856
rect 280212 307844 280218 307896
rect 228450 307776 228456 307828
rect 228508 307816 228514 307828
rect 228910 307816 228916 307828
rect 228508 307788 228916 307816
rect 228508 307776 228514 307788
rect 228910 307776 228916 307788
rect 228968 307816 228974 307828
rect 324406 307816 324412 307828
rect 228968 307788 324412 307816
rect 228968 307776 228974 307788
rect 324406 307776 324412 307788
rect 324464 307776 324470 307828
rect 154758 307708 154764 307760
rect 154816 307748 154822 307760
rect 155310 307748 155316 307760
rect 154816 307720 155316 307748
rect 154816 307708 154822 307720
rect 155310 307708 155316 307720
rect 155368 307708 155374 307760
rect 239214 307708 239220 307760
rect 239272 307748 239278 307760
rect 242526 307748 242532 307760
rect 239272 307720 242532 307748
rect 239272 307708 239278 307720
rect 242526 307708 242532 307720
rect 242584 307708 242590 307760
rect 18598 307028 18604 307080
rect 18656 307068 18662 307080
rect 66714 307068 66720 307080
rect 18656 307040 66720 307068
rect 18656 307028 18662 307040
rect 66714 307028 66720 307040
rect 66772 307028 66778 307080
rect 207750 306416 207756 306468
rect 207808 306456 207814 306468
rect 286410 306456 286416 306468
rect 207808 306428 286416 306456
rect 207808 306416 207814 306428
rect 286410 306416 286416 306428
rect 286468 306416 286474 306468
rect 61746 306348 61752 306400
rect 61804 306388 61810 306400
rect 66990 306388 66996 306400
rect 61804 306360 66996 306388
rect 61804 306348 61810 306360
rect 66990 306348 66996 306360
rect 67048 306348 67054 306400
rect 154758 306348 154764 306400
rect 154816 306388 154822 306400
rect 239490 306388 239496 306400
rect 154816 306360 239496 306388
rect 154816 306348 154822 306360
rect 239490 306348 239496 306360
rect 239548 306348 239554 306400
rect 3418 306280 3424 306332
rect 3476 306320 3482 306332
rect 36538 306320 36544 306332
rect 3476 306292 36544 306320
rect 3476 306280 3482 306292
rect 36538 306280 36544 306292
rect 36596 306280 36602 306332
rect 63218 306280 63224 306332
rect 63276 306320 63282 306332
rect 66898 306320 66904 306332
rect 63276 306292 66904 306320
rect 63276 306280 63282 306292
rect 66898 306280 66904 306292
rect 66956 306280 66962 306332
rect 157242 306280 157248 306332
rect 157300 306320 157306 306332
rect 160186 306320 160192 306332
rect 157300 306292 160192 306320
rect 157300 306280 157306 306292
rect 160186 306280 160192 306292
rect 160244 306280 160250 306332
rect 160186 305668 160192 305720
rect 160244 305708 160250 305720
rect 174722 305708 174728 305720
rect 160244 305680 174728 305708
rect 160244 305668 160250 305680
rect 174722 305668 174728 305680
rect 174780 305668 174786 305720
rect 163682 305600 163688 305652
rect 163740 305640 163746 305652
rect 245746 305640 245752 305652
rect 163740 305612 245752 305640
rect 163740 305600 163746 305612
rect 245746 305600 245752 305612
rect 245804 305600 245810 305652
rect 184382 304988 184388 305040
rect 184440 305028 184446 305040
rect 258074 305028 258080 305040
rect 184440 305000 258080 305028
rect 184440 304988 184446 305000
rect 258074 304988 258080 305000
rect 258132 304988 258138 305040
rect 157242 304240 157248 304292
rect 157300 304280 157306 304292
rect 183462 304280 183468 304292
rect 157300 304252 183468 304280
rect 157300 304240 157306 304252
rect 183462 304240 183468 304252
rect 183520 304240 183526 304292
rect 224310 304240 224316 304292
rect 224368 304280 224374 304292
rect 247034 304280 247040 304292
rect 224368 304252 247040 304280
rect 224368 304240 224374 304252
rect 247034 304240 247040 304252
rect 247092 304240 247098 304292
rect 157242 303696 157248 303748
rect 157300 303736 157306 303748
rect 215938 303736 215944 303748
rect 157300 303708 215944 303736
rect 157300 303696 157306 303708
rect 215938 303696 215944 303708
rect 215996 303696 216002 303748
rect 57882 303628 57888 303680
rect 57940 303668 57946 303680
rect 66254 303668 66260 303680
rect 57940 303640 66260 303668
rect 57940 303628 57946 303640
rect 66254 303628 66260 303640
rect 66312 303628 66318 303680
rect 197170 303628 197176 303680
rect 197228 303668 197234 303680
rect 198182 303668 198188 303680
rect 197228 303640 198188 303668
rect 197228 303628 197234 303640
rect 198182 303628 198188 303640
rect 198240 303668 198246 303680
rect 262950 303668 262956 303680
rect 198240 303640 262956 303668
rect 198240 303628 198246 303640
rect 262950 303628 262956 303640
rect 263008 303628 263014 303680
rect 60458 303560 60464 303612
rect 60516 303600 60522 303612
rect 66806 303600 66812 303612
rect 60516 303572 66812 303600
rect 60516 303560 60522 303572
rect 66806 303560 66812 303572
rect 66864 303560 66870 303612
rect 183462 302268 183468 302320
rect 183520 302308 183526 302320
rect 261478 302308 261484 302320
rect 183520 302280 261484 302308
rect 183520 302268 183526 302280
rect 261478 302268 261484 302280
rect 261536 302268 261542 302320
rect 157242 302200 157248 302252
rect 157300 302240 157306 302252
rect 243906 302240 243912 302252
rect 157300 302212 243912 302240
rect 157300 302200 157306 302212
rect 243906 302200 243912 302212
rect 243964 302200 243970 302252
rect 64690 302132 64696 302184
rect 64748 302172 64754 302184
rect 66806 302172 66812 302184
rect 64748 302144 66812 302172
rect 64748 302132 64754 302144
rect 66806 302132 66812 302144
rect 66864 302132 66870 302184
rect 197262 301520 197268 301572
rect 197320 301560 197326 301572
rect 198090 301560 198096 301572
rect 197320 301532 198096 301560
rect 197320 301520 197326 301532
rect 198090 301520 198096 301532
rect 198148 301520 198154 301572
rect 193858 301316 193864 301368
rect 193916 301356 193922 301368
rect 194502 301356 194508 301368
rect 193916 301328 194508 301356
rect 193916 301316 193922 301328
rect 194502 301316 194508 301328
rect 194560 301316 194566 301368
rect 215294 300908 215300 300960
rect 215352 300948 215358 300960
rect 216030 300948 216036 300960
rect 215352 300920 216036 300948
rect 215352 300908 215358 300920
rect 216030 300908 216036 300920
rect 216088 300948 216094 300960
rect 266998 300948 267004 300960
rect 216088 300920 267004 300948
rect 216088 300908 216094 300920
rect 266998 300908 267004 300920
rect 267056 300908 267062 300960
rect 194502 300840 194508 300892
rect 194560 300880 194566 300892
rect 246298 300880 246304 300892
rect 194560 300852 246304 300880
rect 194560 300840 194566 300852
rect 246298 300840 246304 300852
rect 246356 300840 246362 300892
rect 60550 300772 60556 300824
rect 60608 300812 60614 300824
rect 66806 300812 66812 300824
rect 60608 300784 66812 300812
rect 60608 300772 60614 300784
rect 66806 300772 66812 300784
rect 66864 300772 66870 300824
rect 63310 299548 63316 299600
rect 63368 299588 63374 299600
rect 66254 299588 66260 299600
rect 63368 299560 66260 299588
rect 63368 299548 63374 299560
rect 66254 299548 66260 299560
rect 66312 299548 66318 299600
rect 157242 299548 157248 299600
rect 157300 299588 157306 299600
rect 244458 299588 244464 299600
rect 157300 299560 244464 299588
rect 157300 299548 157306 299560
rect 244458 299548 244464 299560
rect 244516 299548 244522 299600
rect 162394 299480 162400 299532
rect 162452 299520 162458 299532
rect 256694 299520 256700 299532
rect 162452 299492 256700 299520
rect 162452 299480 162458 299492
rect 256694 299480 256700 299492
rect 256752 299480 256758 299532
rect 157242 299412 157248 299464
rect 157300 299452 157306 299464
rect 165706 299452 165712 299464
rect 157300 299424 165712 299452
rect 157300 299412 157306 299424
rect 165706 299412 165712 299424
rect 165764 299452 165770 299464
rect 166074 299452 166080 299464
rect 165764 299424 166080 299452
rect 165764 299412 165770 299424
rect 166074 299412 166080 299424
rect 166132 299412 166138 299464
rect 231118 299412 231124 299464
rect 231176 299452 231182 299464
rect 233142 299452 233148 299464
rect 231176 299424 233148 299452
rect 231176 299412 231182 299424
rect 233142 299412 233148 299424
rect 233200 299412 233206 299464
rect 214558 298800 214564 298852
rect 214616 298840 214622 298852
rect 227438 298840 227444 298852
rect 214616 298812 227444 298840
rect 214616 298800 214622 298812
rect 227438 298800 227444 298812
rect 227496 298800 227502 298852
rect 50798 298732 50804 298784
rect 50856 298772 50862 298784
rect 66898 298772 66904 298784
rect 50856 298744 66904 298772
rect 50856 298732 50862 298744
rect 66898 298732 66904 298744
rect 66956 298732 66962 298784
rect 166074 298732 166080 298784
rect 166132 298772 166138 298784
rect 216582 298772 216588 298784
rect 166132 298744 216588 298772
rect 166132 298732 166138 298744
rect 216582 298732 216588 298744
rect 216640 298732 216646 298784
rect 233142 298120 233148 298172
rect 233200 298160 233206 298172
rect 583754 298160 583760 298172
rect 233200 298132 583760 298160
rect 233200 298120 233206 298132
rect 583754 298120 583760 298132
rect 583812 298120 583818 298172
rect 238202 298052 238208 298104
rect 238260 298092 238266 298104
rect 238662 298092 238668 298104
rect 238260 298064 238668 298092
rect 238260 298052 238266 298064
rect 238662 298052 238668 298064
rect 238720 298052 238726 298104
rect 156782 296760 156788 296812
rect 156840 296800 156846 296812
rect 252738 296800 252744 296812
rect 156840 296772 252744 296800
rect 156840 296760 156846 296772
rect 252738 296760 252744 296772
rect 252796 296760 252802 296812
rect 238662 296692 238668 296744
rect 238720 296732 238726 296744
rect 582558 296732 582564 296744
rect 238720 296704 582564 296732
rect 238720 296692 238726 296704
rect 582558 296692 582564 296704
rect 582616 296692 582622 296744
rect 39942 296624 39948 296676
rect 40000 296664 40006 296676
rect 66438 296664 66444 296676
rect 40000 296636 66444 296664
rect 40000 296624 40006 296636
rect 66438 296624 66444 296636
rect 66496 296624 66502 296676
rect 157242 295944 157248 295996
rect 157300 295984 157306 295996
rect 161474 295984 161480 295996
rect 157300 295956 161480 295984
rect 157300 295944 157306 295956
rect 161474 295944 161480 295956
rect 161532 295984 161538 295996
rect 162762 295984 162768 295996
rect 161532 295956 162768 295984
rect 161532 295944 161538 295956
rect 162762 295944 162768 295956
rect 162820 295944 162826 295996
rect 203702 295400 203708 295452
rect 203760 295440 203766 295452
rect 277394 295440 277400 295452
rect 203760 295412 277400 295440
rect 203760 295400 203766 295412
rect 277394 295400 277400 295412
rect 277452 295400 277458 295452
rect 200574 295332 200580 295384
rect 200632 295372 200638 295384
rect 216674 295372 216680 295384
rect 200632 295344 216680 295372
rect 200632 295332 200638 295344
rect 216674 295332 216680 295344
rect 216732 295332 216738 295384
rect 233970 295332 233976 295384
rect 234028 295372 234034 295384
rect 582466 295372 582472 295384
rect 234028 295344 582472 295372
rect 234028 295332 234034 295344
rect 582466 295332 582472 295344
rect 582524 295332 582530 295384
rect 156414 295264 156420 295316
rect 156472 295304 156478 295316
rect 169754 295304 169760 295316
rect 156472 295276 169760 295304
rect 156472 295264 156478 295276
rect 169754 295264 169760 295276
rect 169812 295264 169818 295316
rect 216582 294652 216588 294704
rect 216640 294692 216646 294704
rect 228358 294692 228364 294704
rect 216640 294664 228364 294692
rect 216640 294652 216646 294664
rect 228358 294652 228364 294664
rect 228416 294652 228422 294704
rect 169754 294584 169760 294636
rect 169812 294624 169818 294636
rect 204346 294624 204352 294636
rect 169812 294596 204352 294624
rect 169812 294584 169818 294596
rect 204346 294584 204352 294596
rect 204404 294584 204410 294636
rect 218698 294584 218704 294636
rect 218756 294624 218762 294636
rect 245838 294624 245844 294636
rect 218756 294596 245844 294624
rect 218756 294584 218762 294596
rect 245838 294584 245844 294596
rect 245896 294584 245902 294636
rect 246298 294584 246304 294636
rect 246356 294624 246362 294636
rect 297358 294624 297364 294636
rect 246356 294596 297364 294624
rect 246356 294584 246362 294596
rect 297358 294584 297364 294596
rect 297416 294584 297422 294636
rect 46842 294040 46848 294092
rect 46900 294080 46906 294092
rect 66254 294080 66260 294092
rect 46900 294052 66260 294080
rect 46900 294040 46906 294052
rect 66254 294040 66260 294052
rect 66312 294040 66318 294092
rect 33778 293972 33784 294024
rect 33836 294012 33842 294024
rect 67542 294012 67548 294024
rect 33836 293984 67548 294012
rect 33836 293972 33842 293984
rect 67542 293972 67548 293984
rect 67600 293972 67606 294024
rect 199470 293972 199476 294024
rect 199528 294012 199534 294024
rect 218054 294012 218060 294024
rect 199528 293984 218060 294012
rect 199528 293972 199534 293984
rect 218054 293972 218060 293984
rect 218112 293972 218118 294024
rect 240870 293972 240876 294024
rect 240928 294012 240934 294024
rect 583202 294012 583208 294024
rect 240928 293984 583208 294012
rect 240928 293972 240934 293984
rect 583202 293972 583208 293984
rect 583260 293972 583266 294024
rect 215938 293292 215944 293344
rect 215996 293332 216002 293344
rect 236730 293332 236736 293344
rect 215996 293304 236736 293332
rect 215996 293292 216002 293304
rect 236730 293292 236736 293304
rect 236788 293292 236794 293344
rect 170398 293224 170404 293276
rect 170456 293264 170462 293276
rect 202782 293264 202788 293276
rect 170456 293236 202788 293264
rect 170456 293224 170462 293236
rect 202782 293224 202788 293236
rect 202840 293264 202846 293276
rect 209958 293264 209964 293276
rect 202840 293236 209964 293264
rect 202840 293224 202846 293236
rect 209958 293224 209964 293236
rect 210016 293224 210022 293276
rect 235166 293224 235172 293276
rect 235224 293264 235230 293276
rect 241514 293264 241520 293276
rect 235224 293236 241520 293264
rect 235224 293224 235230 293236
rect 241514 293224 241520 293236
rect 241572 293264 241578 293276
rect 291838 293264 291844 293276
rect 241572 293236 291844 293264
rect 241572 293224 241578 293236
rect 291838 293224 291844 293236
rect 291896 293224 291902 293276
rect 2774 292816 2780 292868
rect 2832 292856 2838 292868
rect 4798 292856 4804 292868
rect 2832 292828 4804 292856
rect 2832 292816 2838 292828
rect 4798 292816 4804 292828
rect 4856 292816 4862 292868
rect 157242 292544 157248 292596
rect 157300 292584 157306 292596
rect 215478 292584 215484 292596
rect 157300 292556 215484 292584
rect 157300 292544 157306 292556
rect 215478 292544 215484 292556
rect 215536 292544 215542 292596
rect 40678 292476 40684 292528
rect 40736 292516 40742 292528
rect 66806 292516 66812 292528
rect 40736 292488 66812 292516
rect 40736 292476 40742 292488
rect 66806 292476 66812 292488
rect 66864 292476 66870 292528
rect 218054 291796 218060 291848
rect 218112 291836 218118 291848
rect 244366 291836 244372 291848
rect 218112 291808 244372 291836
rect 218112 291796 218118 291808
rect 244366 291796 244372 291808
rect 244424 291796 244430 291848
rect 204346 291592 204352 291644
rect 204404 291632 204410 291644
rect 208578 291632 208584 291644
rect 204404 291604 208584 291632
rect 204404 291592 204410 291604
rect 208578 291592 208584 291604
rect 208636 291592 208642 291644
rect 157242 291252 157248 291304
rect 157300 291292 157306 291304
rect 193950 291292 193956 291304
rect 157300 291264 193956 291292
rect 157300 291252 157306 291264
rect 193950 291252 193956 291264
rect 194008 291252 194014 291304
rect 193858 291184 193864 291236
rect 193916 291224 193922 291236
rect 223022 291224 223028 291236
rect 193916 291196 223028 291224
rect 193916 291184 193922 291196
rect 223022 291184 223028 291196
rect 223080 291184 223086 291236
rect 223574 291184 223580 291236
rect 223632 291224 223638 291236
rect 265618 291224 265624 291236
rect 223632 291196 265624 291224
rect 223632 291184 223638 291196
rect 265618 291184 265624 291196
rect 265676 291184 265682 291236
rect 64690 291116 64696 291168
rect 64748 291156 64754 291168
rect 65518 291156 65524 291168
rect 64748 291128 65524 291156
rect 64748 291116 64754 291128
rect 65518 291116 65524 291128
rect 65576 291116 65582 291168
rect 158070 291116 158076 291168
rect 158128 291156 158134 291168
rect 160738 291156 160744 291168
rect 158128 291128 160744 291156
rect 158128 291116 158134 291128
rect 160738 291116 160744 291128
rect 160796 291116 160802 291168
rect 64690 289892 64696 289944
rect 64748 289932 64754 289944
rect 66806 289932 66812 289944
rect 64748 289904 66812 289932
rect 64748 289892 64754 289904
rect 66806 289892 66812 289904
rect 66864 289892 66870 289944
rect 174538 289892 174544 289944
rect 174596 289932 174602 289944
rect 247218 289932 247224 289944
rect 174596 289904 247224 289932
rect 174596 289892 174602 289904
rect 247218 289892 247224 289904
rect 247276 289892 247282 289944
rect 157242 289824 157248 289876
rect 157300 289864 157306 289876
rect 244550 289864 244556 289876
rect 157300 289836 244556 289864
rect 157300 289824 157306 289836
rect 244550 289824 244556 289836
rect 244608 289824 244614 289876
rect 233878 289756 233884 289808
rect 233936 289796 233942 289808
rect 235534 289796 235540 289808
rect 233936 289768 235540 289796
rect 233936 289756 233942 289768
rect 235534 289756 235540 289768
rect 235592 289756 235598 289808
rect 61838 289212 61844 289264
rect 61896 289252 61902 289264
rect 66254 289252 66260 289264
rect 61896 289224 66260 289252
rect 61896 289212 61902 289224
rect 66254 289212 66260 289224
rect 66312 289212 66318 289264
rect 157242 288464 157248 288516
rect 157300 288504 157306 288516
rect 208394 288504 208400 288516
rect 157300 288476 208400 288504
rect 157300 288464 157306 288476
rect 208394 288464 208400 288476
rect 208452 288464 208458 288516
rect 218054 288464 218060 288516
rect 218112 288504 218118 288516
rect 220630 288504 220636 288516
rect 218112 288476 220636 288504
rect 218112 288464 218118 288476
rect 220630 288464 220636 288476
rect 220688 288504 220694 288516
rect 264238 288504 264244 288516
rect 220688 288476 264244 288504
rect 220688 288464 220694 288476
rect 264238 288464 264244 288476
rect 264296 288464 264302 288516
rect 163682 288396 163688 288448
rect 163740 288436 163746 288448
rect 223574 288436 223580 288448
rect 163740 288408 223580 288436
rect 163740 288396 163746 288408
rect 223574 288396 223580 288408
rect 223632 288396 223638 288448
rect 236730 288396 236736 288448
rect 236788 288436 236794 288448
rect 262858 288436 262864 288448
rect 236788 288408 262864 288436
rect 236788 288396 236794 288408
rect 262858 288396 262864 288408
rect 262916 288396 262922 288448
rect 215478 288328 215484 288380
rect 215536 288368 215542 288380
rect 218054 288368 218060 288380
rect 215536 288340 218060 288368
rect 215536 288328 215542 288340
rect 218054 288328 218060 288340
rect 218112 288328 218118 288380
rect 208394 287648 208400 287700
rect 208452 287688 208458 287700
rect 224678 287688 224684 287700
rect 208452 287660 224684 287688
rect 208452 287648 208458 287660
rect 224678 287648 224684 287660
rect 224736 287648 224742 287700
rect 208394 287512 208400 287564
rect 208452 287552 208458 287564
rect 208578 287552 208584 287564
rect 208452 287524 208584 287552
rect 208452 287512 208458 287524
rect 208578 287512 208584 287524
rect 208636 287512 208642 287564
rect 224678 287104 224684 287156
rect 224736 287144 224742 287156
rect 253198 287144 253204 287156
rect 224736 287116 253204 287144
rect 224736 287104 224742 287116
rect 253198 287104 253204 287116
rect 253256 287104 253262 287156
rect 60550 287036 60556 287088
rect 60608 287076 60614 287088
rect 66806 287076 66812 287088
rect 60608 287048 66812 287076
rect 60608 287036 60614 287048
rect 66806 287036 66812 287048
rect 66864 287036 66870 287088
rect 164878 287036 164884 287088
rect 164936 287076 164942 287088
rect 210878 287076 210884 287088
rect 164936 287048 210884 287076
rect 164936 287036 164942 287048
rect 210878 287036 210884 287048
rect 210936 287036 210942 287088
rect 219434 287036 219440 287088
rect 219492 287076 219498 287088
rect 267734 287076 267740 287088
rect 219492 287048 267740 287076
rect 219492 287036 219498 287048
rect 267734 287036 267740 287048
rect 267792 287036 267798 287088
rect 159450 286288 159456 286340
rect 159508 286328 159514 286340
rect 187050 286328 187056 286340
rect 159508 286300 187056 286328
rect 159508 286288 159514 286300
rect 187050 286288 187056 286300
rect 187108 286288 187114 286340
rect 187602 286288 187608 286340
rect 187660 286328 187666 286340
rect 200758 286328 200764 286340
rect 187660 286300 200764 286328
rect 187660 286288 187666 286300
rect 200758 286288 200764 286300
rect 200816 286288 200822 286340
rect 218698 286288 218704 286340
rect 218756 286328 218762 286340
rect 236454 286328 236460 286340
rect 218756 286300 236460 286328
rect 218756 286288 218762 286300
rect 236454 286288 236460 286300
rect 236512 286288 236518 286340
rect 156138 285880 156144 285932
rect 156196 285920 156202 285932
rect 158070 285920 158076 285932
rect 156196 285892 158076 285920
rect 156196 285880 156202 285892
rect 158070 285880 158076 285892
rect 158128 285880 158134 285932
rect 219342 285880 219348 285932
rect 219400 285920 219406 285932
rect 221182 285920 221188 285932
rect 219400 285892 221188 285920
rect 219400 285880 219406 285892
rect 221182 285880 221188 285892
rect 221240 285880 221246 285932
rect 55122 285744 55128 285796
rect 55180 285784 55186 285796
rect 66990 285784 66996 285796
rect 55180 285756 66996 285784
rect 55180 285744 55186 285756
rect 66990 285744 66996 285756
rect 67048 285744 67054 285796
rect 205542 285784 205548 285796
rect 200086 285756 205548 285784
rect 48222 285676 48228 285728
rect 48280 285716 48286 285728
rect 66806 285716 66812 285728
rect 48280 285688 66812 285716
rect 48280 285676 48286 285688
rect 66806 285676 66812 285688
rect 66864 285676 66870 285728
rect 162302 285676 162308 285728
rect 162360 285716 162366 285728
rect 164234 285716 164240 285728
rect 162360 285688 164240 285716
rect 162360 285676 162366 285688
rect 164234 285676 164240 285688
rect 164292 285676 164298 285728
rect 195514 285676 195520 285728
rect 195572 285716 195578 285728
rect 200086 285716 200114 285756
rect 205542 285744 205548 285756
rect 205600 285744 205606 285796
rect 250438 285784 250444 285796
rect 234264 285756 250444 285784
rect 234264 285728 234292 285756
rect 250438 285744 250444 285756
rect 250496 285744 250502 285796
rect 195572 285688 200114 285716
rect 195572 285676 195578 285688
rect 203150 285676 203156 285728
rect 203208 285716 203214 285728
rect 204162 285716 204168 285728
rect 203208 285688 204168 285716
rect 203208 285676 203214 285688
rect 204162 285676 204168 285688
rect 204220 285676 204226 285728
rect 204898 285676 204904 285728
rect 204956 285716 204962 285728
rect 208118 285716 208124 285728
rect 204956 285688 208124 285716
rect 204956 285676 204962 285688
rect 208118 285676 208124 285688
rect 208176 285676 208182 285728
rect 232590 285676 232596 285728
rect 232648 285716 232654 285728
rect 234246 285716 234252 285728
rect 232648 285688 234252 285716
rect 232648 285676 232654 285688
rect 234246 285676 234252 285688
rect 234304 285676 234310 285728
rect 237558 285676 237564 285728
rect 237616 285716 237622 285728
rect 237926 285716 237932 285728
rect 237616 285688 237932 285716
rect 237616 285676 237622 285688
rect 237926 285676 237932 285688
rect 237984 285716 237990 285728
rect 300118 285716 300124 285728
rect 237984 285688 300124 285716
rect 237984 285676 237990 285688
rect 300118 285676 300124 285688
rect 300176 285676 300182 285728
rect 156782 285608 156788 285660
rect 156840 285648 156846 285660
rect 174538 285648 174544 285660
rect 156840 285620 174544 285648
rect 156840 285608 156846 285620
rect 174538 285608 174544 285620
rect 174596 285608 174602 285660
rect 201494 285268 201500 285320
rect 201552 285308 201558 285320
rect 202414 285308 202420 285320
rect 201552 285280 202420 285308
rect 201552 285268 201558 285280
rect 202414 285268 202420 285280
rect 202472 285268 202478 285320
rect 208394 285268 208400 285320
rect 208452 285308 208458 285320
rect 208670 285308 208676 285320
rect 208452 285280 208676 285308
rect 208452 285268 208458 285280
rect 208670 285268 208676 285280
rect 208728 285268 208734 285320
rect 177482 284996 177488 285048
rect 177540 285036 177546 285048
rect 184290 285036 184296 285048
rect 177540 285008 184296 285036
rect 177540 284996 177546 285008
rect 184290 284996 184296 285008
rect 184348 284996 184354 285048
rect 159542 284928 159548 284980
rect 159600 284968 159606 284980
rect 196710 284968 196716 284980
rect 159600 284940 196716 284968
rect 159600 284928 159606 284940
rect 196710 284928 196716 284940
rect 196768 284928 196774 284980
rect 216674 284928 216680 284980
rect 216732 284968 216738 284980
rect 240042 284968 240048 284980
rect 216732 284940 240048 284968
rect 216732 284928 216738 284940
rect 240042 284928 240048 284940
rect 240100 284928 240106 284980
rect 216766 284724 216772 284776
rect 216824 284764 216830 284776
rect 219434 284764 219440 284776
rect 216824 284736 219440 284764
rect 216824 284724 216830 284736
rect 219434 284724 219440 284736
rect 219492 284724 219498 284776
rect 200114 284384 200120 284436
rect 200172 284424 200178 284436
rect 216766 284424 216772 284436
rect 200172 284396 216772 284424
rect 200172 284384 200178 284396
rect 216766 284384 216772 284396
rect 216824 284384 216830 284436
rect 230750 284384 230756 284436
rect 230808 284424 230814 284436
rect 231118 284424 231124 284436
rect 230808 284396 231124 284424
rect 230808 284384 230814 284396
rect 231118 284384 231124 284396
rect 231176 284424 231182 284436
rect 243906 284424 243912 284436
rect 231176 284396 243912 284424
rect 231176 284384 231182 284396
rect 243906 284384 243912 284396
rect 243964 284384 243970 284436
rect 199562 284316 199568 284368
rect 199620 284356 199626 284368
rect 217318 284356 217324 284368
rect 199620 284328 217324 284356
rect 199620 284316 199626 284328
rect 217318 284316 217324 284328
rect 217376 284316 217382 284368
rect 241974 284316 241980 284368
rect 242032 284356 242038 284368
rect 313918 284356 313924 284368
rect 242032 284328 313924 284356
rect 242032 284316 242038 284328
rect 313918 284316 313924 284328
rect 313976 284316 313982 284368
rect 157242 284248 157248 284300
rect 157300 284288 157306 284300
rect 191282 284288 191288 284300
rect 157300 284260 191288 284288
rect 157300 284248 157306 284260
rect 191282 284248 191288 284260
rect 191340 284248 191346 284300
rect 195974 283908 195980 283960
rect 196032 283948 196038 283960
rect 204346 283948 204352 283960
rect 196032 283920 204352 283948
rect 196032 283908 196038 283920
rect 204346 283908 204352 283920
rect 204404 283908 204410 283960
rect 178770 283840 178776 283892
rect 178828 283880 178834 283892
rect 200114 283880 200120 283892
rect 178828 283852 200120 283880
rect 178828 283840 178834 283852
rect 200114 283840 200120 283852
rect 200172 283840 200178 283892
rect 243906 283840 243912 283892
rect 243964 283880 243970 283892
rect 282914 283880 282920 283892
rect 243964 283852 282920 283880
rect 243964 283840 243970 283852
rect 282914 283840 282920 283852
rect 282972 283840 282978 283892
rect 50982 282888 50988 282940
rect 51040 282928 51046 282940
rect 66622 282928 66628 282940
rect 51040 282900 66628 282928
rect 51040 282888 51046 282900
rect 66622 282888 66628 282900
rect 66680 282888 66686 282940
rect 245378 282888 245384 282940
rect 245436 282928 245442 282940
rect 273254 282928 273260 282940
rect 245436 282900 273260 282928
rect 245436 282888 245442 282900
rect 273254 282888 273260 282900
rect 273312 282888 273318 282940
rect 246114 282820 246120 282872
rect 246172 282860 246178 282872
rect 251358 282860 251364 282872
rect 246172 282832 251364 282860
rect 246172 282820 246178 282832
rect 251358 282820 251364 282832
rect 251416 282860 251422 282872
rect 582834 282860 582840 282872
rect 251416 282832 582840 282860
rect 251416 282820 251422 282832
rect 582834 282820 582840 282832
rect 582892 282820 582898 282872
rect 157242 282616 157248 282668
rect 157300 282656 157306 282668
rect 162394 282656 162400 282668
rect 157300 282628 162400 282656
rect 157300 282616 157306 282628
rect 162394 282616 162400 282628
rect 162452 282616 162458 282668
rect 173342 282208 173348 282260
rect 173400 282248 173406 282260
rect 198734 282248 198740 282260
rect 173400 282220 198740 282248
rect 173400 282208 173406 282220
rect 198734 282208 198740 282220
rect 198792 282208 198798 282260
rect 157150 282140 157156 282192
rect 157208 282180 157214 282192
rect 185762 282180 185768 282192
rect 157208 282152 185768 282180
rect 157208 282140 157214 282152
rect 185762 282140 185768 282152
rect 185820 282140 185826 282192
rect 56410 281528 56416 281580
rect 56468 281568 56474 281580
rect 66346 281568 66352 281580
rect 56468 281540 66352 281568
rect 56468 281528 56474 281540
rect 66346 281528 66352 281540
rect 66404 281528 66410 281580
rect 185762 281528 185768 281580
rect 185820 281568 185826 281580
rect 186222 281568 186228 281580
rect 185820 281540 186228 281568
rect 185820 281528 185826 281540
rect 186222 281528 186228 281540
rect 186280 281568 186286 281580
rect 197354 281568 197360 281580
rect 186280 281540 197360 281568
rect 186280 281528 186286 281540
rect 197354 281528 197360 281540
rect 197412 281528 197418 281580
rect 245654 281528 245660 281580
rect 245712 281568 245718 281580
rect 249702 281568 249708 281580
rect 245712 281540 249708 281568
rect 245712 281528 245718 281540
rect 249702 281528 249708 281540
rect 249760 281528 249766 281580
rect 157242 281460 157248 281512
rect 157300 281500 157306 281512
rect 184382 281500 184388 281512
rect 157300 281472 184388 281500
rect 157300 281460 157306 281472
rect 184382 281460 184388 281472
rect 184440 281460 184446 281512
rect 246114 281460 246120 281512
rect 246172 281500 246178 281512
rect 258166 281500 258172 281512
rect 246172 281472 258172 281500
rect 246172 281460 246178 281472
rect 258166 281460 258172 281472
rect 258224 281500 258230 281512
rect 259362 281500 259368 281512
rect 258224 281472 259368 281500
rect 258224 281460 258230 281472
rect 259362 281460 259368 281472
rect 259420 281460 259426 281512
rect 174722 281392 174728 281444
rect 174780 281432 174786 281444
rect 197354 281432 197360 281444
rect 174780 281404 197360 281432
rect 174780 281392 174786 281404
rect 197354 281392 197360 281404
rect 197412 281392 197418 281444
rect 259362 280780 259368 280832
rect 259420 280820 259426 280832
rect 286318 280820 286324 280832
rect 259420 280792 286324 280820
rect 259420 280780 259426 280792
rect 286318 280780 286324 280792
rect 286376 280780 286382 280832
rect 63126 280168 63132 280220
rect 63184 280208 63190 280220
rect 66806 280208 66812 280220
rect 63184 280180 66812 280208
rect 63184 280168 63190 280180
rect 66806 280168 66812 280180
rect 66864 280168 66870 280220
rect 245654 280168 245660 280220
rect 245712 280208 245718 280220
rect 298738 280208 298744 280220
rect 245712 280180 298744 280208
rect 245712 280168 245718 280180
rect 298738 280168 298744 280180
rect 298796 280168 298802 280220
rect 183462 280100 183468 280152
rect 183520 280140 183526 280152
rect 197354 280140 197360 280152
rect 183520 280112 197360 280140
rect 183520 280100 183526 280112
rect 197354 280100 197360 280112
rect 197412 280100 197418 280152
rect 156966 279624 156972 279676
rect 157024 279664 157030 279676
rect 160922 279664 160928 279676
rect 157024 279636 160928 279664
rect 157024 279624 157030 279636
rect 160922 279624 160928 279636
rect 160980 279624 160986 279676
rect 173434 279420 173440 279472
rect 173492 279460 173498 279472
rect 197446 279460 197452 279472
rect 173492 279432 197452 279460
rect 173492 279420 173498 279432
rect 197446 279420 197452 279432
rect 197504 279420 197510 279472
rect 249702 279420 249708 279472
rect 249760 279460 249766 279472
rect 266354 279460 266360 279472
rect 249760 279432 266360 279460
rect 249760 279420 249766 279432
rect 266354 279420 266360 279432
rect 266412 279420 266418 279472
rect 29638 278740 29644 278792
rect 29696 278780 29702 278792
rect 60458 278780 60464 278792
rect 29696 278752 60464 278780
rect 29696 278740 29702 278752
rect 60458 278740 60464 278752
rect 60516 278780 60522 278792
rect 66622 278780 66628 278792
rect 60516 278752 66628 278780
rect 60516 278740 60522 278752
rect 66622 278740 66628 278752
rect 66680 278740 66686 278792
rect 157058 278740 157064 278792
rect 157116 278780 157122 278792
rect 175182 278780 175188 278792
rect 157116 278752 175188 278780
rect 157116 278740 157122 278752
rect 175182 278740 175188 278752
rect 175240 278740 175246 278792
rect 246114 278740 246120 278792
rect 246172 278780 246178 278792
rect 251358 278780 251364 278792
rect 246172 278752 251364 278780
rect 246172 278740 246178 278752
rect 251358 278740 251364 278752
rect 251416 278780 251422 278792
rect 583570 278780 583576 278792
rect 251416 278752 583576 278780
rect 251416 278740 251422 278752
rect 583570 278740 583576 278752
rect 583628 278740 583634 278792
rect 173250 277992 173256 278044
rect 173308 278032 173314 278044
rect 197262 278032 197268 278044
rect 173308 278004 197268 278032
rect 173308 277992 173314 278004
rect 197262 277992 197268 278004
rect 197320 277992 197326 278044
rect 246114 277992 246120 278044
rect 246172 278032 246178 278044
rect 249978 278032 249984 278044
rect 246172 278004 249984 278032
rect 246172 277992 246178 278004
rect 249978 277992 249984 278004
rect 250036 278032 250042 278044
rect 583386 278032 583392 278044
rect 250036 278004 583392 278032
rect 250036 277992 250042 278004
rect 583386 277992 583392 278004
rect 583444 277992 583450 278044
rect 156506 277380 156512 277432
rect 156564 277420 156570 277432
rect 187050 277420 187056 277432
rect 156564 277392 187056 277420
rect 156564 277380 156570 277392
rect 187050 277380 187056 277392
rect 187108 277380 187114 277432
rect 175182 277312 175188 277364
rect 175240 277352 175246 277364
rect 193122 277352 193128 277364
rect 175240 277324 193128 277352
rect 175240 277312 175246 277324
rect 193122 277312 193128 277324
rect 193180 277312 193186 277364
rect 193122 277108 193128 277160
rect 193180 277148 193186 277160
rect 197354 277148 197360 277160
rect 193180 277120 197360 277148
rect 193180 277108 193186 277120
rect 197354 277108 197360 277120
rect 197412 277108 197418 277160
rect 155310 276632 155316 276684
rect 155368 276672 155374 276684
rect 197998 276672 198004 276684
rect 155368 276644 198004 276672
rect 155368 276632 155374 276644
rect 197998 276632 198004 276644
rect 198056 276632 198062 276684
rect 246022 276632 246028 276684
rect 246080 276672 246086 276684
rect 282178 276672 282184 276684
rect 246080 276644 282184 276672
rect 246080 276632 246086 276644
rect 282178 276632 282184 276644
rect 282236 276632 282242 276684
rect 245838 276224 245844 276276
rect 245896 276264 245902 276276
rect 246022 276264 246028 276276
rect 245896 276236 246028 276264
rect 245896 276224 245902 276236
rect 246022 276224 246028 276236
rect 246080 276224 246086 276276
rect 244274 276088 244280 276140
rect 244332 276128 244338 276140
rect 245654 276128 245660 276140
rect 244332 276100 245660 276128
rect 244332 276088 244338 276100
rect 245654 276088 245660 276100
rect 245712 276088 245718 276140
rect 157242 275952 157248 276004
rect 157300 275992 157306 276004
rect 198274 275992 198280 276004
rect 157300 275964 198280 275992
rect 157300 275952 157306 275964
rect 198274 275952 198280 275964
rect 198332 275952 198338 276004
rect 245930 275952 245936 276004
rect 245988 275992 245994 276004
rect 249886 275992 249892 276004
rect 245988 275964 249892 275992
rect 245988 275952 245994 275964
rect 249886 275952 249892 275964
rect 249944 275992 249950 276004
rect 582650 275992 582656 276004
rect 249944 275964 582656 275992
rect 249944 275952 249950 275964
rect 582650 275952 582656 275964
rect 582708 275952 582714 276004
rect 157242 274660 157248 274712
rect 157300 274700 157306 274712
rect 169202 274700 169208 274712
rect 157300 274672 169208 274700
rect 157300 274660 157306 274672
rect 169202 274660 169208 274672
rect 169260 274660 169266 274712
rect 183094 274660 183100 274712
rect 183152 274700 183158 274712
rect 197446 274700 197452 274712
rect 183152 274672 197452 274700
rect 183152 274660 183158 274672
rect 197446 274660 197452 274672
rect 197504 274660 197510 274712
rect 168282 274592 168288 274644
rect 168340 274632 168346 274644
rect 197354 274632 197360 274644
rect 168340 274604 197360 274632
rect 168340 274592 168346 274604
rect 197354 274592 197360 274604
rect 197412 274592 197418 274644
rect 57606 273912 57612 273964
rect 57664 273952 57670 273964
rect 66254 273952 66260 273964
rect 57664 273924 66260 273952
rect 57664 273912 57670 273924
rect 66254 273912 66260 273924
rect 66312 273912 66318 273964
rect 245930 273912 245936 273964
rect 245988 273952 245994 273964
rect 327166 273952 327172 273964
rect 245988 273924 327172 273952
rect 245988 273912 245994 273924
rect 327166 273912 327172 273924
rect 327224 273912 327230 273964
rect 157242 273232 157248 273284
rect 157300 273272 157306 273284
rect 166442 273272 166448 273284
rect 157300 273244 166448 273272
rect 157300 273232 157306 273244
rect 166442 273232 166448 273244
rect 166500 273232 166506 273284
rect 180242 273232 180248 273284
rect 180300 273272 180306 273284
rect 197354 273272 197360 273284
rect 180300 273244 197360 273272
rect 180300 273232 180306 273244
rect 197354 273232 197360 273244
rect 197412 273232 197418 273284
rect 245838 273232 245844 273284
rect 245896 273272 245902 273284
rect 249886 273272 249892 273284
rect 245896 273244 249892 273272
rect 245896 273232 245902 273244
rect 249886 273232 249892 273244
rect 249944 273232 249950 273284
rect 245930 272552 245936 272604
rect 245988 272592 245994 272604
rect 251266 272592 251272 272604
rect 245988 272564 251272 272592
rect 245988 272552 245994 272564
rect 251266 272552 251272 272564
rect 251324 272592 251330 272604
rect 251818 272592 251824 272604
rect 251324 272564 251824 272592
rect 251324 272552 251330 272564
rect 251818 272552 251824 272564
rect 251876 272552 251882 272604
rect 169110 272484 169116 272536
rect 169168 272524 169174 272536
rect 195882 272524 195888 272536
rect 169168 272496 195888 272524
rect 169168 272484 169174 272496
rect 195882 272484 195888 272496
rect 195940 272484 195946 272536
rect 245838 272484 245844 272536
rect 245896 272524 245902 272536
rect 325694 272524 325700 272536
rect 245896 272496 325700 272524
rect 245896 272484 245902 272496
rect 325694 272484 325700 272496
rect 325752 272484 325758 272536
rect 61746 271940 61752 271992
rect 61804 271980 61810 271992
rect 66990 271980 66996 271992
rect 61804 271952 66996 271980
rect 61804 271940 61810 271952
rect 66990 271940 66996 271952
rect 67048 271940 67054 271992
rect 52178 271872 52184 271924
rect 52236 271912 52242 271924
rect 66806 271912 66812 271924
rect 52236 271884 66812 271912
rect 52236 271872 52242 271884
rect 66806 271872 66812 271884
rect 66864 271872 66870 271924
rect 157242 271872 157248 271924
rect 157300 271912 157306 271924
rect 192478 271912 192484 271924
rect 157300 271884 192484 271912
rect 157300 271872 157306 271884
rect 192478 271872 192484 271884
rect 192536 271872 192542 271924
rect 195882 271872 195888 271924
rect 195940 271912 195946 271924
rect 197354 271912 197360 271924
rect 195940 271884 197360 271912
rect 195940 271872 195946 271884
rect 197354 271872 197360 271884
rect 197412 271872 197418 271924
rect 162486 271124 162492 271176
rect 162544 271164 162550 271176
rect 178770 271164 178776 271176
rect 162544 271136 178776 271164
rect 162544 271124 162550 271136
rect 178770 271124 178776 271136
rect 178828 271124 178834 271176
rect 245746 271124 245752 271176
rect 245804 271164 245810 271176
rect 248598 271164 248604 271176
rect 245804 271136 248604 271164
rect 245804 271124 245810 271136
rect 248598 271124 248604 271136
rect 248656 271124 248662 271176
rect 253198 271124 253204 271176
rect 253256 271164 253262 271176
rect 274634 271164 274640 271176
rect 253256 271136 274640 271164
rect 253256 271124 253262 271136
rect 274634 271124 274640 271136
rect 274692 271124 274698 271176
rect 193030 270580 193036 270632
rect 193088 270620 193094 270632
rect 197446 270620 197452 270632
rect 193088 270592 197452 270620
rect 193088 270580 193094 270592
rect 197446 270580 197452 270592
rect 197504 270580 197510 270632
rect 53742 270512 53748 270564
rect 53800 270552 53806 270564
rect 66806 270552 66812 270564
rect 53800 270524 66812 270552
rect 53800 270512 53806 270524
rect 66806 270512 66812 270524
rect 66864 270512 66870 270564
rect 157242 270512 157248 270564
rect 157300 270552 157306 270564
rect 174538 270552 174544 270564
rect 157300 270524 174544 270552
rect 157300 270512 157306 270524
rect 174538 270512 174544 270524
rect 174596 270512 174602 270564
rect 183002 270512 183008 270564
rect 183060 270552 183066 270564
rect 197354 270552 197360 270564
rect 183060 270524 197360 270552
rect 183060 270512 183066 270524
rect 197354 270512 197360 270524
rect 197412 270512 197418 270564
rect 249058 270552 249064 270564
rect 248386 270524 249064 270552
rect 245654 270444 245660 270496
rect 245712 270484 245718 270496
rect 248386 270484 248414 270524
rect 249058 270512 249064 270524
rect 249116 270552 249122 270564
rect 280246 270552 280252 270564
rect 249116 270524 280252 270552
rect 249116 270512 249122 270524
rect 280246 270512 280252 270524
rect 280304 270512 280310 270564
rect 245712 270456 248414 270484
rect 245712 270444 245718 270456
rect 4062 269764 4068 269816
rect 4120 269804 4126 269816
rect 35894 269804 35900 269816
rect 4120 269776 35900 269804
rect 4120 269764 4126 269776
rect 35894 269764 35900 269776
rect 35952 269764 35958 269816
rect 245930 269764 245936 269816
rect 245988 269804 245994 269816
rect 312170 269804 312176 269816
rect 245988 269776 312176 269804
rect 245988 269764 245994 269776
rect 312170 269764 312176 269776
rect 312228 269764 312234 269816
rect 157242 269152 157248 269204
rect 157300 269192 157306 269204
rect 166258 269192 166264 269204
rect 157300 269164 166264 269192
rect 157300 269152 157306 269164
rect 166258 269152 166264 269164
rect 166316 269152 166322 269204
rect 178862 269152 178868 269204
rect 178920 269192 178926 269204
rect 197354 269192 197360 269204
rect 178920 269164 197360 269192
rect 178920 269152 178926 269164
rect 197354 269152 197360 269164
rect 197412 269152 197418 269204
rect 64506 269084 64512 269136
rect 64564 269124 64570 269136
rect 66438 269124 66444 269136
rect 64564 269096 66444 269124
rect 64564 269084 64570 269096
rect 66438 269084 66444 269096
rect 66496 269084 66502 269136
rect 156782 269084 156788 269136
rect 156840 269124 156846 269136
rect 199654 269124 199660 269136
rect 156840 269096 199660 269124
rect 156840 269084 156846 269096
rect 199654 269084 199660 269096
rect 199712 269084 199718 269136
rect 156506 269016 156512 269068
rect 156564 269056 156570 269068
rect 163682 269056 163688 269068
rect 156564 269028 163688 269056
rect 156564 269016 156570 269028
rect 163682 269016 163688 269028
rect 163740 269016 163746 269068
rect 165062 269016 165068 269068
rect 165120 269056 165126 269068
rect 197354 269056 197360 269068
rect 165120 269028 197360 269056
rect 165120 269016 165126 269028
rect 197354 269016 197360 269028
rect 197412 269016 197418 269068
rect 158162 268336 158168 268388
rect 158220 268376 158226 268388
rect 171226 268376 171232 268388
rect 158220 268348 171232 268376
rect 158220 268336 158226 268348
rect 171226 268336 171232 268348
rect 171284 268376 171290 268388
rect 172422 268376 172428 268388
rect 171284 268348 172428 268376
rect 171284 268336 171290 268348
rect 172422 268336 172428 268348
rect 172480 268336 172486 268388
rect 185578 268336 185584 268388
rect 185636 268376 185642 268388
rect 199562 268376 199568 268388
rect 185636 268348 199568 268376
rect 185636 268336 185642 268348
rect 199562 268336 199568 268348
rect 199620 268336 199626 268388
rect 245930 268336 245936 268388
rect 245988 268376 245994 268388
rect 256786 268376 256792 268388
rect 245988 268348 256792 268376
rect 245988 268336 245994 268348
rect 256786 268336 256792 268348
rect 256844 268336 256850 268388
rect 244458 267724 244464 267776
rect 244516 267764 244522 267776
rect 331306 267764 331312 267776
rect 244516 267736 331312 267764
rect 244516 267724 244522 267736
rect 331306 267724 331312 267736
rect 331364 267724 331370 267776
rect 62022 267656 62028 267708
rect 62080 267696 62086 267708
rect 66438 267696 66444 267708
rect 62080 267668 66444 267696
rect 62080 267656 62086 267668
rect 66438 267656 66444 267668
rect 66496 267656 66502 267708
rect 157242 267656 157248 267708
rect 157300 267696 157306 267708
rect 199470 267696 199476 267708
rect 157300 267668 199476 267696
rect 157300 267656 157306 267668
rect 199470 267656 199476 267668
rect 199528 267656 199534 267708
rect 195422 267452 195428 267504
rect 195480 267492 195486 267504
rect 197354 267492 197360 267504
rect 195480 267464 197360 267492
rect 195480 267452 195486 267464
rect 197354 267452 197360 267464
rect 197412 267452 197418 267504
rect 3418 266976 3424 267028
rect 3476 267016 3482 267028
rect 15838 267016 15844 267028
rect 3476 266988 15844 267016
rect 3476 266976 3482 266988
rect 15838 266976 15844 266988
rect 15896 266976 15902 267028
rect 52086 266976 52092 267028
rect 52144 267016 52150 267028
rect 66898 267016 66904 267028
rect 52144 266988 66904 267016
rect 52144 266976 52150 266988
rect 66898 266976 66904 266988
rect 66956 266976 66962 267028
rect 177390 266976 177396 267028
rect 177448 267016 177454 267028
rect 195054 267016 195060 267028
rect 177448 266988 195060 267016
rect 177448 266976 177454 266988
rect 195054 266976 195060 266988
rect 195112 266976 195118 267028
rect 245930 266976 245936 267028
rect 245988 267016 245994 267028
rect 262214 267016 262220 267028
rect 245988 266988 262220 267016
rect 245988 266976 245994 266988
rect 262214 266976 262220 266988
rect 262272 266976 262278 267028
rect 246022 266364 246028 266416
rect 246080 266404 246086 266416
rect 250070 266404 250076 266416
rect 246080 266376 250076 266404
rect 246080 266364 246086 266376
rect 250070 266364 250076 266376
rect 250128 266364 250134 266416
rect 186958 266296 186964 266348
rect 187016 266336 187022 266348
rect 197354 266336 197360 266348
rect 187016 266308 197360 266336
rect 187016 266296 187022 266308
rect 197354 266296 197360 266308
rect 197412 266296 197418 266348
rect 245746 266296 245752 266348
rect 245804 266336 245810 266348
rect 254118 266336 254124 266348
rect 245804 266308 254124 266336
rect 245804 266296 245810 266308
rect 254118 266296 254124 266308
rect 254176 266336 254182 266348
rect 583110 266336 583116 266348
rect 254176 266308 583116 266336
rect 254176 266296 254182 266308
rect 583110 266296 583116 266308
rect 583168 266296 583174 266348
rect 245838 266228 245844 266280
rect 245896 266268 245902 266280
rect 255406 266268 255412 266280
rect 245896 266240 255412 266268
rect 245896 266228 245902 266240
rect 255406 266228 255412 266240
rect 255464 266228 255470 266280
rect 162394 265616 162400 265668
rect 162452 265656 162458 265668
rect 192570 265656 192576 265668
rect 162452 265628 192576 265656
rect 162452 265616 162458 265628
rect 192570 265616 192576 265628
rect 192628 265616 192634 265668
rect 255406 265616 255412 265668
rect 255464 265656 255470 265668
rect 274726 265656 274732 265668
rect 255464 265628 274732 265656
rect 255464 265616 255470 265628
rect 274726 265616 274732 265628
rect 274784 265616 274790 265668
rect 177850 265140 177856 265192
rect 177908 265180 177914 265192
rect 183094 265180 183100 265192
rect 177908 265152 183100 265180
rect 177908 265140 177914 265152
rect 183094 265140 183100 265152
rect 183152 265140 183158 265192
rect 41322 264936 41328 264988
rect 41380 264976 41386 264988
rect 66806 264976 66812 264988
rect 41380 264948 66812 264976
rect 41380 264936 41386 264948
rect 66806 264936 66812 264948
rect 66864 264936 66870 264988
rect 157242 264936 157248 264988
rect 157300 264976 157306 264988
rect 171870 264976 171876 264988
rect 157300 264948 171876 264976
rect 157300 264936 157306 264948
rect 171870 264936 171876 264948
rect 171928 264936 171934 264988
rect 184198 264868 184204 264920
rect 184256 264908 184262 264920
rect 197354 264908 197360 264920
rect 184256 264880 197360 264908
rect 184256 264868 184262 264880
rect 197354 264868 197360 264880
rect 197412 264868 197418 264920
rect 245930 264868 245936 264920
rect 245988 264908 245994 264920
rect 251174 264908 251180 264920
rect 245988 264880 251180 264908
rect 245988 264868 245994 264880
rect 251174 264868 251180 264880
rect 251232 264868 251238 264920
rect 55030 264188 55036 264240
rect 55088 264228 55094 264240
rect 65978 264228 65984 264240
rect 55088 264200 65984 264228
rect 55088 264188 55094 264200
rect 65978 264188 65984 264200
rect 66036 264228 66042 264240
rect 66438 264228 66444 264240
rect 66036 264200 66444 264228
rect 66036 264188 66042 264200
rect 66438 264188 66444 264200
rect 66496 264188 66502 264240
rect 159542 264188 159548 264240
rect 159600 264228 159606 264240
rect 178678 264228 178684 264240
rect 159600 264200 178684 264228
rect 159600 264188 159606 264200
rect 178678 264188 178684 264200
rect 178736 264188 178742 264240
rect 55030 263644 55036 263696
rect 55088 263684 55094 263696
rect 66806 263684 66812 263696
rect 55088 263656 66812 263684
rect 55088 263644 55094 263656
rect 66806 263644 66812 263656
rect 66864 263644 66870 263696
rect 163682 263576 163688 263628
rect 163740 263616 163746 263628
rect 193122 263616 193128 263628
rect 163740 263588 193128 263616
rect 163740 263576 163746 263588
rect 193122 263576 193128 263588
rect 193180 263616 193186 263628
rect 197354 263616 197360 263628
rect 193180 263588 197360 263616
rect 193180 263576 193186 263588
rect 197354 263576 197360 263588
rect 197412 263576 197418 263628
rect 245838 263576 245844 263628
rect 245896 263616 245902 263628
rect 262214 263616 262220 263628
rect 245896 263588 262220 263616
rect 245896 263576 245902 263588
rect 262214 263576 262220 263588
rect 262272 263576 262278 263628
rect 194042 262896 194048 262948
rect 194100 262936 194106 262948
rect 195514 262936 195520 262948
rect 194100 262908 195520 262936
rect 194100 262896 194106 262908
rect 195514 262896 195520 262908
rect 195572 262896 195578 262948
rect 52270 262828 52276 262880
rect 52328 262868 52334 262880
rect 62114 262868 62120 262880
rect 52328 262840 62120 262868
rect 52328 262828 52334 262840
rect 62114 262828 62120 262840
rect 62172 262828 62178 262880
rect 256786 262828 256792 262880
rect 256844 262868 256850 262880
rect 582650 262868 582656 262880
rect 256844 262840 582656 262868
rect 256844 262828 256850 262840
rect 582650 262828 582656 262840
rect 582708 262828 582714 262880
rect 178678 262284 178684 262336
rect 178736 262324 178742 262336
rect 197354 262324 197360 262336
rect 178736 262296 197360 262324
rect 178736 262284 178742 262296
rect 197354 262284 197360 262296
rect 197412 262284 197418 262336
rect 62114 262216 62120 262268
rect 62172 262256 62178 262268
rect 63218 262256 63224 262268
rect 62172 262228 63224 262256
rect 62172 262216 62178 262228
rect 63218 262216 63224 262228
rect 63276 262256 63282 262268
rect 66806 262256 66812 262268
rect 63276 262228 66812 262256
rect 63276 262216 63282 262228
rect 66806 262216 66812 262228
rect 66864 262216 66870 262268
rect 157242 262216 157248 262268
rect 157300 262256 157306 262268
rect 184198 262256 184204 262268
rect 157300 262228 184204 262256
rect 157300 262216 157306 262228
rect 184198 262216 184204 262228
rect 184256 262216 184262 262268
rect 245930 262216 245936 262268
rect 245988 262256 245994 262268
rect 251174 262256 251180 262268
rect 245988 262228 251180 262256
rect 245988 262216 245994 262228
rect 251174 262216 251180 262228
rect 251232 262216 251238 262268
rect 156782 262148 156788 262200
rect 156840 262188 156846 262200
rect 165614 262188 165620 262200
rect 156840 262160 165620 262188
rect 156840 262148 156846 262160
rect 165614 262148 165620 262160
rect 165672 262148 165678 262200
rect 35894 261468 35900 261520
rect 35952 261508 35958 261520
rect 58986 261508 58992 261520
rect 35952 261480 58992 261508
rect 35952 261468 35958 261480
rect 58986 261468 58992 261480
rect 59044 261468 59050 261520
rect 250438 261468 250444 261520
rect 250496 261508 250502 261520
rect 303614 261508 303620 261520
rect 250496 261480 303620 261508
rect 250496 261468 250502 261480
rect 303614 261468 303620 261480
rect 303672 261468 303678 261520
rect 185670 260924 185676 260976
rect 185728 260964 185734 260976
rect 197354 260964 197360 260976
rect 185728 260936 197360 260964
rect 185728 260924 185734 260936
rect 197354 260924 197360 260936
rect 197412 260924 197418 260976
rect 58986 260856 58992 260908
rect 59044 260896 59050 260908
rect 66806 260896 66812 260908
rect 59044 260868 66812 260896
rect 59044 260856 59050 260868
rect 66806 260856 66812 260868
rect 66864 260856 66870 260908
rect 173250 260856 173256 260908
rect 173308 260896 173314 260908
rect 197446 260896 197452 260908
rect 173308 260868 197452 260896
rect 173308 260856 173314 260868
rect 197446 260856 197452 260868
rect 197504 260856 197510 260908
rect 244918 260856 244924 260908
rect 244976 260896 244982 260908
rect 288526 260896 288532 260908
rect 244976 260868 288532 260896
rect 244976 260856 244982 260868
rect 288526 260856 288532 260868
rect 288584 260856 288590 260908
rect 245930 260788 245936 260840
rect 245988 260828 245994 260840
rect 252738 260828 252744 260840
rect 245988 260800 252744 260828
rect 245988 260788 245994 260800
rect 252738 260788 252744 260800
rect 252796 260828 252802 260840
rect 253014 260828 253020 260840
rect 252796 260800 253020 260828
rect 252796 260788 252802 260800
rect 253014 260788 253020 260800
rect 253072 260788 253078 260840
rect 245838 260176 245844 260228
rect 245896 260216 245902 260228
rect 276014 260216 276020 260228
rect 245896 260188 276020 260216
rect 245896 260176 245902 260188
rect 276014 260176 276020 260188
rect 276072 260176 276078 260228
rect 162210 260108 162216 260160
rect 162268 260148 162274 260160
rect 189902 260148 189908 260160
rect 162268 260120 189908 260148
rect 162268 260108 162274 260120
rect 189902 260108 189908 260120
rect 189960 260108 189966 260160
rect 253014 260108 253020 260160
rect 253072 260148 253078 260160
rect 306650 260148 306656 260160
rect 253072 260120 306656 260148
rect 253072 260108 253078 260120
rect 306650 260108 306656 260120
rect 306708 260108 306714 260160
rect 155402 259428 155408 259480
rect 155460 259468 155466 259480
rect 182082 259468 182088 259480
rect 155460 259440 182088 259468
rect 155460 259428 155466 259440
rect 182082 259428 182088 259440
rect 182140 259468 182146 259480
rect 197354 259468 197360 259480
rect 182140 259440 197360 259468
rect 182140 259428 182146 259440
rect 197354 259428 197360 259440
rect 197412 259428 197418 259480
rect 195054 259360 195060 259412
rect 195112 259400 195118 259412
rect 197446 259400 197452 259412
rect 195112 259372 197452 259400
rect 195112 259360 195118 259372
rect 197446 259360 197452 259372
rect 197504 259360 197510 259412
rect 245838 259360 245844 259412
rect 245896 259400 245902 259412
rect 258074 259400 258080 259412
rect 245896 259372 258080 259400
rect 245896 259360 245902 259372
rect 258074 259360 258080 259372
rect 258132 259400 258138 259412
rect 259362 259400 259368 259412
rect 258132 259372 259368 259400
rect 258132 259360 258138 259372
rect 259362 259360 259368 259372
rect 259420 259360 259426 259412
rect 245930 258680 245936 258732
rect 245988 258720 245994 258732
rect 254026 258720 254032 258732
rect 245988 258692 254032 258720
rect 245988 258680 245994 258692
rect 254026 258680 254032 258692
rect 254084 258680 254090 258732
rect 259362 258680 259368 258732
rect 259420 258720 259426 258732
rect 293218 258720 293224 258732
rect 259420 258692 293224 258720
rect 259420 258680 259426 258692
rect 293218 258680 293224 258692
rect 293276 258680 293282 258732
rect 191742 258476 191748 258528
rect 191800 258516 191806 258528
rect 197354 258516 197360 258528
rect 191800 258488 197360 258516
rect 191800 258476 191806 258488
rect 197354 258476 197360 258488
rect 197412 258476 197418 258528
rect 56318 258136 56324 258188
rect 56376 258176 56382 258188
rect 66346 258176 66352 258188
rect 56376 258148 66352 258176
rect 56376 258136 56382 258148
rect 66346 258136 66352 258148
rect 66404 258136 66410 258188
rect 43898 258068 43904 258120
rect 43956 258108 43962 258120
rect 66806 258108 66812 258120
rect 43956 258080 66812 258108
rect 43956 258068 43962 258080
rect 66806 258068 66812 258080
rect 66864 258068 66870 258120
rect 156598 258068 156604 258120
rect 156656 258108 156662 258120
rect 162118 258108 162124 258120
rect 156656 258080 162124 258108
rect 156656 258068 156662 258080
rect 162118 258068 162124 258080
rect 162176 258068 162182 258120
rect 189718 258068 189724 258120
rect 189776 258108 189782 258120
rect 191742 258108 191748 258120
rect 189776 258080 191748 258108
rect 189776 258068 189782 258080
rect 191742 258068 191748 258080
rect 191800 258068 191806 258120
rect 66346 258000 66352 258052
rect 66404 258040 66410 258052
rect 68094 258040 68100 258052
rect 66404 258012 68100 258040
rect 66404 258000 66410 258012
rect 68094 258000 68100 258012
rect 68152 258000 68158 258052
rect 157242 257932 157248 257984
rect 157300 257972 157306 257984
rect 162486 257972 162492 257984
rect 157300 257944 162492 257972
rect 157300 257932 157306 257944
rect 162486 257932 162492 257944
rect 162544 257932 162550 257984
rect 247218 257320 247224 257372
rect 247276 257360 247282 257372
rect 322934 257360 322940 257372
rect 247276 257332 322940 257360
rect 247276 257320 247282 257332
rect 322934 257320 322940 257332
rect 322992 257320 322998 257372
rect 61838 256708 61844 256760
rect 61896 256748 61902 256760
rect 66438 256748 66444 256760
rect 61896 256720 66444 256748
rect 61896 256708 61902 256720
rect 66438 256708 66444 256720
rect 66496 256708 66502 256760
rect 157242 256708 157248 256760
rect 157300 256748 157306 256760
rect 171042 256748 171048 256760
rect 157300 256720 171048 256748
rect 157300 256708 157306 256720
rect 171042 256708 171048 256720
rect 171100 256748 171106 256760
rect 173434 256748 173440 256760
rect 171100 256720 173440 256748
rect 171100 256708 171106 256720
rect 173434 256708 173440 256720
rect 173492 256708 173498 256760
rect 175826 256708 175832 256760
rect 175884 256748 175890 256760
rect 183462 256748 183468 256760
rect 175884 256720 183468 256748
rect 175884 256708 175890 256720
rect 183462 256708 183468 256720
rect 183520 256748 183526 256760
rect 197354 256748 197360 256760
rect 183520 256720 197360 256748
rect 183520 256708 183526 256720
rect 197354 256708 197360 256720
rect 197412 256708 197418 256760
rect 178770 256028 178776 256080
rect 178828 256068 178834 256080
rect 183002 256068 183008 256080
rect 178828 256040 183008 256068
rect 178828 256028 178834 256040
rect 183002 256028 183008 256040
rect 183060 256028 183066 256080
rect 159634 255960 159640 256012
rect 159692 256000 159698 256012
rect 181622 256000 181628 256012
rect 159692 255972 181628 256000
rect 159692 255960 159698 255972
rect 181622 255960 181628 255972
rect 181680 255960 181686 256012
rect 157242 255280 157248 255332
rect 157300 255320 157306 255332
rect 165522 255320 165528 255332
rect 157300 255292 165528 255320
rect 157300 255280 157306 255292
rect 165522 255280 165528 255292
rect 165580 255280 165586 255332
rect 187234 255280 187240 255332
rect 187292 255320 187298 255332
rect 197354 255320 197360 255332
rect 187292 255292 197360 255320
rect 187292 255280 187298 255292
rect 197354 255280 197360 255292
rect 197412 255280 197418 255332
rect 3418 255212 3424 255264
rect 3476 255252 3482 255264
rect 14458 255252 14464 255264
rect 3476 255224 14464 255252
rect 3476 255212 3482 255224
rect 14458 255212 14464 255224
rect 14516 255212 14522 255264
rect 157242 254532 157248 254584
rect 157300 254572 157306 254584
rect 189718 254572 189724 254584
rect 157300 254544 189724 254572
rect 157300 254532 157306 254544
rect 189718 254532 189724 254544
rect 189776 254532 189782 254584
rect 254026 254532 254032 254584
rect 254084 254572 254090 254584
rect 305086 254572 305092 254584
rect 254084 254544 305092 254572
rect 254084 254532 254090 254544
rect 305086 254532 305092 254544
rect 305144 254532 305150 254584
rect 52270 253920 52276 253972
rect 52328 253960 52334 253972
rect 66438 253960 66444 253972
rect 52328 253932 66444 253960
rect 52328 253920 52334 253932
rect 66438 253920 66444 253932
rect 66496 253920 66502 253972
rect 188522 253920 188528 253972
rect 188580 253960 188586 253972
rect 197354 253960 197360 253972
rect 188580 253932 197360 253960
rect 188580 253920 188586 253932
rect 197354 253920 197360 253932
rect 197412 253920 197418 253972
rect 246022 253920 246028 253972
rect 246080 253960 246086 253972
rect 249978 253960 249984 253972
rect 246080 253932 249984 253960
rect 246080 253920 246086 253932
rect 249978 253920 249984 253932
rect 250036 253920 250042 253972
rect 157242 253852 157248 253904
rect 157300 253892 157306 253904
rect 175826 253892 175832 253904
rect 157300 253864 175832 253892
rect 157300 253852 157306 253864
rect 175826 253852 175832 253864
rect 175884 253852 175890 253904
rect 194502 253852 194508 253904
rect 194560 253892 194566 253904
rect 197446 253892 197452 253904
rect 194560 253864 197452 253892
rect 194560 253852 194566 253864
rect 197446 253852 197452 253864
rect 197504 253852 197510 253904
rect 245930 253852 245936 253904
rect 245988 253892 245994 253904
rect 256694 253892 256700 253904
rect 245988 253864 256700 253892
rect 245988 253852 245994 253864
rect 256694 253852 256700 253864
rect 256752 253892 256758 253904
rect 256878 253892 256884 253904
rect 256752 253864 256884 253892
rect 256752 253852 256758 253864
rect 256878 253852 256884 253864
rect 256936 253852 256942 253904
rect 167638 253172 167644 253224
rect 167696 253212 167702 253224
rect 177390 253212 177396 253224
rect 167696 253184 177396 253212
rect 167696 253172 167702 253184
rect 177390 253172 177396 253184
rect 177448 253172 177454 253224
rect 256878 253172 256884 253224
rect 256936 253212 256942 253224
rect 327258 253212 327264 253224
rect 256936 253184 327264 253212
rect 256936 253172 256942 253184
rect 327258 253172 327264 253184
rect 327316 253172 327322 253224
rect 245930 252832 245936 252884
rect 245988 252872 245994 252884
rect 248506 252872 248512 252884
rect 245988 252844 248512 252872
rect 245988 252832 245994 252844
rect 248506 252832 248512 252844
rect 248564 252872 248570 252884
rect 249058 252872 249064 252884
rect 248564 252844 249064 252872
rect 248564 252832 248570 252844
rect 249058 252832 249064 252844
rect 249116 252832 249122 252884
rect 59170 252628 59176 252680
rect 59228 252668 59234 252680
rect 64598 252668 64604 252680
rect 59228 252640 64604 252668
rect 59228 252628 59234 252640
rect 64598 252628 64604 252640
rect 64656 252668 64662 252680
rect 66622 252668 66628 252680
rect 64656 252640 66628 252668
rect 64656 252628 64662 252640
rect 66622 252628 66628 252640
rect 66680 252628 66686 252680
rect 245746 252424 245752 252476
rect 245804 252464 245810 252476
rect 255314 252464 255320 252476
rect 245804 252436 255320 252464
rect 245804 252424 245810 252436
rect 255314 252424 255320 252436
rect 255372 252424 255378 252476
rect 165522 251812 165528 251864
rect 165580 251852 165586 251864
rect 184842 251852 184848 251864
rect 165580 251824 184848 251852
rect 165580 251812 165586 251824
rect 184842 251812 184848 251824
rect 184900 251812 184906 251864
rect 255314 251812 255320 251864
rect 255372 251852 255378 251864
rect 522298 251852 522304 251864
rect 255372 251824 522304 251852
rect 255372 251812 255378 251824
rect 522298 251812 522304 251824
rect 522356 251812 522362 251864
rect 192570 251268 192576 251320
rect 192628 251308 192634 251320
rect 197446 251308 197452 251320
rect 192628 251280 197452 251308
rect 192628 251268 192634 251280
rect 197446 251268 197452 251280
rect 197504 251268 197510 251320
rect 157242 251200 157248 251252
rect 157300 251240 157306 251252
rect 168374 251240 168380 251252
rect 157300 251212 168380 251240
rect 157300 251200 157306 251212
rect 168374 251200 168380 251212
rect 168432 251200 168438 251252
rect 184842 251200 184848 251252
rect 184900 251240 184906 251252
rect 197354 251240 197360 251252
rect 184900 251212 197360 251240
rect 184900 251200 184906 251212
rect 197354 251200 197360 251212
rect 197412 251200 197418 251252
rect 156138 250452 156144 250504
rect 156196 250492 156202 250504
rect 174722 250492 174728 250504
rect 156196 250464 174728 250492
rect 156196 250452 156202 250464
rect 174722 250452 174728 250464
rect 174780 250452 174786 250504
rect 287698 250452 287704 250504
rect 287756 250492 287762 250504
rect 317506 250492 317512 250504
rect 287756 250464 317512 250492
rect 287756 250452 287762 250464
rect 317506 250452 317512 250464
rect 317564 250452 317570 250504
rect 195330 249908 195336 249960
rect 195388 249948 195394 249960
rect 197446 249948 197452 249960
rect 195388 249920 197452 249948
rect 195388 249908 195394 249920
rect 197446 249908 197452 249920
rect 197504 249908 197510 249960
rect 157242 249772 157248 249824
rect 157300 249812 157306 249824
rect 176102 249812 176108 249824
rect 157300 249784 176108 249812
rect 157300 249772 157306 249784
rect 176102 249772 176108 249784
rect 176160 249772 176166 249824
rect 178954 249772 178960 249824
rect 179012 249812 179018 249824
rect 197354 249812 197360 249824
rect 179012 249784 197360 249812
rect 179012 249772 179018 249784
rect 197354 249772 197360 249784
rect 197412 249772 197418 249824
rect 245746 249772 245752 249824
rect 245804 249812 245810 249824
rect 255314 249812 255320 249824
rect 245804 249784 255320 249812
rect 245804 249772 245810 249784
rect 255314 249772 255320 249784
rect 255372 249772 255378 249824
rect 192478 249704 192484 249756
rect 192536 249744 192542 249756
rect 193030 249744 193036 249756
rect 192536 249716 193036 249744
rect 192536 249704 192542 249716
rect 193030 249704 193036 249716
rect 193088 249744 193094 249756
rect 197446 249744 197452 249756
rect 193088 249716 197452 249744
rect 193088 249704 193094 249716
rect 197446 249704 197452 249716
rect 197504 249704 197510 249756
rect 245930 249500 245936 249552
rect 245988 249540 245994 249552
rect 249794 249540 249800 249552
rect 245988 249512 249800 249540
rect 245988 249500 245994 249512
rect 249794 249500 249800 249512
rect 249852 249500 249858 249552
rect 157242 249432 157248 249484
rect 157300 249472 157306 249484
rect 163682 249472 163688 249484
rect 157300 249444 163688 249472
rect 157300 249432 157306 249444
rect 163682 249432 163688 249444
rect 163740 249432 163746 249484
rect 181990 249024 181996 249076
rect 182048 249064 182054 249076
rect 195330 249064 195336 249076
rect 182048 249036 195336 249064
rect 182048 249024 182054 249036
rect 195330 249024 195336 249036
rect 195388 249024 195394 249076
rect 268378 249024 268384 249076
rect 268436 249064 268442 249076
rect 334066 249064 334072 249076
rect 268436 249036 334072 249064
rect 268436 249024 268442 249036
rect 334066 249024 334072 249036
rect 334124 249024 334130 249076
rect 173158 248888 173164 248940
rect 173216 248928 173222 248940
rect 178862 248928 178868 248940
rect 173216 248900 178868 248928
rect 173216 248888 173222 248900
rect 178862 248888 178868 248900
rect 178920 248888 178926 248940
rect 62022 248412 62028 248464
rect 62080 248452 62086 248464
rect 66806 248452 66812 248464
rect 62080 248424 66812 248452
rect 62080 248412 62086 248424
rect 66806 248412 66812 248424
rect 66864 248412 66870 248464
rect 157150 248412 157156 248464
rect 157208 248452 157214 248464
rect 174170 248452 174176 248464
rect 157208 248424 174176 248452
rect 157208 248412 157214 248424
rect 174170 248412 174176 248424
rect 174228 248412 174234 248464
rect 157242 247732 157248 247784
rect 157300 247772 157306 247784
rect 165522 247772 165528 247784
rect 157300 247744 165528 247772
rect 157300 247732 157306 247744
rect 165522 247732 165528 247744
rect 165580 247732 165586 247784
rect 169202 247732 169208 247784
rect 169260 247772 169266 247784
rect 191282 247772 191288 247784
rect 169260 247744 191288 247772
rect 169260 247732 169266 247744
rect 191282 247732 191288 247744
rect 191340 247732 191346 247784
rect 158070 247664 158076 247716
rect 158128 247704 158134 247716
rect 192570 247704 192576 247716
rect 158128 247676 192576 247704
rect 158128 247664 158134 247676
rect 192570 247664 192576 247676
rect 192628 247664 192634 247716
rect 245930 247664 245936 247716
rect 245988 247704 245994 247716
rect 246114 247704 246120 247716
rect 245988 247676 246120 247704
rect 245988 247664 245994 247676
rect 246114 247664 246120 247676
rect 246172 247704 246178 247716
rect 583294 247704 583300 247716
rect 246172 247676 583300 247704
rect 246172 247664 246178 247676
rect 583294 247664 583300 247676
rect 583352 247664 583358 247716
rect 59170 247052 59176 247104
rect 59228 247092 59234 247104
rect 66806 247092 66812 247104
rect 59228 247064 66812 247092
rect 59228 247052 59234 247064
rect 66806 247052 66812 247064
rect 66864 247052 66870 247104
rect 166350 247052 166356 247104
rect 166408 247092 166414 247104
rect 167730 247092 167736 247104
rect 166408 247064 167736 247092
rect 166408 247052 166414 247064
rect 167730 247052 167736 247064
rect 167788 247052 167794 247104
rect 194134 247052 194140 247104
rect 194192 247092 194198 247104
rect 197354 247092 197360 247104
rect 194192 247064 197360 247092
rect 194192 247052 194198 247064
rect 197354 247052 197360 247064
rect 197412 247052 197418 247104
rect 191098 246984 191104 247036
rect 191156 247024 191162 247036
rect 197446 247024 197452 247036
rect 191156 246996 197452 247024
rect 191156 246984 191162 246996
rect 197446 246984 197452 246996
rect 197504 246984 197510 247036
rect 244918 246304 244924 246356
rect 244976 246344 244982 246356
rect 269114 246344 269120 246356
rect 244976 246316 269120 246344
rect 244976 246304 244982 246316
rect 269114 246304 269120 246316
rect 269172 246304 269178 246356
rect 166534 245692 166540 245744
rect 166592 245732 166598 245744
rect 188982 245732 188988 245744
rect 166592 245704 188988 245732
rect 166592 245692 166598 245704
rect 188982 245692 188988 245704
rect 189040 245732 189046 245744
rect 197354 245732 197360 245744
rect 189040 245704 197360 245732
rect 189040 245692 189046 245704
rect 197354 245692 197360 245704
rect 197412 245692 197418 245744
rect 157242 245624 157248 245676
rect 157300 245664 157306 245676
rect 180058 245664 180064 245676
rect 157300 245636 180064 245664
rect 157300 245624 157306 245636
rect 180058 245624 180064 245636
rect 180116 245624 180122 245676
rect 246390 245624 246396 245676
rect 246448 245664 246454 245676
rect 247034 245664 247040 245676
rect 246448 245636 247040 245664
rect 246448 245624 246454 245636
rect 247034 245624 247040 245636
rect 247092 245664 247098 245676
rect 302234 245664 302240 245676
rect 247092 245636 302240 245664
rect 247092 245624 247098 245636
rect 302234 245624 302240 245636
rect 302292 245624 302298 245676
rect 57698 244876 57704 244928
rect 57756 244916 57762 244928
rect 67174 244916 67180 244928
rect 57756 244888 67180 244916
rect 57756 244876 57762 244888
rect 67174 244876 67180 244888
rect 67232 244876 67238 244928
rect 280798 244876 280804 244928
rect 280856 244916 280862 244928
rect 310514 244916 310520 244928
rect 280856 244888 310520 244916
rect 280856 244876 280862 244888
rect 310514 244876 310520 244888
rect 310572 244876 310578 244928
rect 188430 244332 188436 244384
rect 188488 244372 188494 244384
rect 188488 244344 189764 244372
rect 188488 244332 188494 244344
rect 157978 244264 157984 244316
rect 158036 244304 158042 244316
rect 189074 244304 189080 244316
rect 158036 244276 189080 244304
rect 158036 244264 158042 244276
rect 189074 244264 189080 244276
rect 189132 244264 189138 244316
rect 189736 244304 189764 244344
rect 189902 244332 189908 244384
rect 189960 244372 189966 244384
rect 191650 244372 191656 244384
rect 189960 244344 191656 244372
rect 189960 244332 189966 244344
rect 191650 244332 191656 244344
rect 191708 244372 191714 244384
rect 197446 244372 197452 244384
rect 191708 244344 197452 244372
rect 191708 244332 191714 244344
rect 197446 244332 197452 244344
rect 197504 244332 197510 244384
rect 190362 244304 190368 244316
rect 189736 244276 190368 244304
rect 190362 244264 190368 244276
rect 190420 244304 190426 244316
rect 197354 244304 197360 244316
rect 190420 244276 197360 244304
rect 190420 244264 190426 244276
rect 197354 244264 197360 244276
rect 197412 244264 197418 244316
rect 245930 244264 245936 244316
rect 245988 244304 245994 244316
rect 258074 244304 258080 244316
rect 245988 244276 258080 244304
rect 245988 244264 245994 244276
rect 258074 244264 258080 244276
rect 258132 244264 258138 244316
rect 174170 243516 174176 243568
rect 174228 243556 174234 243568
rect 199562 243556 199568 243568
rect 174228 243528 199568 243556
rect 174228 243516 174234 243528
rect 199562 243516 199568 243528
rect 199620 243516 199626 243568
rect 286410 243516 286416 243568
rect 286468 243556 286474 243568
rect 321646 243556 321652 243568
rect 286468 243528 321652 243556
rect 286468 243516 286474 243528
rect 321646 243516 321652 243528
rect 321704 243516 321710 243568
rect 156138 242972 156144 243024
rect 156196 243012 156202 243024
rect 158070 243012 158076 243024
rect 156196 242984 158076 243012
rect 156196 242972 156202 242984
rect 158070 242972 158076 242984
rect 158128 242972 158134 243024
rect 157242 242904 157248 242956
rect 157300 242944 157306 242956
rect 189902 242944 189908 242956
rect 157300 242916 189908 242944
rect 157300 242904 157306 242916
rect 189902 242904 189908 242916
rect 189960 242904 189966 242956
rect 246390 242904 246396 242956
rect 246448 242944 246454 242956
rect 247218 242944 247224 242956
rect 246448 242916 247224 242944
rect 246448 242904 246454 242916
rect 247218 242904 247224 242916
rect 247276 242944 247282 242956
rect 286502 242944 286508 242956
rect 247276 242916 286508 242944
rect 247276 242904 247282 242916
rect 286502 242904 286508 242916
rect 286560 242904 286566 242956
rect 166442 242156 166448 242208
rect 166500 242196 166506 242208
rect 184382 242196 184388 242208
rect 166500 242168 184388 242196
rect 166500 242156 166506 242168
rect 184382 242156 184388 242168
rect 184440 242156 184446 242208
rect 244274 242156 244280 242208
rect 244332 242196 244338 242208
rect 329926 242196 329932 242208
rect 244332 242168 329932 242196
rect 244332 242156 244338 242168
rect 329926 242156 329932 242168
rect 329984 242156 329990 242208
rect 65978 242020 65984 242072
rect 66036 242060 66042 242072
rect 71038 242060 71044 242072
rect 66036 242032 71044 242060
rect 66036 242020 66042 242032
rect 71038 242020 71044 242032
rect 71096 242020 71102 242072
rect 152458 242020 152464 242072
rect 152516 242060 152522 242072
rect 155218 242060 155224 242072
rect 152516 242032 155224 242060
rect 152516 242020 152522 242032
rect 155218 242020 155224 242032
rect 155276 242020 155282 242072
rect 69750 241816 69756 241868
rect 69808 241856 69814 241868
rect 72418 241856 72424 241868
rect 69808 241828 72424 241856
rect 69808 241816 69814 241828
rect 72418 241816 72424 241828
rect 72476 241816 72482 241868
rect 153838 241476 153844 241528
rect 153896 241516 153902 241528
rect 192938 241516 192944 241528
rect 153896 241488 192944 241516
rect 153896 241476 153902 241488
rect 192938 241476 192944 241488
rect 192996 241476 193002 241528
rect 195790 241476 195796 241528
rect 195848 241516 195854 241528
rect 197906 241516 197912 241528
rect 195848 241488 197912 241516
rect 195848 241476 195854 241488
rect 197906 241476 197912 241488
rect 197964 241476 197970 241528
rect 246298 241476 246304 241528
rect 246356 241516 246362 241528
rect 247126 241516 247132 241528
rect 246356 241488 247132 241516
rect 246356 241476 246362 241488
rect 247126 241476 247132 241488
rect 247184 241516 247190 241528
rect 320266 241516 320272 241528
rect 247184 241488 320272 241516
rect 247184 241476 247190 241488
rect 320266 241476 320272 241488
rect 320324 241476 320330 241528
rect 3418 241408 3424 241460
rect 3476 241448 3482 241460
rect 32398 241448 32404 241460
rect 3476 241420 32404 241448
rect 3476 241408 3482 241420
rect 32398 241408 32404 241420
rect 32456 241408 32462 241460
rect 105032 241408 105038 241460
rect 105090 241448 105096 241460
rect 155402 241448 155408 241460
rect 105090 241420 155408 241448
rect 105090 241408 105096 241420
rect 155402 241408 155408 241420
rect 155460 241408 155466 241460
rect 67450 240796 67456 240848
rect 67508 240836 67514 240848
rect 81250 240836 81256 240848
rect 67508 240808 81256 240836
rect 67508 240796 67514 240808
rect 81250 240796 81256 240808
rect 81308 240796 81314 240848
rect 258718 240796 258724 240848
rect 258776 240836 258782 240848
rect 278038 240836 278044 240848
rect 258776 240808 278044 240836
rect 258776 240796 258782 240808
rect 278038 240796 278044 240808
rect 278096 240796 278102 240848
rect 64506 240728 64512 240780
rect 64564 240768 64570 240780
rect 103606 240768 103612 240780
rect 64564 240740 103612 240768
rect 64564 240728 64570 240740
rect 103606 240728 103612 240740
rect 103664 240728 103670 240780
rect 120994 240728 121000 240780
rect 121052 240768 121058 240780
rect 200114 240768 200120 240780
rect 121052 240740 200120 240768
rect 121052 240728 121058 240740
rect 200114 240728 200120 240740
rect 200172 240728 200178 240780
rect 244090 240728 244096 240780
rect 244148 240768 244154 240780
rect 580258 240768 580264 240780
rect 244148 240740 580264 240768
rect 244148 240728 244154 240740
rect 580258 240728 580264 240740
rect 580316 240728 580322 240780
rect 199930 240456 199936 240508
rect 199988 240496 199994 240508
rect 199988 240468 201172 240496
rect 199988 240456 199994 240468
rect 196618 240388 196624 240440
rect 196676 240428 196682 240440
rect 196676 240400 201080 240428
rect 196676 240388 196682 240400
rect 200114 240320 200120 240372
rect 200172 240360 200178 240372
rect 200172 240332 200344 240360
rect 200172 240320 200178 240332
rect 200316 240168 200344 240332
rect 201052 240168 201080 240400
rect 200298 240116 200304 240168
rect 200356 240116 200362 240168
rect 201034 240116 201040 240168
rect 201092 240116 201098 240168
rect 201144 240156 201172 240468
rect 201402 240156 201408 240168
rect 201144 240128 201408 240156
rect 201402 240116 201408 240128
rect 201460 240116 201466 240168
rect 231946 240116 231952 240168
rect 232004 240156 232010 240168
rect 235810 240156 235816 240168
rect 232004 240128 235816 240156
rect 232004 240116 232010 240128
rect 235810 240116 235816 240128
rect 235868 240116 235874 240168
rect 245746 240116 245752 240168
rect 245804 240156 245810 240168
rect 256694 240156 256700 240168
rect 245804 240128 256700 240156
rect 245804 240116 245810 240128
rect 256694 240116 256700 240128
rect 256752 240116 256758 240168
rect 86034 240048 86040 240100
rect 86092 240088 86098 240100
rect 86862 240088 86868 240100
rect 86092 240060 86868 240088
rect 86092 240048 86098 240060
rect 86862 240048 86868 240060
rect 86920 240048 86926 240100
rect 91922 240048 91928 240100
rect 91980 240088 91986 240100
rect 92382 240088 92388 240100
rect 91980 240060 92388 240088
rect 91980 240048 91986 240060
rect 92382 240048 92388 240060
rect 92440 240048 92446 240100
rect 101122 240048 101128 240100
rect 101180 240088 101186 240100
rect 101950 240088 101956 240100
rect 101180 240060 101956 240088
rect 101180 240048 101186 240060
rect 101950 240048 101956 240060
rect 102008 240048 102014 240100
rect 115290 240048 115296 240100
rect 115348 240088 115354 240100
rect 115842 240088 115848 240100
rect 115348 240060 115848 240088
rect 115348 240048 115354 240060
rect 115842 240048 115848 240060
rect 115900 240048 115906 240100
rect 118786 240048 118792 240100
rect 118844 240088 118850 240100
rect 119982 240088 119988 240100
rect 118844 240060 119988 240088
rect 118844 240048 118850 240060
rect 119982 240048 119988 240060
rect 120040 240048 120046 240100
rect 121730 240048 121736 240100
rect 121788 240088 121794 240100
rect 122742 240088 122748 240100
rect 121788 240060 122748 240088
rect 121788 240048 121794 240060
rect 122742 240048 122748 240060
rect 122800 240048 122806 240100
rect 124674 240048 124680 240100
rect 124732 240088 124738 240100
rect 125502 240088 125508 240100
rect 124732 240060 125508 240088
rect 124732 240048 124738 240060
rect 125502 240048 125508 240060
rect 125560 240048 125566 240100
rect 128906 240048 128912 240100
rect 128964 240088 128970 240100
rect 129642 240088 129648 240100
rect 128964 240060 129648 240088
rect 128964 240048 128970 240060
rect 129642 240048 129648 240060
rect 129700 240048 129706 240100
rect 130378 240048 130384 240100
rect 130436 240088 130442 240100
rect 130930 240088 130936 240100
rect 130436 240060 130936 240088
rect 130436 240048 130442 240060
rect 130930 240048 130936 240060
rect 130988 240048 130994 240100
rect 249702 240048 249708 240100
rect 249760 240088 249766 240100
rect 250070 240088 250076 240100
rect 249760 240060 250076 240088
rect 249760 240048 249766 240060
rect 250070 240048 250076 240060
rect 250128 240048 250134 240100
rect 96890 239980 96896 240032
rect 96948 240020 96954 240032
rect 101490 240020 101496 240032
rect 96948 239992 101496 240020
rect 96948 239980 96954 239992
rect 101490 239980 101496 239992
rect 101548 239980 101554 240032
rect 114646 239980 114652 240032
rect 114704 240020 114710 240032
rect 115382 240020 115388 240032
rect 114704 239992 115388 240020
rect 114704 239980 114710 239992
rect 115382 239980 115388 239992
rect 115440 239980 115446 240032
rect 116762 239980 116768 240032
rect 116820 240020 116826 240032
rect 124306 240020 124312 240032
rect 116820 239992 124312 240020
rect 116820 239980 116826 239992
rect 124306 239980 124312 239992
rect 124364 239980 124370 240032
rect 75362 239912 75368 239964
rect 75420 239952 75426 239964
rect 75822 239952 75828 239964
rect 75420 239924 75828 239952
rect 75420 239912 75426 239924
rect 75822 239912 75828 239924
rect 75880 239912 75886 239964
rect 88978 239912 88984 239964
rect 89036 239952 89042 239964
rect 89530 239952 89536 239964
rect 89036 239924 89536 239952
rect 89036 239912 89042 239924
rect 89530 239912 89536 239924
rect 89588 239912 89594 239964
rect 90450 239912 90456 239964
rect 90508 239952 90514 239964
rect 90910 239952 90916 239964
rect 90508 239924 90916 239952
rect 90508 239912 90514 239924
rect 90910 239912 90916 239924
rect 90968 239912 90974 239964
rect 147766 239912 147772 239964
rect 147824 239952 147830 239964
rect 148318 239952 148324 239964
rect 147824 239924 148324 239952
rect 147824 239912 147830 239924
rect 148318 239912 148324 239924
rect 148376 239912 148382 239964
rect 106826 239776 106832 239828
rect 106884 239816 106890 239828
rect 107562 239816 107568 239828
rect 106884 239788 107568 239816
rect 106884 239776 106890 239788
rect 107562 239776 107568 239788
rect 107620 239776 107626 239828
rect 109586 239776 109592 239828
rect 109644 239816 109650 239828
rect 110322 239816 110328 239828
rect 109644 239788 110328 239816
rect 109644 239776 109650 239788
rect 110322 239776 110328 239788
rect 110380 239776 110386 239828
rect 68922 239504 68928 239556
rect 68980 239544 68986 239556
rect 70302 239544 70308 239556
rect 68980 239516 70308 239544
rect 68980 239504 68986 239516
rect 70302 239504 70308 239516
rect 70360 239504 70366 239556
rect 81526 239504 81532 239556
rect 81584 239544 81590 239556
rect 82722 239544 82728 239556
rect 81584 239516 82728 239544
rect 81584 239504 81590 239516
rect 82722 239504 82728 239516
rect 82780 239504 82786 239556
rect 99374 239504 99380 239556
rect 99432 239544 99438 239556
rect 100662 239544 100668 239556
rect 99432 239516 100668 239544
rect 99432 239504 99438 239516
rect 100662 239504 100668 239516
rect 100720 239504 100726 239556
rect 70210 239436 70216 239488
rect 70268 239476 70274 239488
rect 108298 239476 108304 239488
rect 70268 239448 108304 239476
rect 70268 239436 70274 239448
rect 108298 239436 108304 239448
rect 108356 239436 108362 239488
rect 110230 239436 110236 239488
rect 110288 239476 110294 239488
rect 115198 239476 115204 239488
rect 110288 239448 115204 239476
rect 110288 239436 110294 239448
rect 115198 239436 115204 239448
rect 115256 239436 115262 239488
rect 149698 239436 149704 239488
rect 149756 239476 149762 239488
rect 240318 239476 240324 239488
rect 149756 239448 240324 239476
rect 149756 239436 149762 239448
rect 240318 239436 240324 239448
rect 240376 239436 240382 239488
rect 79042 239368 79048 239420
rect 79100 239408 79106 239420
rect 79962 239408 79968 239420
rect 79100 239380 79968 239408
rect 79100 239368 79106 239380
rect 79962 239368 79968 239380
rect 80020 239368 80026 239420
rect 80514 239368 80520 239420
rect 80572 239408 80578 239420
rect 88978 239408 88984 239420
rect 80572 239380 88984 239408
rect 80572 239368 80578 239380
rect 88978 239368 88984 239380
rect 89036 239368 89042 239420
rect 108206 239368 108212 239420
rect 108264 239408 108270 239420
rect 208394 239408 208400 239420
rect 108264 239380 208400 239408
rect 108264 239368 108270 239380
rect 208394 239368 208400 239380
rect 208452 239368 208458 239420
rect 102594 239232 102600 239284
rect 102652 239272 102658 239284
rect 103330 239272 103336 239284
rect 102652 239244 103336 239272
rect 102652 239232 102658 239244
rect 103330 239232 103336 239244
rect 103388 239232 103394 239284
rect 107746 239232 107752 239284
rect 107804 239272 107810 239284
rect 108390 239272 108396 239284
rect 107804 239244 108396 239272
rect 107804 239232 107810 239244
rect 108390 239232 108396 239244
rect 108448 239232 108454 239284
rect 111058 239232 111064 239284
rect 111116 239272 111122 239284
rect 111702 239272 111708 239284
rect 111116 239244 111708 239272
rect 111116 239232 111122 239244
rect 111702 239232 111708 239244
rect 111760 239232 111766 239284
rect 131850 239232 131856 239284
rect 131908 239272 131914 239284
rect 132310 239272 132316 239284
rect 131908 239244 132316 239272
rect 131908 239232 131914 239244
rect 132310 239232 132316 239244
rect 132368 239232 132374 239284
rect 143994 239232 144000 239284
rect 144052 239272 144058 239284
rect 144730 239272 144736 239284
rect 144052 239244 144736 239272
rect 144052 239232 144058 239244
rect 144730 239232 144736 239244
rect 144788 239232 144794 239284
rect 153930 239232 153936 239284
rect 153988 239272 153994 239284
rect 154482 239272 154488 239284
rect 153988 239244 154488 239272
rect 153988 239232 153994 239244
rect 154482 239232 154488 239244
rect 154540 239232 154546 239284
rect 145282 239096 145288 239148
rect 145340 239136 145346 239148
rect 145926 239136 145932 239148
rect 145340 239108 145932 239136
rect 145340 239096 145346 239108
rect 145926 239096 145932 239108
rect 145984 239096 145990 239148
rect 148226 239096 148232 239148
rect 148284 239136 148290 239148
rect 148962 239136 148968 239148
rect 148284 239108 148968 239136
rect 148284 239096 148290 239108
rect 148962 239096 148968 239108
rect 149020 239096 149026 239148
rect 133138 238960 133144 239012
rect 133196 239000 133202 239012
rect 133690 239000 133696 239012
rect 133196 238972 133696 239000
rect 133196 238960 133202 238972
rect 133690 238960 133696 238972
rect 133748 238960 133754 239012
rect 134610 238960 134616 239012
rect 134668 239000 134674 239012
rect 135162 239000 135168 239012
rect 134668 238972 135168 239000
rect 134668 238960 134674 238972
rect 135162 238960 135168 238972
rect 135220 238960 135226 239012
rect 74442 238756 74448 238808
rect 74500 238796 74506 238808
rect 75454 238796 75460 238808
rect 74500 238768 75460 238796
rect 74500 238756 74506 238768
rect 75454 238756 75460 238768
rect 75512 238756 75518 238808
rect 83090 238688 83096 238740
rect 83148 238728 83154 238740
rect 207658 238728 207664 238740
rect 83148 238700 207664 238728
rect 83148 238688 83154 238700
rect 207658 238688 207664 238700
rect 207716 238688 207722 238740
rect 208394 238688 208400 238740
rect 208452 238728 208458 238740
rect 219894 238728 219900 238740
rect 208452 238700 219900 238728
rect 208452 238688 208458 238700
rect 219894 238688 219900 238700
rect 219952 238688 219958 238740
rect 220814 238688 220820 238740
rect 220872 238728 220878 238740
rect 222286 238728 222292 238740
rect 220872 238700 222292 238728
rect 220872 238688 220878 238700
rect 222286 238688 222292 238700
rect 222344 238688 222350 238740
rect 101490 238620 101496 238672
rect 101548 238660 101554 238672
rect 214190 238660 214196 238672
rect 101548 238632 214196 238660
rect 101548 238620 101554 238632
rect 214190 238620 214196 238632
rect 214248 238620 214254 238672
rect 216582 238348 216588 238400
rect 216640 238388 216646 238400
rect 218054 238388 218060 238400
rect 216640 238360 218060 238388
rect 216640 238348 216646 238360
rect 218054 238348 218060 238360
rect 218112 238348 218118 238400
rect 67910 238076 67916 238128
rect 67968 238116 67974 238128
rect 79318 238116 79324 238128
rect 67968 238088 79324 238116
rect 67968 238076 67974 238088
rect 79318 238076 79324 238088
rect 79376 238076 79382 238128
rect 224770 238076 224776 238128
rect 224828 238116 224834 238128
rect 226702 238116 226708 238128
rect 224828 238088 226708 238116
rect 224828 238076 224834 238088
rect 226702 238076 226708 238088
rect 226760 238076 226766 238128
rect 67358 238008 67364 238060
rect 67416 238048 67422 238060
rect 98546 238048 98552 238060
rect 67416 238020 98552 238048
rect 67416 238008 67422 238020
rect 98546 238008 98552 238020
rect 98604 238008 98610 238060
rect 226978 238008 226984 238060
rect 227036 238048 227042 238060
rect 238846 238048 238852 238060
rect 227036 238020 238852 238048
rect 227036 238008 227042 238020
rect 238846 238008 238852 238020
rect 238904 238008 238910 238060
rect 240318 238008 240324 238060
rect 240376 238048 240382 238060
rect 301498 238048 301504 238060
rect 240376 238020 301504 238048
rect 240376 238008 240382 238020
rect 301498 238008 301504 238020
rect 301556 238008 301562 238060
rect 218146 237464 218152 237516
rect 218204 237504 218210 237516
rect 218698 237504 218704 237516
rect 218204 237476 218704 237504
rect 218204 237464 218210 237476
rect 218698 237464 218704 237476
rect 218756 237504 218762 237516
rect 218756 237476 219434 237504
rect 218756 237464 218762 237476
rect 219406 237436 219434 237476
rect 220078 237464 220084 237516
rect 220136 237504 220142 237516
rect 221918 237504 221924 237516
rect 220136 237476 221924 237504
rect 220136 237464 220142 237476
rect 221918 237464 221924 237476
rect 221976 237464 221982 237516
rect 222286 237464 222292 237516
rect 222344 237504 222350 237516
rect 222838 237504 222844 237516
rect 222344 237476 222844 237504
rect 222344 237464 222350 237476
rect 222838 237464 222844 237476
rect 222896 237464 222902 237516
rect 222930 237464 222936 237516
rect 222988 237504 222994 237516
rect 223758 237504 223764 237516
rect 222988 237476 223764 237504
rect 222988 237464 222994 237476
rect 223758 237464 223764 237476
rect 223816 237464 223822 237516
rect 233878 237436 233884 237448
rect 219406 237408 233884 237436
rect 233878 237396 233884 237408
rect 233936 237396 233942 237448
rect 237374 237396 237380 237448
rect 237432 237436 237438 237448
rect 240778 237436 240784 237448
rect 237432 237408 240784 237436
rect 237432 237396 237438 237408
rect 240778 237396 240784 237408
rect 240836 237396 240842 237448
rect 243262 237396 243268 237448
rect 243320 237436 243326 237448
rect 244274 237436 244280 237448
rect 243320 237408 244280 237436
rect 243320 237396 243326 237408
rect 244274 237396 244280 237408
rect 244332 237396 244338 237448
rect 4798 237328 4804 237380
rect 4856 237368 4862 237380
rect 54846 237368 54852 237380
rect 4856 237340 54852 237368
rect 4856 237328 4862 237340
rect 54846 237328 54852 237340
rect 54904 237368 54910 237380
rect 136634 237368 136640 237380
rect 54904 237340 136640 237368
rect 54904 237328 54910 237340
rect 136634 237328 136640 237340
rect 136692 237328 136698 237380
rect 138106 237328 138112 237380
rect 138164 237368 138170 237380
rect 160922 237368 160928 237380
rect 138164 237340 160928 237368
rect 138164 237328 138170 237340
rect 160922 237328 160928 237340
rect 160980 237328 160986 237380
rect 189718 237328 189724 237380
rect 189776 237368 189782 237380
rect 242710 237368 242716 237380
rect 189776 237340 242716 237368
rect 189776 237328 189782 237340
rect 242710 237328 242716 237340
rect 242768 237328 242774 237380
rect 81250 236648 81256 236700
rect 81308 236688 81314 236700
rect 248322 236688 248328 236700
rect 81308 236660 248328 236688
rect 81308 236648 81314 236660
rect 248322 236648 248328 236660
rect 248380 236648 248386 236700
rect 136634 235968 136640 236020
rect 136692 236008 136698 236020
rect 137278 236008 137284 236020
rect 136692 235980 137284 236008
rect 136692 235968 136698 235980
rect 137278 235968 137284 235980
rect 137336 235968 137342 236020
rect 103606 235900 103612 235952
rect 103664 235940 103670 235952
rect 180242 235940 180248 235952
rect 103664 235912 180248 235940
rect 103664 235900 103670 235912
rect 180242 235900 180248 235912
rect 180300 235900 180306 235952
rect 199562 235900 199568 235952
rect 199620 235940 199626 235952
rect 243630 235940 243636 235952
rect 199620 235912 243636 235940
rect 199620 235900 199626 235912
rect 243630 235900 243636 235912
rect 243688 235900 243694 235952
rect 146018 235424 146024 235476
rect 146076 235464 146082 235476
rect 153838 235464 153844 235476
rect 146076 235436 153844 235464
rect 146076 235424 146082 235436
rect 153838 235424 153844 235436
rect 153896 235424 153902 235476
rect 61930 235288 61936 235340
rect 61988 235328 61994 235340
rect 75178 235328 75184 235340
rect 61988 235300 75184 235328
rect 61988 235288 61994 235300
rect 75178 235288 75184 235300
rect 75236 235288 75242 235340
rect 61746 235220 61752 235272
rect 61804 235260 61810 235272
rect 124582 235260 124588 235272
rect 61804 235232 124588 235260
rect 61804 235220 61810 235232
rect 124582 235220 124588 235232
rect 124640 235220 124646 235272
rect 126790 235220 126796 235272
rect 126848 235260 126854 235272
rect 135254 235260 135260 235272
rect 126848 235232 135260 235260
rect 126848 235220 126854 235232
rect 135254 235220 135260 235232
rect 135312 235220 135318 235272
rect 176102 235220 176108 235272
rect 176160 235260 176166 235272
rect 198734 235260 198740 235272
rect 176160 235232 198740 235260
rect 176160 235220 176166 235232
rect 198734 235220 198740 235232
rect 198792 235220 198798 235272
rect 243630 235220 243636 235272
rect 243688 235260 243694 235272
rect 260098 235260 260104 235272
rect 243688 235232 260104 235260
rect 243688 235220 243694 235232
rect 260098 235220 260104 235232
rect 260156 235220 260162 235272
rect 284938 235220 284944 235272
rect 284996 235260 285002 235272
rect 301590 235260 301596 235272
rect 284996 235232 301596 235260
rect 284996 235220 285002 235232
rect 301590 235220 301596 235232
rect 301648 235220 301654 235272
rect 234062 234608 234068 234660
rect 234120 234648 234126 234660
rect 321554 234648 321560 234660
rect 234120 234620 321560 234648
rect 234120 234608 234126 234620
rect 321554 234608 321560 234620
rect 321612 234608 321618 234660
rect 153010 234540 153016 234592
rect 153068 234580 153074 234592
rect 159358 234580 159364 234592
rect 153068 234552 159364 234580
rect 153068 234540 153074 234552
rect 159358 234540 159364 234552
rect 159416 234540 159422 234592
rect 198734 234540 198740 234592
rect 198792 234580 198798 234592
rect 247218 234580 247224 234592
rect 198792 234552 247224 234580
rect 198792 234540 198798 234552
rect 247218 234540 247224 234552
rect 247276 234540 247282 234592
rect 191190 234472 191196 234524
rect 191248 234512 191254 234524
rect 204162 234512 204168 234524
rect 191248 234484 204168 234512
rect 191248 234472 191254 234484
rect 204162 234472 204168 234484
rect 204220 234472 204226 234524
rect 114646 233928 114652 233980
rect 114704 233968 114710 233980
rect 139210 233968 139216 233980
rect 114704 233940 139216 233968
rect 114704 233928 114710 233940
rect 139210 233928 139216 233940
rect 139268 233928 139274 233980
rect 139394 233928 139400 233980
rect 139452 233968 139458 233980
rect 147674 233968 147680 233980
rect 139452 233940 147680 233968
rect 139452 233928 139458 233940
rect 147674 233928 147680 233940
rect 147732 233928 147738 233980
rect 63126 233860 63132 233912
rect 63184 233900 63190 233912
rect 104158 233900 104164 233912
rect 63184 233872 104164 233900
rect 63184 233860 63190 233872
rect 104158 233860 104164 233872
rect 104216 233860 104222 233912
rect 107746 233860 107752 233912
rect 107804 233900 107810 233912
rect 146938 233900 146944 233912
rect 107804 233872 146944 233900
rect 107804 233860 107810 233872
rect 146938 233860 146944 233872
rect 146996 233860 147002 233912
rect 147766 233860 147772 233912
rect 147824 233900 147830 233912
rect 177942 233900 177948 233912
rect 147824 233872 177948 233900
rect 147824 233860 147830 233872
rect 177942 233860 177948 233872
rect 178000 233900 178006 233912
rect 178770 233900 178776 233912
rect 178000 233872 178776 233900
rect 178000 233860 178006 233872
rect 178770 233860 178776 233872
rect 178828 233860 178834 233912
rect 204162 233860 204168 233912
rect 204220 233900 204226 233912
rect 214650 233900 214656 233912
rect 204220 233872 214656 233900
rect 204220 233860 204226 233872
rect 214650 233860 214656 233872
rect 214708 233860 214714 233912
rect 215938 233792 215944 233844
rect 215996 233832 216002 233844
rect 220998 233832 221004 233844
rect 215996 233804 221004 233832
rect 215996 233792 216002 233804
rect 220998 233792 221004 233804
rect 221056 233832 221062 233844
rect 222102 233832 222108 233844
rect 221056 233804 222108 233832
rect 221056 233792 221062 233804
rect 222102 233792 222108 233804
rect 222160 233792 222166 233844
rect 159450 233248 159456 233300
rect 159508 233288 159514 233300
rect 185670 233288 185676 233300
rect 159508 233260 185676 233288
rect 159508 233248 159514 233260
rect 185670 233248 185676 233260
rect 185728 233248 185734 233300
rect 240778 233248 240784 233300
rect 240836 233288 240842 233300
rect 331398 233288 331404 233300
rect 240836 233260 331404 233288
rect 240836 233248 240842 233260
rect 331398 233248 331404 233260
rect 331456 233248 331462 233300
rect 98546 233180 98552 233232
rect 98604 233220 98610 233232
rect 155586 233220 155592 233232
rect 98604 233192 155592 233220
rect 98604 233180 98610 233192
rect 155586 233180 155592 233192
rect 155644 233180 155650 233232
rect 187050 233180 187056 233232
rect 187108 233220 187114 233232
rect 220446 233220 220452 233232
rect 187108 233192 220452 233220
rect 187108 233180 187114 233192
rect 220446 233180 220452 233192
rect 220504 233220 220510 233232
rect 220722 233220 220728 233232
rect 220504 233192 220728 233220
rect 220504 233180 220510 233192
rect 220722 233180 220728 233192
rect 220780 233180 220786 233232
rect 124582 233112 124588 233164
rect 124640 233152 124646 233164
rect 139394 233152 139400 233164
rect 124640 233124 139400 233152
rect 124640 233112 124646 233124
rect 139394 233112 139400 233124
rect 139452 233112 139458 233164
rect 146938 233112 146944 233164
rect 146996 233152 147002 233164
rect 159542 233152 159548 233164
rect 146996 233124 159548 233152
rect 146996 233112 147002 233124
rect 159542 233112 159548 233124
rect 159600 233112 159606 233164
rect 199378 233112 199384 233164
rect 199436 233152 199442 233164
rect 214558 233152 214564 233164
rect 199436 233124 214564 233152
rect 199436 233112 199442 233124
rect 214558 233112 214564 233124
rect 214616 233152 214622 233164
rect 215110 233152 215116 233164
rect 214616 233124 215116 233152
rect 214616 233112 214622 233124
rect 215110 233112 215116 233124
rect 215168 233112 215174 233164
rect 58986 232500 58992 232552
rect 59044 232540 59050 232552
rect 123478 232540 123484 232552
rect 59044 232512 123484 232540
rect 59044 232500 59050 232512
rect 123478 232500 123484 232512
rect 123536 232500 123542 232552
rect 214190 232500 214196 232552
rect 214248 232540 214254 232552
rect 258810 232540 258816 232552
rect 214248 232512 258816 232540
rect 214248 232500 214254 232512
rect 258810 232500 258816 232512
rect 258868 232500 258874 232552
rect 232038 231888 232044 231940
rect 232096 231928 232102 231940
rect 233142 231928 233148 231940
rect 232096 231900 233148 231928
rect 232096 231888 232102 231900
rect 233142 231888 233148 231900
rect 233200 231928 233206 231940
rect 233200 231900 238754 231928
rect 233200 231888 233206 231900
rect 238726 231860 238754 231900
rect 314654 231860 314660 231872
rect 238726 231832 314660 231860
rect 314654 231820 314660 231832
rect 314712 231820 314718 231872
rect 15838 231752 15844 231804
rect 15896 231792 15902 231804
rect 92474 231792 92480 231804
rect 15896 231764 92480 231792
rect 15896 231752 15902 231764
rect 92474 231752 92480 231764
rect 92532 231752 92538 231804
rect 93854 231752 93860 231804
rect 93912 231792 93918 231804
rect 94498 231792 94504 231804
rect 93912 231764 94504 231792
rect 93912 231752 93918 231764
rect 94498 231752 94504 231764
rect 94556 231792 94562 231804
rect 135990 231792 135996 231804
rect 94556 231764 135996 231792
rect 94556 231752 94562 231764
rect 135990 231752 135996 231764
rect 136048 231752 136054 231804
rect 147582 231752 147588 231804
rect 147640 231792 147646 231804
rect 155310 231792 155316 231804
rect 147640 231764 155316 231792
rect 147640 231752 147646 231764
rect 155310 231752 155316 231764
rect 155368 231752 155374 231804
rect 155862 231752 155868 231804
rect 155920 231792 155926 231804
rect 216674 231792 216680 231804
rect 155920 231764 216680 231792
rect 155920 231752 155926 231764
rect 216674 231752 216680 231764
rect 216732 231752 216738 231804
rect 136542 231684 136548 231736
rect 136600 231724 136606 231736
rect 176654 231724 176660 231736
rect 136600 231696 176660 231724
rect 136600 231684 136606 231696
rect 176654 231684 176660 231696
rect 176712 231684 176718 231736
rect 189902 231684 189908 231736
rect 189960 231724 189966 231736
rect 241238 231724 241244 231736
rect 189960 231696 241244 231724
rect 189960 231684 189966 231696
rect 241238 231684 241244 231696
rect 241296 231724 241302 231736
rect 241422 231724 241428 231736
rect 241296 231696 241428 231724
rect 241296 231684 241302 231696
rect 241422 231684 241428 231696
rect 241480 231684 241486 231736
rect 128354 231616 128360 231668
rect 128412 231656 128418 231668
rect 146018 231656 146024 231668
rect 128412 231628 146024 231656
rect 128412 231616 128418 231628
rect 146018 231616 146024 231628
rect 146076 231616 146082 231668
rect 220722 231140 220728 231192
rect 220780 231180 220786 231192
rect 253290 231180 253296 231192
rect 220780 231152 253296 231180
rect 220780 231140 220786 231152
rect 253290 231140 253296 231152
rect 253348 231140 253354 231192
rect 92474 231072 92480 231124
rect 92532 231112 92538 231124
rect 93118 231112 93124 231124
rect 92532 231084 93124 231112
rect 92532 231072 92538 231084
rect 93118 231072 93124 231084
rect 93176 231072 93182 231124
rect 176654 231072 176660 231124
rect 176712 231112 176718 231124
rect 177850 231112 177856 231124
rect 176712 231084 177856 231112
rect 176712 231072 176718 231084
rect 177850 231072 177856 231084
rect 177908 231112 177914 231124
rect 188430 231112 188436 231124
rect 177908 231084 188436 231112
rect 177908 231072 177914 231084
rect 188430 231072 188436 231084
rect 188488 231072 188494 231124
rect 241422 231072 241428 231124
rect 241480 231112 241486 231124
rect 318886 231112 318892 231124
rect 241480 231084 318892 231112
rect 241480 231072 241486 231084
rect 318886 231072 318892 231084
rect 318944 231072 318950 231124
rect 71038 230392 71044 230444
rect 71096 230432 71102 230444
rect 176010 230432 176016 230444
rect 71096 230404 176016 230432
rect 71096 230392 71102 230404
rect 176010 230392 176016 230404
rect 176068 230392 176074 230444
rect 200298 230392 200304 230444
rect 200356 230432 200362 230444
rect 202138 230432 202144 230444
rect 200356 230404 202144 230432
rect 200356 230392 200362 230404
rect 202138 230392 202144 230404
rect 202196 230392 202202 230444
rect 137922 230324 137928 230376
rect 137980 230364 137986 230376
rect 233142 230364 233148 230376
rect 137980 230336 233148 230364
rect 137980 230324 137986 230336
rect 233142 230324 233148 230336
rect 233200 230324 233206 230376
rect 66070 229712 66076 229764
rect 66128 229752 66134 229764
rect 97258 229752 97264 229764
rect 66128 229724 97264 229752
rect 66128 229712 66134 229724
rect 97258 229712 97264 229724
rect 97316 229712 97322 229764
rect 184382 229712 184388 229764
rect 184440 229752 184446 229764
rect 200114 229752 200120 229764
rect 184440 229724 200120 229752
rect 184440 229712 184446 229724
rect 200114 229712 200120 229724
rect 200172 229712 200178 229764
rect 221458 229712 221464 229764
rect 221516 229752 221522 229764
rect 229646 229752 229652 229764
rect 221516 229724 229652 229752
rect 221516 229712 221522 229724
rect 229646 229712 229652 229724
rect 229704 229712 229710 229764
rect 249058 229712 249064 229764
rect 249116 229752 249122 229764
rect 328546 229752 328552 229764
rect 249116 229724 328552 229752
rect 249116 229712 249122 229724
rect 328546 229712 328552 229724
rect 328604 229712 328610 229764
rect 57606 229032 57612 229084
rect 57664 229072 57670 229084
rect 178678 229072 178684 229084
rect 57664 229044 178684 229072
rect 57664 229032 57670 229044
rect 178678 229032 178684 229044
rect 178736 229032 178742 229084
rect 180150 229032 180156 229084
rect 180208 229072 180214 229084
rect 206830 229072 206836 229084
rect 180208 229044 206836 229072
rect 180208 229032 180214 229044
rect 206830 229032 206836 229044
rect 206888 229032 206894 229084
rect 79870 228964 79876 229016
rect 79928 229004 79934 229016
rect 173342 229004 173348 229016
rect 79928 228976 173348 229004
rect 79928 228964 79934 228976
rect 173342 228964 173348 228976
rect 173400 228964 173406 229016
rect 211062 228420 211068 228472
rect 211120 228460 211126 228472
rect 247126 228460 247132 228472
rect 211120 228432 247132 228460
rect 211120 228420 211126 228432
rect 247126 228420 247132 228432
rect 247184 228420 247190 228472
rect 220170 228352 220176 228404
rect 220228 228392 220234 228404
rect 316218 228392 316224 228404
rect 220228 228364 316224 228392
rect 220228 228352 220234 228364
rect 316218 228352 316224 228364
rect 316276 228352 316282 228404
rect 206922 227916 206928 227928
rect 200086 227888 206928 227916
rect 200086 227780 200114 227888
rect 206922 227876 206928 227888
rect 206980 227916 206986 227928
rect 208302 227916 208308 227928
rect 206980 227888 208308 227916
rect 206980 227876 206986 227888
rect 208302 227876 208308 227888
rect 208360 227876 208366 227928
rect 195256 227752 200114 227780
rect 106918 227672 106924 227724
rect 106976 227712 106982 227724
rect 195256 227712 195284 227752
rect 206278 227740 206284 227792
rect 206336 227780 206342 227792
rect 206830 227780 206836 227792
rect 206336 227752 206836 227780
rect 206336 227740 206342 227752
rect 206830 227740 206836 227752
rect 206888 227740 206894 227792
rect 106976 227684 195284 227712
rect 106976 227672 106982 227684
rect 48130 227604 48136 227656
rect 48188 227644 48194 227656
rect 118878 227644 118884 227656
rect 48188 227616 118884 227644
rect 48188 227604 48194 227616
rect 118878 227604 118884 227616
rect 118936 227604 118942 227656
rect 142062 227604 142068 227656
rect 142120 227644 142126 227656
rect 155494 227644 155500 227656
rect 142120 227616 155500 227644
rect 142120 227604 142126 227616
rect 155494 227604 155500 227616
rect 155552 227604 155558 227656
rect 192570 227604 192576 227656
rect 192628 227644 192634 227656
rect 222930 227644 222936 227656
rect 192628 227616 222936 227644
rect 192628 227604 192634 227616
rect 222930 227604 222936 227616
rect 222988 227604 222994 227656
rect 211798 226312 211804 226364
rect 211856 226352 211862 226364
rect 582650 226352 582656 226364
rect 211856 226324 582656 226352
rect 211856 226312 211862 226324
rect 582650 226312 582656 226324
rect 582708 226312 582714 226364
rect 123018 226244 123024 226296
rect 123076 226284 123082 226296
rect 173158 226284 173164 226296
rect 123076 226256 173164 226284
rect 123076 226244 123082 226256
rect 173158 226244 173164 226256
rect 173216 226284 173222 226296
rect 173342 226284 173348 226296
rect 173216 226256 173348 226284
rect 173216 226244 173222 226256
rect 173342 226244 173348 226256
rect 173400 226244 173406 226296
rect 184290 226244 184296 226296
rect 184348 226284 184354 226296
rect 222378 226284 222384 226296
rect 184348 226256 222384 226284
rect 184348 226244 184354 226256
rect 222378 226244 222384 226256
rect 222436 226244 222442 226296
rect 174722 226176 174728 226228
rect 174780 226216 174786 226228
rect 211062 226216 211068 226228
rect 174780 226188 211068 226216
rect 174780 226176 174786 226188
rect 211062 226176 211068 226188
rect 211120 226176 211126 226228
rect 146110 225564 146116 225616
rect 146168 225604 146174 225616
rect 178678 225604 178684 225616
rect 146168 225576 178684 225604
rect 146168 225564 146174 225576
rect 178678 225564 178684 225576
rect 178736 225564 178742 225616
rect 222378 225020 222384 225072
rect 222436 225060 222442 225072
rect 223022 225060 223028 225072
rect 222436 225032 223028 225060
rect 222436 225020 222442 225032
rect 223022 225020 223028 225032
rect 223080 225020 223086 225072
rect 229094 225020 229100 225072
rect 229152 225060 229158 225072
rect 229738 225060 229744 225072
rect 229152 225032 229744 225060
rect 229152 225020 229158 225032
rect 229738 225020 229744 225032
rect 229796 225060 229802 225072
rect 313366 225060 313372 225072
rect 229796 225032 313372 225060
rect 229796 225020 229802 225032
rect 313366 225020 313372 225032
rect 313424 225020 313430 225072
rect 580902 225020 580908 225072
rect 580960 225060 580966 225072
rect 583570 225060 583576 225072
rect 580960 225032 583576 225060
rect 580960 225020 580966 225032
rect 583570 225020 583576 225032
rect 583628 225020 583634 225072
rect 209866 224952 209872 225004
rect 209924 224992 209930 225004
rect 583018 224992 583024 225004
rect 209924 224964 583024 224992
rect 209924 224952 209930 224964
rect 583018 224952 583024 224964
rect 583076 224952 583082 225004
rect 130930 224884 130936 224936
rect 130988 224924 130994 224936
rect 185578 224924 185584 224936
rect 130988 224896 185584 224924
rect 130988 224884 130994 224896
rect 185578 224884 185584 224896
rect 185636 224884 185642 224936
rect 194502 224272 194508 224324
rect 194560 224312 194566 224324
rect 307754 224312 307760 224324
rect 194560 224284 307760 224312
rect 194560 224272 194566 224284
rect 307754 224272 307760 224284
rect 307812 224272 307818 224324
rect 82722 224204 82728 224256
rect 82780 224244 82786 224256
rect 195146 224244 195152 224256
rect 82780 224216 195152 224244
rect 82780 224204 82786 224216
rect 195146 224204 195152 224216
rect 195204 224204 195210 224256
rect 204990 224204 204996 224256
rect 205048 224244 205054 224256
rect 582742 224244 582748 224256
rect 205048 224216 582748 224244
rect 205048 224204 205054 224216
rect 582742 224204 582748 224216
rect 582800 224204 582806 224256
rect 86954 223524 86960 223576
rect 87012 223564 87018 223576
rect 164878 223564 164884 223576
rect 87012 223536 164884 223564
rect 87012 223524 87018 223536
rect 164878 223524 164884 223536
rect 164936 223524 164942 223576
rect 195146 223524 195152 223576
rect 195204 223564 195210 223576
rect 276014 223564 276020 223576
rect 195204 223536 276020 223564
rect 195204 223524 195210 223536
rect 276014 223524 276020 223536
rect 276072 223524 276078 223576
rect 119982 223456 119988 223508
rect 120040 223496 120046 223508
rect 187234 223496 187240 223508
rect 120040 223468 187240 223496
rect 120040 223456 120046 223468
rect 187234 223456 187240 223468
rect 187292 223456 187298 223508
rect 193030 222912 193036 222964
rect 193088 222952 193094 222964
rect 218698 222952 218704 222964
rect 193088 222924 218704 222952
rect 193088 222912 193094 222924
rect 218698 222912 218704 222924
rect 218756 222912 218762 222964
rect 169018 222844 169024 222896
rect 169076 222884 169082 222896
rect 195146 222884 195152 222896
rect 169076 222856 195152 222884
rect 169076 222844 169082 222856
rect 195146 222844 195152 222856
rect 195204 222844 195210 222896
rect 97258 222096 97264 222148
rect 97316 222136 97322 222148
rect 195054 222136 195060 222148
rect 97316 222108 195060 222136
rect 97316 222096 97322 222108
rect 195054 222096 195060 222108
rect 195112 222096 195118 222148
rect 195146 222096 195152 222148
rect 195204 222136 195210 222148
rect 219618 222136 219624 222148
rect 195204 222108 219624 222136
rect 195204 222096 195210 222108
rect 219618 222096 219624 222108
rect 219676 222096 219682 222148
rect 214650 221484 214656 221536
rect 214708 221524 214714 221536
rect 233970 221524 233976 221536
rect 214708 221496 233976 221524
rect 214708 221484 214714 221496
rect 233970 221484 233976 221496
rect 234028 221484 234034 221536
rect 238662 221484 238668 221536
rect 238720 221524 238726 221536
rect 267826 221524 267832 221536
rect 238720 221496 267832 221524
rect 238720 221484 238726 221496
rect 267826 221484 267832 221496
rect 267884 221484 267890 221536
rect 133874 221416 133880 221468
rect 133932 221456 133938 221468
rect 215202 221456 215208 221468
rect 133932 221428 215208 221456
rect 133932 221416 133938 221428
rect 215202 221416 215208 221428
rect 215260 221416 215266 221468
rect 232682 221416 232688 221468
rect 232740 221456 232746 221468
rect 282086 221456 282092 221468
rect 232740 221428 282092 221456
rect 232740 221416 232746 221428
rect 282086 221416 282092 221428
rect 282144 221416 282150 221468
rect 75822 220736 75828 220788
rect 75880 220776 75886 220788
rect 172422 220776 172428 220788
rect 75880 220748 172428 220776
rect 75880 220736 75886 220748
rect 172422 220736 172428 220748
rect 172480 220736 172486 220788
rect 191282 220736 191288 220788
rect 191340 220776 191346 220788
rect 249978 220776 249984 220788
rect 191340 220748 249984 220776
rect 191340 220736 191346 220748
rect 249978 220736 249984 220748
rect 250036 220776 250042 220788
rect 251082 220776 251088 220788
rect 250036 220748 251088 220776
rect 250036 220736 250042 220748
rect 251082 220736 251088 220748
rect 251140 220736 251146 220788
rect 49602 220668 49608 220720
rect 49660 220708 49666 220720
rect 94498 220708 94504 220720
rect 49660 220680 94504 220708
rect 49660 220668 49666 220680
rect 94498 220668 94504 220680
rect 94556 220668 94562 220720
rect 251082 220124 251088 220176
rect 251140 220164 251146 220176
rect 281534 220164 281540 220176
rect 251140 220136 281540 220164
rect 251140 220124 251146 220136
rect 281534 220124 281540 220136
rect 281592 220124 281598 220176
rect 14458 220056 14464 220108
rect 14516 220096 14522 220108
rect 49602 220096 49608 220108
rect 14516 220068 49608 220096
rect 14516 220056 14522 220068
rect 49602 220056 49608 220068
rect 49660 220056 49666 220108
rect 104158 220056 104164 220108
rect 104216 220096 104222 220108
rect 191834 220096 191840 220108
rect 104216 220068 191840 220096
rect 104216 220056 104222 220068
rect 191834 220056 191840 220068
rect 191892 220056 191898 220108
rect 200022 220056 200028 220108
rect 200080 220096 200086 220108
rect 266538 220096 266544 220108
rect 200080 220068 266544 220096
rect 200080 220056 200086 220068
rect 266538 220056 266544 220068
rect 266596 220056 266602 220108
rect 282086 220056 282092 220108
rect 282144 220096 282150 220108
rect 298830 220096 298836 220108
rect 282144 220068 298836 220096
rect 282144 220056 282150 220068
rect 298830 220056 298836 220068
rect 298888 220056 298894 220108
rect 195790 219444 195796 219496
rect 195848 219484 195854 219496
rect 198090 219484 198096 219496
rect 195848 219456 198096 219484
rect 195848 219444 195854 219456
rect 198090 219444 198096 219456
rect 198148 219444 198154 219496
rect 99466 219376 99472 219428
rect 99524 219416 99530 219428
rect 212626 219416 212632 219428
rect 99524 219388 212632 219416
rect 99524 219376 99530 219388
rect 212626 219376 212632 219388
rect 212684 219376 212690 219428
rect 215202 218832 215208 218884
rect 215260 218872 215266 218884
rect 245562 218872 245568 218884
rect 215260 218844 245568 218872
rect 215260 218832 215266 218844
rect 245562 218832 245568 218844
rect 245620 218832 245626 218884
rect 224218 218764 224224 218816
rect 224276 218804 224282 218816
rect 270770 218804 270776 218816
rect 224276 218776 270776 218804
rect 224276 218764 224282 218776
rect 270770 218764 270776 218776
rect 270828 218764 270834 218816
rect 122650 218696 122656 218748
rect 122708 218736 122714 218748
rect 224862 218736 224868 218748
rect 122708 218708 224868 218736
rect 122708 218696 122714 218708
rect 224862 218696 224868 218708
rect 224920 218696 224926 218748
rect 52178 217948 52184 218000
rect 52236 217988 52242 218000
rect 159450 217988 159456 218000
rect 52236 217960 159456 217988
rect 52236 217948 52242 217960
rect 159450 217948 159456 217960
rect 159508 217948 159514 218000
rect 122834 217880 122840 217932
rect 122892 217920 122898 217932
rect 217318 217920 217324 217932
rect 122892 217892 217324 217920
rect 122892 217880 122898 217892
rect 217318 217880 217324 217892
rect 217376 217880 217382 217932
rect 258810 217268 258816 217320
rect 258868 217308 258874 217320
rect 335538 217308 335544 217320
rect 258868 217280 335544 217308
rect 258868 217268 258874 217280
rect 335538 217268 335544 217280
rect 335596 217268 335602 217320
rect 181990 216696 181996 216708
rect 180766 216668 181996 216696
rect 81618 216588 81624 216640
rect 81676 216628 81682 216640
rect 180766 216628 180794 216668
rect 181990 216656 181996 216668
rect 182048 216696 182054 216708
rect 191190 216696 191196 216708
rect 182048 216668 191196 216696
rect 182048 216656 182054 216668
rect 191190 216656 191196 216668
rect 191248 216656 191254 216708
rect 192570 216656 192576 216708
rect 192628 216696 192634 216708
rect 249886 216696 249892 216708
rect 192628 216668 249892 216696
rect 192628 216656 192634 216668
rect 249886 216656 249892 216668
rect 249944 216696 249950 216708
rect 250622 216696 250628 216708
rect 249944 216668 250628 216696
rect 249944 216656 249950 216668
rect 250622 216656 250628 216668
rect 250680 216656 250686 216708
rect 81676 216600 180794 216628
rect 81676 216588 81682 216600
rect 178678 216520 178684 216572
rect 178736 216560 178742 216572
rect 262214 216560 262220 216572
rect 178736 216532 262220 216560
rect 178736 216520 178742 216532
rect 262214 216520 262220 216532
rect 262272 216520 262278 216572
rect 103422 216452 103428 216504
rect 103480 216492 103486 216504
rect 178034 216492 178040 216504
rect 103480 216464 178040 216492
rect 103480 216452 103486 216464
rect 178034 216452 178040 216464
rect 178092 216452 178098 216504
rect 204990 215908 204996 215960
rect 205048 215948 205054 215960
rect 240778 215948 240784 215960
rect 205048 215920 240784 215948
rect 205048 215908 205054 215920
rect 240778 215908 240784 215920
rect 240836 215908 240842 215960
rect 286318 215908 286324 215960
rect 286376 215948 286382 215960
rect 316126 215948 316132 215960
rect 286376 215920 316132 215948
rect 286376 215908 286382 215920
rect 316126 215908 316132 215920
rect 316184 215908 316190 215960
rect 262214 215296 262220 215348
rect 262272 215336 262278 215348
rect 262950 215336 262956 215348
rect 262272 215308 262956 215336
rect 262272 215296 262278 215308
rect 262950 215296 262956 215308
rect 263008 215296 263014 215348
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 22738 215268 22744 215280
rect 3384 215240 22744 215268
rect 3384 215228 3390 215240
rect 22738 215228 22744 215240
rect 22796 215228 22802 215280
rect 132310 215228 132316 215280
rect 132368 215268 132374 215280
rect 256694 215268 256700 215280
rect 132368 215240 256700 215268
rect 132368 215228 132374 215240
rect 256694 215228 256700 215240
rect 256752 215228 256758 215280
rect 144730 215160 144736 215212
rect 144788 215200 144794 215212
rect 235994 215200 236000 215212
rect 144788 215172 236000 215200
rect 144788 215160 144794 215172
rect 235994 215160 236000 215172
rect 236052 215160 236058 215212
rect 256694 214752 256700 214804
rect 256752 214792 256758 214804
rect 257338 214792 257344 214804
rect 256752 214764 257344 214792
rect 256752 214752 256758 214764
rect 257338 214752 257344 214764
rect 257396 214752 257402 214804
rect 158070 213868 158076 213920
rect 158128 213908 158134 213920
rect 269114 213908 269120 213920
rect 158128 213880 269120 213908
rect 158128 213868 158134 213880
rect 269114 213868 269120 213880
rect 269172 213868 269178 213920
rect 171870 213800 171876 213852
rect 171928 213840 171934 213852
rect 247034 213840 247040 213852
rect 171928 213812 247040 213840
rect 171928 213800 171934 213812
rect 247034 213800 247040 213812
rect 247092 213800 247098 213852
rect 46842 213188 46848 213240
rect 46900 213228 46906 213240
rect 171962 213228 171968 213240
rect 46900 213200 171968 213228
rect 46900 213188 46906 213200
rect 171962 213188 171968 213200
rect 172020 213188 172026 213240
rect 113082 211828 113088 211880
rect 113140 211868 113146 211880
rect 194778 211868 194784 211880
rect 113140 211840 194784 211868
rect 113140 211828 113146 211840
rect 194778 211828 194784 211840
rect 194836 211828 194842 211880
rect 39298 211760 39304 211812
rect 39356 211800 39362 211812
rect 164234 211800 164240 211812
rect 39356 211772 164240 211800
rect 39356 211760 39362 211772
rect 164234 211760 164240 211772
rect 164292 211760 164298 211812
rect 193122 211760 193128 211812
rect 193180 211800 193186 211812
rect 242158 211800 242164 211812
rect 193180 211772 242164 211800
rect 193180 211760 193186 211772
rect 242158 211760 242164 211772
rect 242216 211760 242222 211812
rect 288618 211188 288624 211200
rect 213840 211160 288624 211188
rect 191650 211080 191656 211132
rect 191708 211120 191714 211132
rect 213840 211120 213868 211160
rect 288618 211148 288624 211160
rect 288676 211148 288682 211200
rect 191708 211092 213868 211120
rect 191708 211080 191714 211092
rect 193122 211012 193128 211064
rect 193180 211052 193186 211064
rect 194134 211052 194140 211064
rect 193180 211024 194140 211052
rect 193180 211012 193186 211024
rect 194134 211012 194140 211024
rect 194192 211012 194198 211064
rect 151078 210536 151084 210588
rect 151136 210576 151142 210588
rect 191098 210576 191104 210588
rect 151136 210548 191104 210576
rect 151136 210536 151142 210548
rect 191098 210536 191104 210548
rect 191156 210536 191162 210588
rect 131022 210468 131028 210520
rect 131080 210508 131086 210520
rect 193122 210508 193128 210520
rect 131080 210480 193128 210508
rect 131080 210468 131086 210480
rect 193122 210468 193128 210480
rect 193180 210468 193186 210520
rect 70394 210400 70400 210452
rect 70452 210440 70458 210452
rect 150434 210440 150440 210452
rect 70452 210412 150440 210440
rect 70452 210400 70458 210412
rect 150434 210400 150440 210412
rect 150492 210400 150498 210452
rect 212626 210400 212632 210452
rect 212684 210440 212690 210452
rect 258810 210440 258816 210452
rect 212684 210412 258816 210440
rect 212684 210400 212690 210412
rect 258810 210400 258816 210412
rect 258868 210400 258874 210452
rect 278038 210400 278044 210452
rect 278096 210440 278102 210452
rect 294690 210440 294696 210452
rect 278096 210412 294696 210440
rect 278096 210400 278102 210412
rect 294690 210400 294696 210412
rect 294748 210400 294754 210452
rect 69014 209720 69020 209772
rect 69072 209760 69078 209772
rect 231118 209760 231124 209772
rect 69072 209732 231124 209760
rect 69072 209720 69078 209732
rect 231118 209720 231124 209732
rect 231176 209720 231182 209772
rect 92382 209652 92388 209704
rect 92440 209692 92446 209704
rect 209038 209692 209044 209704
rect 92440 209664 209044 209692
rect 92440 209652 92446 209664
rect 209038 209652 209044 209664
rect 209096 209652 209102 209704
rect 231118 209040 231124 209092
rect 231176 209080 231182 209092
rect 277486 209080 277492 209092
rect 231176 209052 277492 209080
rect 231176 209040 231182 209052
rect 277486 209040 277492 209052
rect 277544 209040 277550 209092
rect 208394 208360 208400 208412
rect 208452 208400 208458 208412
rect 209682 208400 209688 208412
rect 208452 208372 209688 208400
rect 208452 208360 208458 208372
rect 209682 208360 209688 208372
rect 209740 208400 209746 208412
rect 281626 208400 281632 208412
rect 209740 208372 281632 208400
rect 209740 208360 209746 208372
rect 281626 208360 281632 208372
rect 281684 208360 281690 208412
rect 53650 208292 53656 208344
rect 53708 208332 53714 208344
rect 244274 208332 244280 208344
rect 53708 208304 244280 208332
rect 53708 208292 53714 208304
rect 244274 208292 244280 208304
rect 244332 208292 244338 208344
rect 85574 207612 85580 207664
rect 85632 207652 85638 207664
rect 214650 207652 214656 207664
rect 85632 207624 214656 207652
rect 85632 207612 85638 207624
rect 214650 207612 214656 207624
rect 214708 207612 214714 207664
rect 218974 207612 218980 207664
rect 219032 207652 219038 207664
rect 311986 207652 311992 207664
rect 219032 207624 311992 207652
rect 219032 207612 219038 207624
rect 311986 207612 311992 207624
rect 312044 207612 312050 207664
rect 244274 207000 244280 207052
rect 244332 207040 244338 207052
rect 244918 207040 244924 207052
rect 244332 207012 244924 207040
rect 244332 207000 244338 207012
rect 244918 207000 244924 207012
rect 244976 207000 244982 207052
rect 89530 206932 89536 206984
rect 89588 206972 89594 206984
rect 192570 206972 192576 206984
rect 89588 206944 192576 206972
rect 89588 206932 89594 206944
rect 192570 206932 192576 206944
rect 192628 206932 192634 206984
rect 194778 206932 194784 206984
rect 194836 206972 194842 206984
rect 258074 206972 258080 206984
rect 194836 206944 258080 206972
rect 194836 206932 194842 206944
rect 258074 206932 258080 206944
rect 258132 206972 258138 206984
rect 259362 206972 259368 206984
rect 258132 206944 259368 206972
rect 258132 206932 258138 206944
rect 259362 206932 259368 206944
rect 259420 206932 259426 206984
rect 110322 206864 110328 206916
rect 110380 206904 110386 206916
rect 184290 206904 184296 206916
rect 110380 206876 184296 206904
rect 110380 206864 110386 206876
rect 184290 206864 184296 206876
rect 184348 206864 184354 206916
rect 259362 206320 259368 206372
rect 259420 206360 259426 206372
rect 278774 206360 278780 206372
rect 259420 206332 278780 206360
rect 259420 206320 259426 206332
rect 278774 206320 278780 206332
rect 278832 206320 278838 206372
rect 222838 206252 222844 206304
rect 222896 206292 222902 206304
rect 308398 206292 308404 206304
rect 222896 206264 308404 206292
rect 222896 206252 222902 206264
rect 308398 206252 308404 206264
rect 308456 206252 308462 206304
rect 125410 205572 125416 205624
rect 125468 205612 125474 205624
rect 251174 205612 251180 205624
rect 125468 205584 251180 205612
rect 125468 205572 125474 205584
rect 251174 205572 251180 205584
rect 251232 205612 251238 205624
rect 252462 205612 252468 205624
rect 251232 205584 252468 205612
rect 251232 205572 251238 205584
rect 252462 205572 252468 205584
rect 252520 205572 252526 205624
rect 72418 204892 72424 204944
rect 72476 204932 72482 204944
rect 233142 204932 233148 204944
rect 72476 204904 233148 204932
rect 72476 204892 72482 204904
rect 233142 204892 233148 204904
rect 233200 204932 233206 204944
rect 234430 204932 234436 204944
rect 233200 204904 234436 204932
rect 233200 204892 233206 204904
rect 234430 204892 234436 204904
rect 234488 204892 234494 204944
rect 252462 204892 252468 204944
rect 252520 204932 252526 204944
rect 273346 204932 273352 204944
rect 252520 204904 273352 204932
rect 252520 204892 252526 204904
rect 273346 204892 273352 204904
rect 273404 204892 273410 204944
rect 67174 204212 67180 204264
rect 67232 204252 67238 204264
rect 213730 204252 213736 204264
rect 67232 204224 213736 204252
rect 67232 204212 67238 204224
rect 213730 204212 213736 204224
rect 213788 204212 213794 204264
rect 150434 204144 150440 204196
rect 150492 204184 150498 204196
rect 215662 204184 215668 204196
rect 150492 204156 215668 204184
rect 150492 204144 150498 204156
rect 215662 204144 215668 204156
rect 215720 204144 215726 204196
rect 214558 203532 214564 203584
rect 214616 203572 214622 203584
rect 264054 203572 264060 203584
rect 214616 203544 264060 203572
rect 214616 203532 214622 203544
rect 264054 203532 264060 203544
rect 264112 203532 264118 203584
rect 3418 202784 3424 202836
rect 3476 202824 3482 202836
rect 126790 202824 126796 202836
rect 3476 202796 126796 202824
rect 3476 202784 3482 202796
rect 126790 202784 126796 202796
rect 126848 202784 126854 202836
rect 97810 202716 97816 202768
rect 97868 202756 97874 202768
rect 157978 202756 157984 202768
rect 97868 202728 157984 202756
rect 97868 202716 97874 202728
rect 157978 202716 157984 202728
rect 158036 202716 158042 202768
rect 154482 202172 154488 202224
rect 154540 202212 154546 202224
rect 173250 202212 173256 202224
rect 154540 202184 173256 202212
rect 154540 202172 154546 202184
rect 173250 202172 173256 202184
rect 173308 202172 173314 202224
rect 201310 202172 201316 202224
rect 201368 202212 201374 202224
rect 276014 202212 276020 202224
rect 201368 202184 276020 202212
rect 201368 202172 201374 202184
rect 276014 202172 276020 202184
rect 276072 202172 276078 202224
rect 171042 202104 171048 202156
rect 171100 202144 171106 202156
rect 292022 202144 292028 202156
rect 171100 202116 292028 202144
rect 171100 202104 171106 202116
rect 292022 202104 292028 202116
rect 292080 202104 292086 202156
rect 77202 201424 77208 201476
rect 77260 201464 77266 201476
rect 221366 201464 221372 201476
rect 77260 201436 221372 201464
rect 77260 201424 77266 201436
rect 221366 201424 221372 201436
rect 221424 201424 221430 201476
rect 144822 201356 144828 201408
rect 144880 201396 144886 201408
rect 204990 201396 204996 201408
rect 144880 201368 204996 201396
rect 144880 201356 144886 201368
rect 204990 201356 204996 201368
rect 205048 201356 205054 201408
rect 226150 200812 226156 200864
rect 226208 200852 226214 200864
rect 314746 200852 314752 200864
rect 226208 200824 314752 200852
rect 226208 200812 226214 200824
rect 314746 200812 314752 200824
rect 314804 200812 314810 200864
rect 206370 200744 206376 200796
rect 206428 200784 206434 200796
rect 304258 200784 304264 200796
rect 206428 200756 304264 200784
rect 206428 200744 206434 200756
rect 304258 200744 304264 200756
rect 304316 200744 304322 200796
rect 139302 200064 139308 200116
rect 139360 200104 139366 200116
rect 166258 200104 166264 200116
rect 139360 200076 166264 200104
rect 139360 200064 139366 200076
rect 166258 200064 166264 200076
rect 166316 200064 166322 200116
rect 203518 199452 203524 199504
rect 203576 199492 203582 199504
rect 320358 199492 320364 199504
rect 203576 199464 320364 199492
rect 203576 199452 203582 199464
rect 320358 199452 320364 199464
rect 320416 199452 320422 199504
rect 111610 199384 111616 199436
rect 111668 199424 111674 199436
rect 233878 199424 233884 199436
rect 111668 199396 233884 199424
rect 111668 199384 111674 199396
rect 233878 199384 233884 199396
rect 233936 199384 233942 199436
rect 115198 198636 115204 198688
rect 115256 198676 115262 198688
rect 186958 198676 186964 198688
rect 115256 198648 186964 198676
rect 115256 198636 115262 198648
rect 186958 198636 186964 198648
rect 187016 198636 187022 198688
rect 207658 198024 207664 198076
rect 207716 198064 207722 198076
rect 297450 198064 297456 198076
rect 207716 198036 297456 198064
rect 207716 198024 207722 198036
rect 297450 198024 297456 198036
rect 297508 198024 297514 198076
rect 183462 197956 183468 198008
rect 183520 197996 183526 198008
rect 306466 197996 306472 198008
rect 183520 197968 306472 197996
rect 183520 197956 183526 197968
rect 306466 197956 306472 197968
rect 306524 197956 306530 198008
rect 74442 197276 74448 197328
rect 74500 197316 74506 197328
rect 200758 197316 200764 197328
rect 74500 197288 200764 197316
rect 74500 197276 74506 197288
rect 200758 197276 200764 197288
rect 200816 197276 200822 197328
rect 201402 196664 201408 196716
rect 201460 196704 201466 196716
rect 300210 196704 300216 196716
rect 201460 196676 300216 196704
rect 201460 196664 201466 196676
rect 300210 196664 300216 196676
rect 300268 196664 300274 196716
rect 148962 196596 148968 196648
rect 149020 196636 149026 196648
rect 182818 196636 182824 196648
rect 149020 196608 182824 196636
rect 149020 196596 149026 196608
rect 182818 196596 182824 196608
rect 182876 196596 182882 196648
rect 186958 196596 186964 196648
rect 187016 196636 187022 196648
rect 314838 196636 314844 196648
rect 187016 196608 314844 196636
rect 187016 196596 187022 196608
rect 314838 196596 314844 196608
rect 314896 196596 314902 196648
rect 52270 195916 52276 195968
rect 52328 195956 52334 195968
rect 207750 195956 207756 195968
rect 52328 195928 207756 195956
rect 52328 195916 52334 195928
rect 207750 195916 207756 195928
rect 207808 195916 207814 195968
rect 122742 195236 122748 195288
rect 122800 195276 122806 195288
rect 185578 195276 185584 195288
rect 122800 195248 185584 195276
rect 122800 195236 122806 195248
rect 185578 195236 185584 195248
rect 185636 195236 185642 195288
rect 186222 195236 186228 195288
rect 186280 195276 186286 195288
rect 264330 195276 264336 195288
rect 186280 195248 264336 195276
rect 186280 195236 186286 195248
rect 264330 195236 264336 195248
rect 264388 195236 264394 195288
rect 247770 194556 247776 194608
rect 247828 194596 247834 194608
rect 284294 194596 284300 194608
rect 247828 194568 284300 194596
rect 247828 194556 247834 194568
rect 284294 194556 284300 194568
rect 284352 194556 284358 194608
rect 93118 194488 93124 194540
rect 93176 194528 93182 194540
rect 212718 194528 212724 194540
rect 93176 194500 212724 194528
rect 93176 194488 93182 194500
rect 212718 194488 212724 194500
rect 212776 194488 212782 194540
rect 233970 193876 233976 193928
rect 234028 193916 234034 193928
rect 285674 193916 285680 193928
rect 234028 193888 285680 193916
rect 234028 193876 234034 193888
rect 285674 193876 285680 193888
rect 285732 193876 285738 193928
rect 100662 193808 100668 193860
rect 100720 193848 100726 193860
rect 236638 193848 236644 193860
rect 100720 193820 236644 193848
rect 100720 193808 100726 193820
rect 236638 193808 236644 193820
rect 236696 193808 236702 193860
rect 156598 192516 156604 192568
rect 156656 192556 156662 192568
rect 202322 192556 202328 192568
rect 156656 192528 202328 192556
rect 156656 192516 156662 192528
rect 202322 192516 202328 192528
rect 202380 192516 202386 192568
rect 242250 192516 242256 192568
rect 242308 192556 242314 192568
rect 325878 192556 325884 192568
rect 242308 192528 325884 192556
rect 242308 192516 242314 192528
rect 325878 192516 325884 192528
rect 325936 192516 325942 192568
rect 132402 192448 132408 192500
rect 132460 192488 132466 192500
rect 178770 192488 178776 192500
rect 132460 192460 178776 192488
rect 132460 192448 132466 192460
rect 178770 192448 178776 192460
rect 178828 192448 178834 192500
rect 201494 192448 201500 192500
rect 201552 192488 201558 192500
rect 310606 192488 310612 192500
rect 201552 192460 310612 192488
rect 201552 192448 201558 192460
rect 310606 192448 310612 192460
rect 310664 192448 310670 192500
rect 97902 191088 97908 191140
rect 97960 191128 97966 191140
rect 251174 191128 251180 191140
rect 97960 191100 251180 191128
rect 97960 191088 97966 191100
rect 251174 191088 251180 191100
rect 251232 191088 251238 191140
rect 106182 190476 106188 190528
rect 106240 190516 106246 190528
rect 217318 190516 217324 190528
rect 106240 190488 217324 190516
rect 106240 190476 106246 190488
rect 217318 190476 217324 190488
rect 217376 190476 217382 190528
rect 242158 189796 242164 189848
rect 242216 189836 242222 189848
rect 269390 189836 269396 189848
rect 242216 189808 269396 189836
rect 242216 189796 242222 189808
rect 269390 189796 269396 189808
rect 269448 189796 269454 189848
rect 217410 189728 217416 189780
rect 217468 189768 217474 189780
rect 305178 189768 305184 189780
rect 217468 189740 305184 189768
rect 217468 189728 217474 189740
rect 305178 189728 305184 189740
rect 305236 189728 305242 189780
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 35158 189020 35164 189032
rect 3568 188992 35164 189020
rect 3568 188980 3574 188992
rect 35158 188980 35164 188992
rect 35216 188980 35222 189032
rect 67542 188980 67548 189032
rect 67600 189020 67606 189032
rect 218422 189020 218428 189032
rect 67600 188992 218428 189020
rect 67600 188980 67606 188992
rect 218422 188980 218428 188992
rect 218480 188980 218486 189032
rect 178862 188300 178868 188352
rect 178920 188340 178926 188352
rect 232590 188340 232596 188352
rect 178920 188312 232596 188340
rect 178920 188300 178926 188312
rect 232590 188300 232596 188312
rect 232648 188300 232654 188352
rect 233142 188300 233148 188352
rect 233200 188340 233206 188352
rect 265066 188340 265072 188352
rect 233200 188312 265072 188340
rect 233200 188300 233206 188312
rect 265066 188300 265072 188312
rect 265124 188300 265130 188352
rect 294690 188300 294696 188352
rect 294748 188340 294754 188352
rect 302326 188340 302332 188352
rect 294748 188312 302332 188340
rect 294748 188300 294754 188312
rect 302326 188300 302332 188312
rect 302384 188300 302390 188352
rect 251818 187688 251824 187740
rect 251876 187728 251882 187740
rect 283098 187728 283104 187740
rect 251876 187700 283104 187728
rect 251876 187688 251882 187700
rect 283098 187688 283104 187700
rect 283156 187688 283162 187740
rect 298830 187076 298836 187128
rect 298888 187116 298894 187128
rect 302418 187116 302424 187128
rect 298888 187088 302424 187116
rect 298888 187076 298894 187088
rect 302418 187076 302424 187088
rect 302476 187076 302482 187128
rect 202138 187008 202144 187060
rect 202196 187048 202202 187060
rect 309410 187048 309416 187060
rect 202196 187020 309416 187048
rect 202196 187008 202202 187020
rect 309410 187008 309416 187020
rect 309468 187008 309474 187060
rect 115842 186940 115848 186992
rect 115900 186980 115906 186992
rect 242158 186980 242164 186992
rect 115900 186952 242164 186980
rect 115900 186940 115906 186952
rect 242158 186940 242164 186952
rect 242216 186940 242222 186992
rect 254578 186940 254584 186992
rect 254636 186980 254642 186992
rect 276106 186980 276112 186992
rect 254636 186952 276112 186980
rect 254636 186940 254642 186952
rect 276106 186940 276112 186952
rect 276164 186940 276170 186992
rect 119982 186328 119988 186380
rect 120040 186368 120046 186380
rect 164878 186368 164884 186380
rect 120040 186340 164884 186368
rect 120040 186328 120046 186340
rect 164878 186328 164884 186340
rect 164936 186328 164942 186380
rect 302326 185784 302332 185836
rect 302384 185824 302390 185836
rect 304442 185824 304448 185836
rect 302384 185796 304448 185824
rect 302384 185784 302390 185796
rect 304442 185784 304448 185796
rect 304500 185784 304506 185836
rect 190362 185648 190368 185700
rect 190420 185688 190426 185700
rect 310790 185688 310796 185700
rect 190420 185660 310796 185688
rect 190420 185648 190426 185660
rect 310790 185648 310796 185660
rect 310848 185648 310854 185700
rect 91002 185580 91008 185632
rect 91060 185620 91066 185632
rect 231118 185620 231124 185632
rect 91060 185592 231124 185620
rect 91060 185580 91066 185592
rect 231118 185580 231124 185592
rect 231176 185580 231182 185632
rect 121362 184900 121368 184952
rect 121420 184940 121426 184952
rect 167914 184940 167920 184952
rect 121420 184912 167920 184940
rect 121420 184900 121426 184912
rect 167914 184900 167920 184912
rect 167972 184900 167978 184952
rect 245562 184220 245568 184272
rect 245620 184260 245626 184272
rect 265250 184260 265256 184272
rect 245620 184232 265256 184260
rect 245620 184220 245626 184232
rect 265250 184220 265256 184232
rect 265308 184220 265314 184272
rect 301590 184220 301596 184272
rect 301648 184260 301654 184272
rect 313458 184260 313464 184272
rect 301648 184232 313464 184260
rect 301648 184220 301654 184232
rect 313458 184220 313464 184232
rect 313516 184220 313522 184272
rect 177942 184152 177948 184204
rect 178000 184192 178006 184204
rect 277578 184192 277584 184204
rect 178000 184164 277584 184192
rect 178000 184152 178006 184164
rect 277578 184152 277584 184164
rect 277636 184152 277642 184204
rect 286502 184152 286508 184204
rect 286560 184192 286566 184204
rect 312078 184192 312084 184204
rect 286560 184164 312084 184192
rect 286560 184152 286566 184164
rect 312078 184152 312084 184164
rect 312136 184152 312142 184204
rect 148962 183608 148968 183660
rect 149020 183648 149026 183660
rect 167638 183648 167644 183660
rect 149020 183620 167644 183648
rect 149020 183608 149026 183620
rect 167638 183608 167644 183620
rect 167696 183608 167702 183660
rect 129642 183540 129648 183592
rect 129700 183580 129706 183592
rect 233970 183580 233976 183592
rect 129700 183552 233976 183580
rect 129700 183540 129706 183552
rect 233970 183540 233976 183552
rect 234028 183540 234034 183592
rect 304350 183472 304356 183524
rect 304408 183512 304414 183524
rect 305270 183512 305276 183524
rect 304408 183484 305276 183512
rect 304408 183472 304414 183484
rect 305270 183472 305276 183484
rect 305328 183472 305334 183524
rect 261570 182860 261576 182912
rect 261628 182900 261634 182912
rect 276198 182900 276204 182912
rect 261628 182872 276204 182900
rect 261628 182860 261634 182872
rect 276198 182860 276204 182872
rect 276256 182860 276262 182912
rect 276658 182860 276664 182912
rect 276716 182900 276722 182912
rect 303798 182900 303804 182912
rect 276716 182872 303804 182900
rect 276716 182860 276722 182872
rect 303798 182860 303804 182872
rect 303856 182860 303862 182912
rect 184842 182792 184848 182844
rect 184900 182832 184906 182844
rect 323118 182832 323124 182844
rect 184900 182804 323124 182832
rect 184900 182792 184906 182804
rect 323118 182792 323124 182804
rect 323176 182792 323182 182844
rect 103330 182248 103336 182300
rect 103388 182288 103394 182300
rect 170490 182288 170496 182300
rect 103388 182260 170496 182288
rect 103388 182248 103394 182260
rect 170490 182248 170496 182260
rect 170548 182248 170554 182300
rect 113726 182180 113732 182232
rect 113784 182220 113790 182232
rect 231210 182220 231216 182232
rect 113784 182192 231216 182220
rect 113784 182180 113790 182192
rect 231210 182180 231216 182192
rect 231268 182180 231274 182232
rect 302418 182112 302424 182164
rect 302476 182152 302482 182164
rect 303706 182152 303712 182164
rect 302476 182124 303712 182152
rect 302476 182112 302482 182124
rect 303706 182112 303712 182124
rect 303764 182112 303770 182164
rect 238018 181500 238024 181552
rect 238076 181540 238082 181552
rect 270586 181540 270592 181552
rect 238076 181512 270592 181540
rect 238076 181500 238082 181512
rect 270586 181500 270592 181512
rect 270644 181500 270650 181552
rect 296070 181500 296076 181552
rect 296128 181540 296134 181552
rect 308030 181540 308036 181552
rect 296128 181512 308036 181540
rect 296128 181500 296134 181512
rect 308030 181500 308036 181512
rect 308088 181500 308094 181552
rect 167822 181432 167828 181484
rect 167880 181472 167886 181484
rect 203518 181472 203524 181484
rect 167880 181444 203524 181472
rect 167880 181432 167886 181444
rect 203518 181432 203524 181444
rect 203576 181432 203582 181484
rect 203610 181432 203616 181484
rect 203668 181472 203674 181484
rect 301038 181472 301044 181484
rect 203668 181444 301044 181472
rect 203668 181432 203674 181444
rect 301038 181432 301044 181444
rect 301096 181432 301102 181484
rect 308398 181432 308404 181484
rect 308456 181472 308462 181484
rect 321738 181472 321744 181484
rect 308456 181444 321744 181472
rect 308456 181432 308462 181444
rect 321738 181432 321744 181444
rect 321796 181432 321802 181484
rect 132494 180888 132500 180940
rect 132552 180928 132558 180940
rect 169110 180928 169116 180940
rect 132552 180900 169116 180928
rect 132552 180888 132558 180900
rect 169110 180888 169116 180900
rect 169168 180888 169174 180940
rect 126054 180820 126060 180872
rect 126112 180860 126118 180872
rect 166442 180860 166448 180872
rect 126112 180832 166448 180860
rect 126112 180820 126118 180832
rect 166442 180820 166448 180832
rect 166500 180820 166506 180872
rect 262858 180140 262864 180192
rect 262916 180180 262922 180192
rect 272058 180180 272064 180192
rect 262916 180152 272064 180180
rect 262916 180140 262922 180152
rect 272058 180140 272064 180152
rect 272116 180140 272122 180192
rect 293218 180140 293224 180192
rect 293276 180180 293282 180192
rect 310698 180180 310704 180192
rect 293276 180152 310704 180180
rect 293276 180140 293282 180152
rect 310698 180140 310704 180152
rect 310756 180140 310762 180192
rect 253290 180072 253296 180124
rect 253348 180112 253354 180124
rect 269298 180112 269304 180124
rect 253348 180084 269304 180112
rect 253348 180072 253354 180084
rect 269298 180072 269304 180084
rect 269356 180072 269362 180124
rect 290458 180072 290464 180124
rect 290516 180112 290522 180124
rect 313550 180112 313556 180124
rect 290516 180084 313556 180112
rect 290516 180072 290522 180084
rect 313550 180072 313556 180084
rect 313608 180072 313614 180124
rect 313918 179868 313924 179920
rect 313976 179908 313982 179920
rect 317690 179908 317696 179920
rect 313976 179880 317696 179908
rect 313976 179868 313982 179880
rect 317690 179868 317696 179880
rect 317748 179868 317754 179920
rect 118510 179460 118516 179512
rect 118568 179500 118574 179512
rect 184382 179500 184388 179512
rect 118568 179472 184388 179500
rect 118568 179460 118574 179472
rect 184382 179460 184388 179472
rect 184440 179460 184446 179512
rect 132402 179392 132408 179444
rect 132460 179432 132466 179444
rect 231578 179432 231584 179444
rect 132460 179404 231584 179432
rect 132460 179392 132466 179404
rect 231578 179392 231584 179404
rect 231636 179392 231642 179444
rect 180242 179324 180248 179376
rect 180300 179364 180306 179376
rect 258074 179364 258080 179376
rect 180300 179336 258080 179364
rect 180300 179324 180306 179336
rect 258074 179324 258080 179336
rect 258132 179324 258138 179376
rect 574738 179324 574744 179376
rect 574796 179364 574802 179376
rect 580166 179364 580172 179376
rect 574796 179336 580172 179364
rect 574796 179324 574802 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 292022 178712 292028 178764
rect 292080 178752 292086 178764
rect 301406 178752 301412 178764
rect 292080 178724 301412 178752
rect 292080 178712 292086 178724
rect 301406 178712 301412 178724
rect 301464 178712 301470 178764
rect 253198 178644 253204 178696
rect 253256 178684 253262 178696
rect 273438 178684 273444 178696
rect 253256 178656 273444 178684
rect 253256 178644 253262 178656
rect 273438 178644 273444 178656
rect 273496 178644 273502 178696
rect 301498 178644 301504 178696
rect 301556 178684 301562 178696
rect 319070 178684 319076 178696
rect 301556 178656 319076 178684
rect 301556 178644 301562 178656
rect 319070 178644 319076 178656
rect 319128 178644 319134 178696
rect 124490 178100 124496 178152
rect 124548 178140 124554 178152
rect 164970 178140 164976 178152
rect 124548 178112 164976 178140
rect 124548 178100 124554 178112
rect 164970 178100 164976 178112
rect 165028 178100 165034 178152
rect 115842 178032 115848 178084
rect 115900 178072 115906 178084
rect 173434 178072 173440 178084
rect 115900 178044 173440 178072
rect 115900 178032 115906 178044
rect 173434 178032 173440 178044
rect 173492 178032 173498 178084
rect 259730 178032 259736 178084
rect 259788 178072 259794 178084
rect 270494 178072 270500 178084
rect 259788 178044 270500 178072
rect 259788 178032 259794 178044
rect 270494 178032 270500 178044
rect 270552 178032 270558 178084
rect 227714 177964 227720 178016
rect 227772 178004 227778 178016
rect 237374 178004 237380 178016
rect 227772 177976 237380 178004
rect 227772 177964 227778 177976
rect 237374 177964 237380 177976
rect 237432 177964 237438 178016
rect 127618 177692 127624 177744
rect 127676 177732 127682 177744
rect 132494 177732 132500 177744
rect 127676 177704 132500 177732
rect 127676 177692 127682 177704
rect 132494 177692 132500 177704
rect 132552 177692 132558 177744
rect 257338 177352 257344 177404
rect 257396 177392 257402 177404
rect 264974 177392 264980 177404
rect 257396 177364 264980 177392
rect 257396 177352 257402 177364
rect 264974 177352 264980 177364
rect 265032 177352 265038 177404
rect 305270 177352 305276 177404
rect 305328 177392 305334 177404
rect 311894 177392 311900 177404
rect 305328 177364 311900 177392
rect 305328 177352 305334 177364
rect 311894 177352 311900 177364
rect 311952 177352 311958 177404
rect 250622 177284 250628 177336
rect 250680 177324 250686 177336
rect 264238 177324 264244 177336
rect 250680 177296 264244 177324
rect 250680 177284 250686 177296
rect 264238 177284 264244 177296
rect 264296 177284 264302 177336
rect 264330 177284 264336 177336
rect 264388 177324 264394 177336
rect 272150 177324 272156 177336
rect 264388 177296 272156 177324
rect 264388 177284 264394 177296
rect 272150 177284 272156 177296
rect 272208 177284 272214 177336
rect 282178 177284 282184 177336
rect 282236 177324 282242 177336
rect 302418 177324 302424 177336
rect 282236 177296 302424 177324
rect 282236 177284 282242 177296
rect 302418 177284 302424 177296
rect 302476 177284 302482 177336
rect 307018 177284 307024 177336
rect 307076 177324 307082 177336
rect 316310 177324 316316 177336
rect 307076 177296 316316 177324
rect 307076 177284 307082 177296
rect 316310 177284 316316 177296
rect 316368 177284 316374 177336
rect 102042 176876 102048 176928
rect 102100 176916 102106 176928
rect 105446 176916 105452 176928
rect 102100 176888 105452 176916
rect 102100 176876 102106 176888
rect 105446 176876 105452 176888
rect 105504 176876 105510 176928
rect 298738 176876 298744 176928
rect 298796 176916 298802 176928
rect 305270 176916 305276 176928
rect 298796 176888 305276 176916
rect 298796 176876 298802 176888
rect 305270 176876 305276 176888
rect 305328 176876 305334 176928
rect 134426 176740 134432 176792
rect 134484 176780 134490 176792
rect 143442 176780 143448 176792
rect 134484 176752 143448 176780
rect 134484 176740 134490 176752
rect 143442 176740 143448 176752
rect 143500 176740 143506 176792
rect 158990 176740 158996 176792
rect 159048 176780 159054 176792
rect 178862 176780 178868 176792
rect 159048 176752 178868 176780
rect 159048 176740 159054 176752
rect 178862 176740 178868 176752
rect 178920 176740 178926 176792
rect 136082 176672 136088 176724
rect 136140 176712 136146 176724
rect 136140 176684 215340 176712
rect 136140 176672 136146 176684
rect 215312 176644 215340 176684
rect 249518 176644 249524 176656
rect 215312 176616 249524 176644
rect 249518 176604 249524 176616
rect 249576 176604 249582 176656
rect 264422 176604 264428 176656
rect 264480 176644 264486 176656
rect 269206 176644 269212 176656
rect 264480 176616 269212 176644
rect 264480 176604 264486 176616
rect 269206 176604 269212 176616
rect 269264 176604 269270 176656
rect 262950 176536 262956 176588
rect 263008 176576 263014 176588
rect 269114 176576 269120 176588
rect 263008 176548 269120 176576
rect 263008 176536 263014 176548
rect 269114 176536 269120 176548
rect 269172 176536 269178 176588
rect 300210 176536 300216 176588
rect 300268 176576 300274 176588
rect 306558 176576 306564 176588
rect 300268 176548 306564 176576
rect 300268 176536 300274 176548
rect 306558 176536 306564 176548
rect 306616 176536 306622 176588
rect 255958 176196 255964 176248
rect 256016 176236 256022 176248
rect 262214 176236 262220 176248
rect 256016 176208 262220 176236
rect 256016 176196 256022 176208
rect 262214 176196 262220 176208
rect 262272 176196 262278 176248
rect 300118 176196 300124 176248
rect 300176 176236 300182 176248
rect 301130 176236 301136 176248
rect 300176 176208 301136 176236
rect 300176 176196 300182 176208
rect 301130 176196 301136 176208
rect 301188 176196 301194 176248
rect 130746 175992 130752 176044
rect 130804 176032 130810 176044
rect 165522 176032 165528 176044
rect 130804 176004 165528 176032
rect 130804 175992 130810 176004
rect 165522 175992 165528 176004
rect 165580 175992 165586 176044
rect 187050 175992 187056 176044
rect 187108 176032 187114 176044
rect 204898 176032 204904 176044
rect 187108 176004 204904 176032
rect 187108 175992 187114 176004
rect 204898 175992 204904 176004
rect 204956 175992 204962 176044
rect 123110 175924 123116 175976
rect 123168 175964 123174 175976
rect 249242 175964 249248 175976
rect 123168 175936 249248 175964
rect 123168 175924 123174 175936
rect 249242 175924 249248 175936
rect 249300 175924 249306 175976
rect 298186 175788 298192 175840
rect 298244 175788 298250 175840
rect 249702 175312 249708 175364
rect 249760 175352 249766 175364
rect 264422 175352 264428 175364
rect 249760 175324 264428 175352
rect 249760 175312 249766 175324
rect 264422 175312 264428 175324
rect 264480 175312 264486 175364
rect 143442 175176 143448 175228
rect 143500 175216 143506 175228
rect 249702 175216 249708 175228
rect 143500 175188 249708 175216
rect 143500 175176 143506 175188
rect 249702 175176 249708 175188
rect 249760 175176 249766 175228
rect 298204 175216 298232 175788
rect 298204 175188 301452 175216
rect 301424 175160 301452 175188
rect 185670 175108 185676 175160
rect 185728 175148 185734 175160
rect 264330 175148 264336 175160
rect 185728 175120 249794 175148
rect 185728 175108 185734 175120
rect 249766 175080 249794 175120
rect 259426 175120 264336 175148
rect 259426 175080 259454 175120
rect 264330 175108 264336 175120
rect 264388 175108 264394 175160
rect 301406 175108 301412 175160
rect 301464 175108 301470 175160
rect 249766 175052 259454 175080
rect 283742 174020 283748 174072
rect 283800 174060 283806 174072
rect 287790 174060 287796 174072
rect 283800 174032 287796 174060
rect 283800 174020 283806 174032
rect 287790 174020 287796 174032
rect 287848 174020 287854 174072
rect 276658 173884 276664 173936
rect 276716 173924 276722 173936
rect 288342 173924 288348 173936
rect 276716 173896 288348 173924
rect 276716 173884 276722 173896
rect 288342 173884 288348 173896
rect 288400 173884 288406 173936
rect 165522 173816 165528 173868
rect 165580 173856 165586 173868
rect 248598 173856 248604 173868
rect 165580 173828 248604 173856
rect 165580 173816 165586 173828
rect 248598 173816 248604 173828
rect 248656 173816 248662 173868
rect 266630 173816 266636 173868
rect 266688 173856 266694 173868
rect 280246 173856 280252 173868
rect 266688 173828 280252 173856
rect 266688 173816 266694 173828
rect 280246 173816 280252 173828
rect 280304 173816 280310 173868
rect 231578 173748 231584 173800
rect 231636 173788 231642 173800
rect 249702 173788 249708 173800
rect 231636 173760 249708 173788
rect 231636 173748 231642 173760
rect 249702 173748 249708 173760
rect 249760 173748 249766 173800
rect 266354 173748 266360 173800
rect 266412 173788 266418 173800
rect 271966 173788 271972 173800
rect 266412 173760 271972 173788
rect 266412 173748 266418 173760
rect 271966 173748 271972 173760
rect 272024 173748 272030 173800
rect 287790 173340 287796 173392
rect 287848 173380 287854 173392
rect 287974 173380 287980 173392
rect 287848 173352 287980 173380
rect 287848 173340 287854 173352
rect 287974 173340 287980 173352
rect 288032 173340 288038 173392
rect 282270 172592 282276 172644
rect 282328 172632 282334 172644
rect 287606 172632 287612 172644
rect 282328 172604 287612 172632
rect 282328 172592 282334 172604
rect 287606 172592 287612 172604
rect 287664 172592 287670 172644
rect 273898 172524 273904 172576
rect 273956 172564 273962 172576
rect 288342 172564 288348 172576
rect 273956 172536 288348 172564
rect 273956 172524 273962 172536
rect 288342 172524 288348 172536
rect 288400 172524 288406 172576
rect 168466 172456 168472 172508
rect 168524 172496 168530 172508
rect 248598 172496 248604 172508
rect 168524 172468 248604 172496
rect 168524 172456 168530 172468
rect 248598 172456 248604 172468
rect 248656 172456 248662 172508
rect 266630 172456 266636 172508
rect 266688 172496 266694 172508
rect 273346 172496 273352 172508
rect 266688 172468 273352 172496
rect 266688 172456 266694 172468
rect 273346 172456 273352 172468
rect 273404 172456 273410 172508
rect 303890 172456 303896 172508
rect 303948 172496 303954 172508
rect 316218 172496 316224 172508
rect 303948 172468 316224 172496
rect 303948 172456 303954 172468
rect 316218 172456 316224 172468
rect 316276 172456 316282 172508
rect 233970 172388 233976 172440
rect 234028 172428 234034 172440
rect 249334 172428 249340 172440
rect 234028 172400 249340 172428
rect 234028 172388 234034 172400
rect 249334 172388 249340 172400
rect 249392 172388 249398 172440
rect 266354 172388 266360 172440
rect 266412 172428 266418 172440
rect 269114 172428 269120 172440
rect 266412 172400 269120 172428
rect 266412 172388 266418 172400
rect 269114 172388 269120 172400
rect 269172 172388 269178 172440
rect 280890 171164 280896 171216
rect 280948 171204 280954 171216
rect 288342 171204 288348 171216
rect 280948 171176 288348 171204
rect 280948 171164 280954 171176
rect 288342 171164 288348 171176
rect 288400 171164 288406 171216
rect 278314 171096 278320 171148
rect 278372 171136 278378 171148
rect 288250 171136 288256 171148
rect 278372 171108 288256 171136
rect 278372 171096 278378 171108
rect 288250 171096 288256 171108
rect 288308 171096 288314 171148
rect 166442 171028 166448 171080
rect 166500 171068 166506 171080
rect 249610 171068 249616 171080
rect 166500 171040 249616 171068
rect 166500 171028 166506 171040
rect 249610 171028 249616 171040
rect 249668 171028 249674 171080
rect 266722 171028 266728 171080
rect 266780 171068 266786 171080
rect 280154 171068 280160 171080
rect 266780 171040 280160 171068
rect 266780 171028 266786 171040
rect 280154 171028 280160 171040
rect 280212 171028 280218 171080
rect 169110 170960 169116 171012
rect 169168 171000 169174 171012
rect 249702 171000 249708 171012
rect 169168 170972 249708 171000
rect 169168 170960 169174 170972
rect 249702 170960 249708 170972
rect 249760 170960 249766 171012
rect 266354 170960 266360 171012
rect 266412 171000 266418 171012
rect 270494 171000 270500 171012
rect 266412 170972 270500 171000
rect 266412 170960 266418 170972
rect 270494 170960 270500 170972
rect 270552 170960 270558 171012
rect 279602 169736 279608 169788
rect 279660 169776 279666 169788
rect 288342 169776 288348 169788
rect 279660 169748 288348 169776
rect 279660 169736 279666 169748
rect 288342 169736 288348 169748
rect 288400 169736 288406 169788
rect 164970 169668 164976 169720
rect 165028 169708 165034 169720
rect 249702 169708 249708 169720
rect 165028 169680 249708 169708
rect 165028 169668 165034 169680
rect 249702 169668 249708 169680
rect 249760 169668 249766 169720
rect 266354 169668 266360 169720
rect 266412 169708 266418 169720
rect 270770 169708 270776 169720
rect 266412 169680 270776 169708
rect 266412 169668 266418 169680
rect 270770 169668 270776 169680
rect 270828 169668 270834 169720
rect 303890 169668 303896 169720
rect 303948 169708 303954 169720
rect 311894 169708 311900 169720
rect 303948 169680 311900 169708
rect 303948 169668 303954 169680
rect 311894 169668 311900 169680
rect 311952 169668 311958 169720
rect 217318 168988 217324 169040
rect 217376 169028 217382 169040
rect 249150 169028 249156 169040
rect 217376 169000 249156 169028
rect 217376 168988 217382 169000
rect 249150 168988 249156 169000
rect 249208 168988 249214 169040
rect 266354 168988 266360 169040
rect 266412 169028 266418 169040
rect 269298 169028 269304 169040
rect 266412 169000 269304 169028
rect 266412 168988 266418 169000
rect 269298 168988 269304 169000
rect 269356 168988 269362 169040
rect 269942 168988 269948 169040
rect 270000 169028 270006 169040
rect 287238 169028 287244 169040
rect 270000 169000 287244 169028
rect 270000 168988 270006 169000
rect 287238 168988 287244 169000
rect 287296 168988 287302 169040
rect 271414 168376 271420 168428
rect 271472 168416 271478 168428
rect 288158 168416 288164 168428
rect 271472 168388 288164 168416
rect 271472 168376 271478 168388
rect 288158 168376 288164 168388
rect 288216 168376 288222 168428
rect 167914 168308 167920 168360
rect 167972 168348 167978 168360
rect 249610 168348 249616 168360
rect 167972 168320 249616 168348
rect 167972 168308 167978 168320
rect 249610 168308 249616 168320
rect 249668 168308 249674 168360
rect 303890 168308 303896 168360
rect 303948 168348 303954 168360
rect 320450 168348 320456 168360
rect 303948 168320 320456 168348
rect 303948 168308 303954 168320
rect 320450 168308 320456 168320
rect 320508 168308 320514 168360
rect 185762 168240 185768 168292
rect 185820 168280 185826 168292
rect 249702 168280 249708 168292
rect 185820 168252 249708 168280
rect 185820 168240 185826 168252
rect 249702 168240 249708 168252
rect 249760 168240 249766 168292
rect 266354 167968 266360 168020
rect 266412 168008 266418 168020
rect 268010 168008 268016 168020
rect 266412 167980 268016 168008
rect 266412 167968 266418 167980
rect 268010 167968 268016 167980
rect 268068 167968 268074 168020
rect 268654 167084 268660 167136
rect 268712 167124 268718 167136
rect 276014 167124 276020 167136
rect 268712 167096 276020 167124
rect 268712 167084 268718 167096
rect 276014 167084 276020 167096
rect 276072 167084 276078 167136
rect 280798 167084 280804 167136
rect 280856 167124 280862 167136
rect 287974 167124 287980 167136
rect 280856 167096 287980 167124
rect 280856 167084 280862 167096
rect 287974 167084 287980 167096
rect 288032 167084 288038 167136
rect 272610 167016 272616 167068
rect 272668 167056 272674 167068
rect 288342 167056 288348 167068
rect 272668 167028 288348 167056
rect 272668 167016 272674 167028
rect 288342 167016 288348 167028
rect 288400 167016 288406 167068
rect 164878 166948 164884 167000
rect 164936 166988 164942 167000
rect 248414 166988 248420 167000
rect 164936 166960 248420 166988
rect 164936 166948 164942 166960
rect 248414 166948 248420 166960
rect 248472 166948 248478 167000
rect 303890 166948 303896 167000
rect 303948 166988 303954 167000
rect 310790 166988 310796 167000
rect 303948 166960 310796 166988
rect 303948 166948 303954 166960
rect 310790 166948 310796 166960
rect 310848 166948 310854 167000
rect 522298 166948 522304 167000
rect 522356 166988 522362 167000
rect 580166 166988 580172 167000
rect 522356 166960 580172 166988
rect 522356 166948 522362 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 184382 166880 184388 166932
rect 184440 166920 184446 166932
rect 248506 166920 248512 166932
rect 184440 166892 248512 166920
rect 184440 166880 184446 166892
rect 248506 166880 248512 166892
rect 248564 166880 248570 166932
rect 266354 166336 266360 166388
rect 266412 166376 266418 166388
rect 269390 166376 269396 166388
rect 266412 166348 269396 166376
rect 266412 166336 266418 166348
rect 269390 166336 269396 166348
rect 269448 166336 269454 166388
rect 268562 166268 268568 166320
rect 268620 166308 268626 166320
rect 287882 166308 287888 166320
rect 268620 166280 287888 166308
rect 268620 166268 268626 166280
rect 287882 166268 287888 166280
rect 287940 166268 287946 166320
rect 304258 166268 304264 166320
rect 304316 166308 304322 166320
rect 323210 166308 323216 166320
rect 304316 166280 323216 166308
rect 304316 166268 304322 166280
rect 323210 166268 323216 166280
rect 323268 166268 323274 166320
rect 283650 165588 283656 165640
rect 283708 165628 283714 165640
rect 288342 165628 288348 165640
rect 283708 165600 288348 165628
rect 283708 165588 283714 165600
rect 288342 165588 288348 165600
rect 288400 165588 288406 165640
rect 173434 165520 173440 165572
rect 173492 165560 173498 165572
rect 248414 165560 248420 165572
rect 173492 165532 248420 165560
rect 173492 165520 173498 165532
rect 248414 165520 248420 165532
rect 248472 165520 248478 165572
rect 264146 165520 264152 165572
rect 264204 165560 264210 165572
rect 264974 165560 264980 165572
rect 264204 165532 264980 165560
rect 264204 165520 264210 165532
rect 264974 165520 264980 165532
rect 265032 165520 265038 165572
rect 266354 165520 266360 165572
rect 266412 165560 266418 165572
rect 272058 165560 272064 165572
rect 266412 165532 272064 165560
rect 266412 165520 266418 165532
rect 272058 165520 272064 165532
rect 272116 165520 272122 165572
rect 303890 165520 303896 165572
rect 303948 165560 303954 165572
rect 309410 165560 309416 165572
rect 303948 165532 309416 165560
rect 303948 165520 303954 165532
rect 309410 165520 309416 165532
rect 309468 165520 309474 165572
rect 278130 165112 278136 165164
rect 278188 165152 278194 165164
rect 281626 165152 281632 165164
rect 278188 165124 281632 165152
rect 278188 165112 278194 165124
rect 281626 165112 281632 165124
rect 281684 165112 281690 165164
rect 271322 164840 271328 164892
rect 271380 164880 271386 164892
rect 288250 164880 288256 164892
rect 271380 164852 288256 164880
rect 271380 164840 271386 164852
rect 288250 164840 288256 164852
rect 288308 164840 288314 164892
rect 282546 164432 282552 164484
rect 282604 164472 282610 164484
rect 288710 164472 288716 164484
rect 282604 164444 288716 164472
rect 282604 164432 282610 164444
rect 288710 164432 288716 164444
rect 288768 164432 288774 164484
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 33778 164200 33784 164212
rect 3292 164172 33784 164200
rect 3292 164160 3298 164172
rect 33778 164160 33784 164172
rect 33836 164160 33842 164212
rect 182910 164160 182916 164212
rect 182968 164200 182974 164212
rect 248506 164200 248512 164212
rect 182968 164172 248512 164200
rect 182968 164160 182974 164172
rect 248506 164160 248512 164172
rect 248564 164160 248570 164212
rect 266354 164160 266360 164212
rect 266412 164200 266418 164212
rect 277394 164200 277400 164212
rect 266412 164172 277400 164200
rect 266412 164160 266418 164172
rect 277394 164160 277400 164172
rect 277452 164160 277458 164212
rect 303890 164160 303896 164212
rect 303948 164200 303954 164212
rect 325878 164200 325884 164212
rect 303948 164172 325884 164200
rect 303948 164160 303954 164172
rect 325878 164160 325884 164172
rect 325936 164160 325942 164212
rect 231210 164092 231216 164144
rect 231268 164132 231274 164144
rect 248414 164132 248420 164144
rect 231268 164104 248420 164132
rect 231268 164092 231274 164104
rect 248414 164092 248420 164104
rect 248472 164092 248478 164144
rect 271230 164092 271236 164144
rect 271288 164132 271294 164144
rect 273346 164132 273352 164144
rect 271288 164104 273352 164132
rect 271288 164092 271294 164104
rect 273346 164092 273352 164104
rect 273404 164092 273410 164144
rect 170398 163480 170404 163532
rect 170456 163520 170462 163532
rect 221458 163520 221464 163532
rect 170456 163492 221464 163520
rect 170456 163480 170462 163492
rect 221458 163480 221464 163492
rect 221516 163480 221522 163532
rect 303890 163276 303896 163328
rect 303948 163316 303954 163328
rect 307938 163316 307944 163328
rect 303948 163288 307944 163316
rect 303948 163276 303954 163288
rect 307938 163276 307944 163288
rect 307996 163276 308002 163328
rect 276750 162868 276756 162920
rect 276808 162908 276814 162920
rect 288158 162908 288164 162920
rect 276808 162880 288164 162908
rect 276808 162868 276814 162880
rect 288158 162868 288164 162880
rect 288216 162868 288222 162920
rect 171870 162800 171876 162852
rect 171928 162840 171934 162852
rect 248414 162840 248420 162852
rect 171928 162812 248420 162840
rect 171928 162800 171934 162812
rect 248414 162800 248420 162812
rect 248472 162800 248478 162852
rect 266538 162800 266544 162852
rect 266596 162840 266602 162852
rect 270586 162840 270592 162852
rect 266596 162812 270592 162840
rect 266596 162800 266602 162812
rect 270586 162800 270592 162812
rect 270644 162800 270650 162852
rect 303890 162800 303896 162852
rect 303948 162840 303954 162852
rect 317598 162840 317604 162852
rect 303948 162812 317604 162840
rect 303948 162800 303954 162812
rect 317598 162800 317604 162812
rect 317656 162800 317662 162852
rect 181438 162732 181444 162784
rect 181496 162772 181502 162784
rect 248506 162772 248512 162784
rect 181496 162744 248512 162772
rect 181496 162732 181502 162744
rect 248506 162732 248512 162744
rect 248564 162732 248570 162784
rect 266354 162528 266360 162580
rect 266412 162568 266418 162580
rect 269206 162568 269212 162580
rect 266412 162540 269212 162568
rect 266412 162528 266418 162540
rect 269206 162528 269212 162540
rect 269264 162528 269270 162580
rect 269206 162120 269212 162172
rect 269264 162160 269270 162172
rect 283098 162160 283104 162172
rect 269264 162132 283104 162160
rect 269264 162120 269270 162132
rect 283098 162120 283104 162132
rect 283156 162120 283162 162172
rect 282454 161508 282460 161560
rect 282512 161548 282518 161560
rect 288250 161548 288256 161560
rect 282512 161520 288256 161548
rect 282512 161508 282518 161520
rect 288250 161508 288256 161520
rect 288308 161508 288314 161560
rect 285122 161440 285128 161492
rect 285180 161480 285186 161492
rect 288342 161480 288348 161492
rect 285180 161452 288348 161480
rect 285180 161440 285186 161452
rect 288342 161440 288348 161452
rect 288400 161440 288406 161492
rect 167730 161372 167736 161424
rect 167788 161412 167794 161424
rect 248506 161412 248512 161424
rect 167788 161384 248512 161412
rect 167788 161372 167794 161384
rect 248506 161372 248512 161384
rect 248564 161372 248570 161424
rect 266354 161372 266360 161424
rect 266412 161412 266418 161424
rect 274818 161412 274824 161424
rect 266412 161384 274824 161412
rect 266412 161372 266418 161384
rect 274818 161372 274824 161384
rect 274876 161372 274882 161424
rect 303890 161372 303896 161424
rect 303948 161412 303954 161424
rect 319070 161412 319076 161424
rect 303948 161384 319076 161412
rect 303948 161372 303954 161384
rect 319070 161372 319076 161384
rect 319128 161372 319134 161424
rect 238018 161304 238024 161356
rect 238076 161344 238082 161356
rect 248414 161344 248420 161356
rect 238076 161316 248420 161344
rect 238076 161304 238082 161316
rect 248414 161304 248420 161316
rect 248472 161304 248478 161356
rect 269758 160080 269764 160132
rect 269816 160120 269822 160132
rect 287514 160120 287520 160132
rect 269816 160092 287520 160120
rect 269816 160080 269822 160092
rect 287514 160080 287520 160092
rect 287572 160080 287578 160132
rect 177482 160012 177488 160064
rect 177540 160052 177546 160064
rect 248414 160052 248420 160064
rect 177540 160024 248420 160052
rect 177540 160012 177546 160024
rect 248414 160012 248420 160024
rect 248472 160012 248478 160064
rect 303798 159876 303804 159928
rect 303856 159916 303862 159928
rect 306558 159916 306564 159928
rect 303856 159888 306564 159916
rect 303856 159876 303862 159888
rect 306558 159876 306564 159888
rect 306616 159876 306622 159928
rect 265066 159332 265072 159384
rect 265124 159372 265130 159384
rect 271874 159372 271880 159384
rect 265124 159344 271880 159372
rect 265124 159332 265130 159344
rect 271874 159332 271880 159344
rect 271932 159332 271938 159384
rect 281074 158788 281080 158840
rect 281132 158828 281138 158840
rect 288342 158828 288348 158840
rect 281132 158800 288348 158828
rect 281132 158788 281138 158800
rect 288342 158788 288348 158800
rect 288400 158788 288406 158840
rect 279418 158720 279424 158772
rect 279476 158760 279482 158772
rect 287422 158760 287428 158772
rect 279476 158732 287428 158760
rect 279476 158720 279482 158732
rect 287422 158720 287428 158732
rect 287480 158720 287486 158772
rect 170490 158652 170496 158704
rect 170548 158692 170554 158704
rect 248414 158692 248420 158704
rect 170548 158664 248420 158692
rect 170548 158652 170554 158664
rect 248414 158652 248420 158664
rect 248472 158652 248478 158704
rect 266354 158652 266360 158704
rect 266412 158692 266418 158704
rect 274634 158692 274640 158704
rect 266412 158664 274640 158692
rect 266412 158652 266418 158664
rect 274634 158652 274640 158664
rect 274692 158652 274698 158704
rect 303614 158652 303620 158704
rect 303672 158692 303678 158704
rect 310698 158692 310704 158704
rect 303672 158664 310704 158692
rect 303672 158652 303678 158664
rect 310698 158652 310704 158664
rect 310756 158652 310762 158704
rect 275370 158244 275376 158296
rect 275428 158284 275434 158296
rect 279602 158284 279608 158296
rect 275428 158256 279608 158284
rect 275428 158244 275434 158256
rect 279602 158244 279608 158256
rect 279660 158244 279666 158296
rect 178862 157972 178868 158024
rect 178920 158012 178926 158024
rect 249426 158012 249432 158024
rect 178920 157984 249432 158012
rect 178920 157972 178926 157984
rect 249426 157972 249432 157984
rect 249484 157972 249490 158024
rect 266722 157972 266728 158024
rect 266780 158012 266786 158024
rect 276106 158012 276112 158024
rect 266780 157984 276112 158012
rect 266780 157972 266786 157984
rect 276106 157972 276112 157984
rect 276164 157972 276170 158024
rect 277026 157972 277032 158024
rect 277084 158012 277090 158024
rect 280890 158012 280896 158024
rect 277084 157984 280896 158012
rect 277084 157972 277090 157984
rect 280890 157972 280896 157984
rect 280948 157972 280954 158024
rect 283834 157904 283840 157956
rect 283892 157944 283898 157956
rect 287146 157944 287152 157956
rect 283892 157916 287152 157944
rect 283892 157904 283898 157916
rect 287146 157904 287152 157916
rect 287204 157904 287210 157956
rect 176010 157292 176016 157344
rect 176068 157332 176074 157344
rect 249610 157332 249616 157344
rect 176068 157304 249616 157332
rect 176068 157292 176074 157304
rect 249610 157292 249616 157304
rect 249668 157292 249674 157344
rect 266354 157292 266360 157344
rect 266412 157332 266418 157344
rect 270586 157332 270592 157344
rect 266412 157304 270592 157332
rect 266412 157292 266418 157304
rect 270586 157292 270592 157304
rect 270644 157292 270650 157344
rect 303798 157292 303804 157344
rect 303856 157332 303862 157344
rect 313550 157332 313556 157344
rect 303856 157304 313556 157332
rect 303856 157292 303862 157304
rect 313550 157292 313556 157304
rect 313608 157292 313614 157344
rect 188430 157224 188436 157276
rect 188488 157264 188494 157276
rect 249702 157264 249708 157276
rect 188488 157236 249708 157264
rect 188488 157224 188494 157236
rect 249702 157224 249708 157236
rect 249760 157224 249766 157276
rect 283558 156000 283564 156052
rect 283616 156040 283622 156052
rect 288342 156040 288348 156052
rect 283616 156012 288348 156040
rect 283616 156000 283622 156012
rect 288342 156000 288348 156012
rect 288400 156000 288406 156052
rect 279602 155932 279608 155984
rect 279660 155972 279666 155984
rect 288158 155972 288164 155984
rect 279660 155944 288164 155972
rect 279660 155932 279666 155944
rect 288158 155932 288164 155944
rect 288216 155932 288222 155984
rect 166350 155864 166356 155916
rect 166408 155904 166414 155916
rect 249702 155904 249708 155916
rect 166408 155876 249708 155904
rect 166408 155864 166414 155876
rect 249702 155864 249708 155876
rect 249760 155864 249766 155916
rect 266354 155864 266360 155916
rect 266412 155904 266418 155916
rect 280338 155904 280344 155916
rect 266412 155876 280344 155904
rect 266412 155864 266418 155876
rect 280338 155864 280344 155876
rect 280396 155864 280402 155916
rect 303614 155864 303620 155916
rect 303672 155904 303678 155916
rect 331306 155904 331312 155916
rect 303672 155876 331312 155904
rect 303672 155864 303678 155876
rect 331306 155864 331312 155876
rect 331364 155864 331370 155916
rect 220078 155796 220084 155848
rect 220136 155836 220142 155848
rect 249610 155836 249616 155848
rect 220136 155808 249616 155836
rect 220136 155796 220142 155808
rect 249610 155796 249616 155808
rect 249668 155796 249674 155848
rect 303798 155796 303804 155848
rect 303856 155836 303862 155848
rect 321738 155836 321744 155848
rect 303856 155808 321744 155836
rect 303856 155796 303862 155808
rect 321738 155796 321744 155808
rect 321796 155796 321802 155848
rect 266354 155320 266360 155372
rect 266412 155360 266418 155372
rect 270034 155360 270040 155372
rect 266412 155332 270040 155360
rect 266412 155320 266418 155332
rect 270034 155320 270040 155332
rect 270092 155320 270098 155372
rect 177390 155184 177396 155236
rect 177448 155224 177454 155236
rect 213178 155224 213184 155236
rect 177448 155196 213184 155224
rect 177448 155184 177454 155196
rect 213178 155184 213184 155196
rect 213236 155184 213242 155236
rect 287698 155184 287704 155236
rect 287756 155224 287762 155236
rect 288526 155224 288532 155236
rect 287756 155196 288532 155224
rect 287756 155184 287762 155196
rect 288526 155184 288532 155196
rect 288584 155184 288590 155236
rect 281166 155116 281172 155168
rect 281224 155156 281230 155168
rect 287974 155156 287980 155168
rect 281224 155128 287980 155156
rect 281224 155116 281230 155128
rect 287974 155116 287980 155128
rect 288032 155116 288038 155168
rect 269850 154572 269856 154624
rect 269908 154612 269914 154624
rect 288342 154612 288348 154624
rect 269908 154584 288348 154612
rect 269908 154572 269914 154584
rect 288342 154572 288348 154584
rect 288400 154572 288406 154624
rect 303798 154504 303804 154556
rect 303856 154544 303862 154556
rect 335538 154544 335544 154556
rect 303856 154516 335544 154544
rect 303856 154504 303862 154516
rect 335538 154504 335544 154516
rect 335596 154504 335602 154556
rect 303614 154436 303620 154488
rect 303672 154476 303678 154488
rect 332686 154476 332692 154488
rect 303672 154448 332692 154476
rect 303672 154436 303678 154448
rect 332686 154436 332692 154448
rect 332744 154436 332750 154488
rect 265710 153892 265716 153944
rect 265768 153932 265774 153944
rect 283650 153932 283656 153944
rect 265768 153904 283656 153932
rect 265768 153892 265774 153904
rect 283650 153892 283656 153904
rect 283708 153892 283714 153944
rect 268470 153824 268476 153876
rect 268528 153864 268534 153876
rect 287882 153864 287888 153876
rect 268528 153836 287888 153864
rect 268528 153824 268534 153836
rect 287882 153824 287888 153836
rect 287940 153824 287946 153876
rect 266354 153348 266360 153400
rect 266412 153388 266418 153400
rect 268654 153388 268660 153400
rect 266412 153360 268660 153388
rect 266412 153348 266418 153360
rect 268654 153348 268660 153360
rect 268712 153348 268718 153400
rect 246390 153280 246396 153332
rect 246448 153320 246454 153332
rect 249702 153320 249708 153332
rect 246448 153292 249708 153320
rect 246448 153280 246454 153292
rect 249702 153280 249708 153292
rect 249760 153280 249766 153332
rect 214558 153212 214564 153264
rect 214616 153252 214622 153264
rect 249150 153252 249156 153264
rect 214616 153224 249156 153252
rect 214616 153212 214622 153224
rect 249150 153212 249156 153224
rect 249208 153212 249214 153264
rect 303798 153144 303804 153196
rect 303856 153184 303862 153196
rect 324498 153184 324504 153196
rect 303856 153156 324504 153184
rect 303856 153144 303862 153156
rect 324498 153144 324504 153156
rect 324556 153144 324562 153196
rect 303890 153076 303896 153128
rect 303948 153116 303954 153128
rect 312078 153116 312084 153128
rect 303948 153088 312084 153116
rect 303948 153076 303954 153088
rect 312078 153076 312084 153088
rect 312136 153076 312142 153128
rect 174630 152464 174636 152516
rect 174688 152504 174694 152516
rect 217318 152504 217324 152516
rect 174688 152476 217324 152504
rect 174688 152464 174694 152476
rect 217318 152464 217324 152476
rect 217376 152464 217382 152516
rect 267090 152464 267096 152516
rect 267148 152504 267154 152516
rect 282270 152504 282276 152516
rect 267148 152476 282276 152504
rect 267148 152464 267154 152476
rect 282270 152464 282276 152476
rect 282328 152464 282334 152516
rect 222930 151852 222936 151904
rect 222988 151892 222994 151904
rect 249702 151892 249708 151904
rect 222988 151864 249708 151892
rect 222988 151852 222994 151864
rect 249702 151852 249708 151864
rect 249760 151852 249766 151904
rect 283650 151852 283656 151904
rect 283708 151892 283714 151904
rect 288342 151892 288348 151904
rect 283708 151864 288348 151892
rect 283708 151852 283714 151864
rect 288342 151852 288348 151864
rect 288400 151852 288406 151904
rect 214650 151784 214656 151836
rect 214708 151824 214714 151836
rect 248966 151824 248972 151836
rect 214708 151796 248972 151824
rect 214708 151784 214714 151796
rect 248966 151784 248972 151796
rect 249024 151784 249030 151836
rect 266262 151784 266268 151836
rect 266320 151824 266326 151836
rect 288250 151824 288256 151836
rect 266320 151796 288256 151824
rect 266320 151784 266326 151796
rect 288250 151784 288256 151796
rect 288308 151784 288314 151836
rect 266354 151580 266360 151632
rect 266412 151620 266418 151632
rect 269114 151620 269120 151632
rect 266412 151592 269120 151620
rect 266412 151580 266418 151592
rect 269114 151580 269120 151592
rect 269172 151580 269178 151632
rect 169018 151036 169024 151088
rect 169076 151076 169082 151088
rect 248966 151076 248972 151088
rect 169076 151048 248972 151076
rect 169076 151036 169082 151048
rect 248966 151036 248972 151048
rect 249024 151036 249030 151088
rect 278130 150492 278136 150544
rect 278188 150532 278194 150544
rect 288342 150532 288348 150544
rect 278188 150504 288348 150532
rect 278188 150492 278194 150504
rect 288342 150492 288348 150504
rect 288400 150492 288406 150544
rect 178862 150424 178868 150476
rect 178920 150464 178926 150476
rect 249702 150464 249708 150476
rect 178920 150436 249708 150464
rect 178920 150424 178926 150436
rect 249702 150424 249708 150436
rect 249760 150424 249766 150476
rect 275462 150424 275468 150476
rect 275520 150464 275526 150476
rect 287974 150464 287980 150476
rect 275520 150436 287980 150464
rect 275520 150424 275526 150436
rect 287974 150424 287980 150436
rect 288032 150424 288038 150476
rect 3510 150356 3516 150408
rect 3568 150396 3574 150408
rect 14458 150396 14464 150408
rect 3568 150368 14464 150396
rect 3568 150356 3574 150368
rect 14458 150356 14464 150368
rect 14516 150356 14522 150408
rect 167638 150356 167644 150408
rect 167696 150396 167702 150408
rect 249610 150396 249616 150408
rect 167696 150368 249616 150396
rect 167696 150356 167702 150368
rect 249610 150356 249616 150368
rect 249668 150356 249674 150408
rect 266354 150356 266360 150408
rect 266412 150396 266418 150408
rect 278774 150396 278780 150408
rect 266412 150368 278780 150396
rect 266412 150356 266418 150368
rect 278774 150356 278780 150368
rect 278832 150356 278838 150408
rect 303798 150356 303804 150408
rect 303856 150396 303862 150408
rect 316310 150396 316316 150408
rect 303856 150368 316316 150396
rect 303856 150356 303862 150368
rect 316310 150356 316316 150368
rect 316368 150356 316374 150408
rect 180150 149676 180156 149728
rect 180208 149716 180214 149728
rect 249242 149716 249248 149728
rect 180208 149688 249248 149716
rect 180208 149676 180214 149688
rect 249242 149676 249248 149688
rect 249300 149676 249306 149728
rect 280982 149064 280988 149116
rect 281040 149104 281046 149116
rect 288342 149104 288348 149116
rect 281040 149076 288348 149104
rect 281040 149064 281046 149076
rect 288342 149064 288348 149076
rect 288400 149064 288406 149116
rect 303798 148996 303804 149048
rect 303856 149036 303862 149048
rect 320266 149036 320272 149048
rect 303856 149008 320272 149036
rect 303856 148996 303862 149008
rect 320266 148996 320272 149008
rect 320324 148996 320330 149048
rect 267182 148384 267188 148436
rect 267240 148424 267246 148436
rect 279510 148424 279516 148436
rect 267240 148396 279516 148424
rect 267240 148384 267246 148396
rect 279510 148384 279516 148396
rect 279568 148384 279574 148436
rect 181530 148316 181536 148368
rect 181588 148356 181594 148368
rect 226978 148356 226984 148368
rect 181588 148328 226984 148356
rect 181588 148316 181594 148328
rect 226978 148316 226984 148328
rect 227036 148316 227042 148368
rect 270034 148316 270040 148368
rect 270092 148356 270098 148368
rect 284938 148356 284944 148368
rect 270092 148328 284944 148356
rect 270092 148316 270098 148328
rect 284938 148316 284944 148328
rect 284996 148316 285002 148368
rect 279694 147636 279700 147688
rect 279752 147676 279758 147688
rect 288342 147676 288348 147688
rect 279752 147648 288348 147676
rect 279752 147636 279758 147648
rect 288342 147636 288348 147648
rect 288400 147636 288406 147688
rect 266354 147568 266360 147620
rect 266412 147608 266418 147620
rect 275554 147608 275560 147620
rect 266412 147580 275560 147608
rect 266412 147568 266418 147580
rect 275554 147568 275560 147580
rect 275612 147568 275618 147620
rect 303706 147568 303712 147620
rect 303764 147608 303770 147620
rect 327350 147608 327356 147620
rect 303764 147580 327356 147608
rect 303764 147568 303770 147580
rect 327350 147568 327356 147580
rect 327408 147568 327414 147620
rect 276934 146888 276940 146940
rect 276992 146928 276998 146940
rect 287238 146928 287244 146940
rect 276992 146900 287244 146928
rect 276992 146888 276998 146900
rect 287238 146888 287244 146900
rect 287296 146888 287302 146940
rect 246482 146344 246488 146396
rect 246540 146384 246546 146396
rect 249702 146384 249708 146396
rect 246540 146356 249708 146384
rect 246540 146344 246546 146356
rect 249702 146344 249708 146356
rect 249760 146344 249766 146396
rect 177390 146276 177396 146328
rect 177448 146316 177454 146328
rect 249150 146316 249156 146328
rect 177448 146288 249156 146316
rect 177448 146276 177454 146288
rect 249150 146276 249156 146288
rect 249208 146276 249214 146328
rect 264238 146276 264244 146328
rect 264296 146316 264302 146328
rect 288342 146316 288348 146328
rect 264296 146288 288348 146316
rect 264296 146276 264302 146288
rect 288342 146276 288348 146288
rect 288400 146276 288406 146328
rect 303798 146208 303804 146260
rect 303856 146248 303862 146260
rect 317690 146248 317696 146260
rect 303856 146220 317696 146248
rect 303856 146208 303862 146220
rect 317690 146208 317696 146220
rect 317748 146208 317754 146260
rect 303706 145800 303712 145852
rect 303764 145840 303770 145852
rect 308030 145840 308036 145852
rect 303764 145812 308036 145840
rect 303764 145800 303770 145812
rect 308030 145800 308036 145812
rect 308088 145800 308094 145852
rect 274082 145664 274088 145716
rect 274140 145704 274146 145716
rect 277026 145704 277032 145716
rect 274140 145676 277032 145704
rect 274140 145664 274146 145676
rect 277026 145664 277032 145676
rect 277084 145664 277090 145716
rect 197998 145596 198004 145648
rect 198056 145636 198062 145648
rect 218790 145636 218796 145648
rect 198056 145608 218796 145636
rect 198056 145596 198062 145608
rect 218790 145596 218796 145608
rect 218848 145596 218854 145648
rect 171778 145528 171784 145580
rect 171836 145568 171842 145580
rect 204990 145568 204996 145580
rect 171836 145540 204996 145568
rect 171836 145528 171842 145540
rect 204990 145528 204996 145540
rect 205048 145528 205054 145580
rect 231210 144916 231216 144968
rect 231268 144956 231274 144968
rect 249702 144956 249708 144968
rect 231268 144928 249708 144956
rect 231268 144916 231274 144928
rect 249702 144916 249708 144928
rect 249760 144916 249766 144968
rect 284938 144916 284944 144968
rect 284996 144956 285002 144968
rect 287422 144956 287428 144968
rect 284996 144928 287428 144956
rect 284996 144916 285002 144928
rect 287422 144916 287428 144928
rect 287480 144916 287486 144968
rect 266354 144848 266360 144900
rect 266412 144888 266418 144900
rect 271230 144888 271236 144900
rect 266412 144860 271236 144888
rect 266412 144848 266418 144860
rect 271230 144848 271236 144860
rect 271288 144848 271294 144900
rect 303798 144848 303804 144900
rect 303856 144888 303862 144900
rect 323118 144888 323124 144900
rect 303856 144860 323124 144888
rect 303856 144848 303862 144860
rect 323118 144848 323124 144860
rect 323176 144848 323182 144900
rect 275554 144168 275560 144220
rect 275612 144208 275618 144220
rect 287790 144208 287796 144220
rect 275612 144180 287796 144208
rect 275612 144168 275618 144180
rect 287790 144168 287796 144180
rect 287848 144168 287854 144220
rect 303982 144168 303988 144220
rect 304040 144208 304046 144220
rect 316126 144208 316132 144220
rect 304040 144180 316132 144208
rect 304040 144168 304046 144180
rect 316126 144168 316132 144180
rect 316184 144168 316190 144220
rect 238018 143624 238024 143676
rect 238076 143664 238082 143676
rect 249702 143664 249708 143676
rect 238076 143636 249708 143664
rect 238076 143624 238082 143636
rect 249702 143624 249708 143636
rect 249760 143624 249766 143676
rect 196710 143556 196716 143608
rect 196768 143596 196774 143608
rect 249150 143596 249156 143608
rect 196768 143568 249156 143596
rect 196768 143556 196774 143568
rect 249150 143556 249156 143568
rect 249208 143556 249214 143608
rect 265618 143556 265624 143608
rect 265676 143596 265682 143608
rect 288158 143596 288164 143608
rect 265676 143568 288164 143596
rect 265676 143556 265682 143568
rect 288158 143556 288164 143568
rect 288216 143556 288222 143608
rect 266354 143488 266360 143540
rect 266412 143528 266418 143540
rect 273254 143528 273260 143540
rect 266412 143500 273260 143528
rect 266412 143488 266418 143500
rect 273254 143488 273260 143500
rect 273312 143488 273318 143540
rect 175918 142808 175924 142860
rect 175976 142848 175982 142860
rect 249610 142848 249616 142860
rect 175976 142820 249616 142848
rect 175976 142808 175982 142820
rect 249610 142808 249616 142820
rect 249668 142808 249674 142860
rect 274174 142808 274180 142860
rect 274232 142848 274238 142860
rect 287882 142848 287888 142860
rect 274232 142820 287888 142848
rect 274232 142808 274238 142820
rect 287882 142808 287888 142820
rect 287940 142808 287946 142860
rect 242250 142128 242256 142180
rect 242308 142168 242314 142180
rect 249702 142168 249708 142180
rect 242308 142140 249708 142168
rect 242308 142128 242314 142140
rect 249702 142128 249708 142140
rect 249760 142128 249766 142180
rect 272794 142128 272800 142180
rect 272852 142168 272858 142180
rect 279602 142168 279608 142180
rect 272852 142140 279608 142168
rect 272852 142128 272858 142140
rect 279602 142128 279608 142140
rect 279660 142128 279666 142180
rect 282362 142128 282368 142180
rect 282420 142168 282426 142180
rect 287974 142168 287980 142180
rect 282420 142140 287980 142168
rect 282420 142128 282426 142140
rect 287974 142128 287980 142140
rect 288032 142128 288038 142180
rect 303798 142060 303804 142112
rect 303856 142100 303862 142112
rect 322934 142100 322940 142112
rect 303856 142072 322940 142100
rect 303856 142060 303862 142072
rect 322934 142060 322940 142072
rect 322992 142060 322998 142112
rect 191098 141448 191104 141500
rect 191156 141488 191162 141500
rect 209038 141488 209044 141500
rect 191156 141460 209044 141488
rect 191156 141448 191162 141460
rect 209038 141448 209044 141460
rect 209096 141448 209102 141500
rect 271230 141448 271236 141500
rect 271288 141488 271294 141500
rect 288250 141488 288256 141500
rect 271288 141460 288256 141488
rect 271288 141448 271294 141460
rect 288250 141448 288256 141460
rect 288308 141448 288314 141500
rect 178770 141380 178776 141432
rect 178828 141420 178834 141432
rect 199378 141420 199384 141432
rect 178828 141392 199384 141420
rect 178828 141380 178834 141392
rect 199378 141380 199384 141392
rect 199436 141380 199442 141432
rect 266446 141380 266452 141432
rect 266504 141420 266510 141432
rect 285214 141420 285220 141432
rect 266504 141392 285220 141420
rect 266504 141380 266510 141392
rect 285214 141380 285220 141392
rect 285272 141380 285278 141432
rect 229830 140836 229836 140888
rect 229888 140876 229894 140888
rect 249610 140876 249616 140888
rect 229888 140848 249616 140876
rect 229888 140836 229894 140848
rect 249610 140836 249616 140848
rect 249668 140836 249674 140888
rect 224218 140768 224224 140820
rect 224276 140808 224282 140820
rect 249702 140808 249708 140820
rect 224276 140780 249708 140808
rect 224276 140768 224282 140780
rect 249702 140768 249708 140780
rect 249760 140768 249766 140820
rect 284294 139816 284300 139868
rect 284352 139856 284358 139868
rect 288066 139856 288072 139868
rect 284352 139828 288072 139856
rect 284352 139816 284358 139828
rect 288066 139816 288072 139828
rect 288124 139816 288130 139868
rect 303614 139816 303620 139868
rect 303672 139856 303678 139868
rect 305270 139856 305276 139868
rect 303672 139828 305276 139856
rect 303672 139816 303678 139828
rect 305270 139816 305276 139828
rect 305328 139816 305334 139868
rect 232682 139408 232688 139460
rect 232740 139448 232746 139460
rect 249150 139448 249156 139460
rect 232740 139420 249156 139448
rect 232740 139408 232746 139420
rect 249150 139408 249156 139420
rect 249208 139408 249214 139460
rect 266354 139340 266360 139392
rect 266412 139380 266418 139392
rect 267734 139380 267740 139392
rect 266412 139352 267740 139380
rect 266412 139340 266418 139352
rect 267734 139340 267740 139352
rect 267792 139340 267798 139392
rect 303798 139340 303804 139392
rect 303856 139380 303862 139392
rect 314838 139380 314844 139392
rect 303856 139352 314844 139380
rect 303856 139340 303862 139352
rect 314838 139340 314844 139352
rect 314896 139340 314902 139392
rect 264054 138864 264060 138916
rect 264112 138864 264118 138916
rect 173250 138660 173256 138712
rect 173308 138700 173314 138712
rect 198090 138700 198096 138712
rect 173308 138672 198096 138700
rect 173308 138660 173314 138672
rect 198090 138660 198096 138672
rect 198148 138660 198154 138712
rect 233970 138660 233976 138712
rect 234028 138700 234034 138712
rect 249334 138700 249340 138712
rect 234028 138672 249340 138700
rect 234028 138660 234034 138672
rect 249334 138660 249340 138672
rect 249392 138660 249398 138712
rect 264072 138700 264100 138864
rect 280798 138700 280804 138712
rect 264072 138672 280804 138700
rect 280798 138660 280804 138672
rect 280856 138660 280862 138712
rect 280890 138048 280896 138100
rect 280948 138088 280954 138100
rect 288250 138088 288256 138100
rect 280948 138060 288256 138088
rect 280948 138048 280954 138060
rect 288250 138048 288256 138060
rect 288308 138048 288314 138100
rect 181438 137980 181444 138032
rect 181496 138020 181502 138032
rect 249702 138020 249708 138032
rect 181496 137992 249708 138020
rect 181496 137980 181502 137992
rect 249702 137980 249708 137992
rect 249760 137980 249766 138032
rect 268654 137980 268660 138032
rect 268712 138020 268718 138032
rect 269942 138020 269948 138032
rect 268712 137992 269948 138020
rect 268712 137980 268718 137992
rect 269942 137980 269948 137992
rect 270000 137980 270006 138032
rect 279602 137980 279608 138032
rect 279660 138020 279666 138032
rect 288342 138020 288348 138032
rect 279660 137992 288348 138020
rect 279660 137980 279666 137992
rect 288342 137980 288348 137992
rect 288400 137980 288406 138032
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 25498 137952 25504 137964
rect 3568 137924 25504 137952
rect 3568 137912 3574 137924
rect 25498 137912 25504 137924
rect 25556 137912 25562 137964
rect 303798 137912 303804 137964
rect 303856 137952 303862 137964
rect 328546 137952 328552 137964
rect 303856 137924 328552 137952
rect 303856 137912 303862 137924
rect 328546 137912 328552 137924
rect 328604 137912 328610 137964
rect 186958 137300 186964 137352
rect 187016 137340 187022 137352
rect 202138 137340 202144 137352
rect 187016 137312 202144 137340
rect 187016 137300 187022 137312
rect 202138 137300 202144 137312
rect 202196 137300 202202 137352
rect 277118 137300 277124 137352
rect 277176 137340 277182 137352
rect 281166 137340 281172 137352
rect 277176 137312 281172 137340
rect 277176 137300 277182 137312
rect 281166 137300 281172 137312
rect 281224 137300 281230 137352
rect 167730 137232 167736 137284
rect 167788 137272 167794 137284
rect 222930 137272 222936 137284
rect 167788 137244 222936 137272
rect 167788 137232 167794 137244
rect 222930 137232 222936 137244
rect 222988 137232 222994 137284
rect 266354 137232 266360 137284
rect 266412 137272 266418 137284
rect 283742 137272 283748 137284
rect 266412 137244 283748 137272
rect 266412 137232 266418 137244
rect 283742 137232 283748 137244
rect 283800 137232 283806 137284
rect 245010 136688 245016 136740
rect 245068 136728 245074 136740
rect 249150 136728 249156 136740
rect 245068 136700 249156 136728
rect 245068 136688 245074 136700
rect 249150 136688 249156 136700
rect 249208 136688 249214 136740
rect 203610 136620 203616 136672
rect 203668 136660 203674 136672
rect 249702 136660 249708 136672
rect 203668 136632 249708 136660
rect 203668 136620 203674 136632
rect 249702 136620 249708 136632
rect 249760 136620 249766 136672
rect 283834 136620 283840 136672
rect 283892 136660 283898 136672
rect 288342 136660 288348 136672
rect 283892 136632 288348 136660
rect 283892 136620 283898 136632
rect 288342 136620 288348 136632
rect 288400 136620 288406 136672
rect 303614 136552 303620 136604
rect 303672 136592 303678 136604
rect 310606 136592 310612 136604
rect 303672 136564 310612 136592
rect 303672 136552 303678 136564
rect 310606 136552 310612 136564
rect 310664 136552 310670 136604
rect 195330 135872 195336 135924
rect 195388 135912 195394 135924
rect 220078 135912 220084 135924
rect 195388 135884 220084 135912
rect 195388 135872 195394 135884
rect 220078 135872 220084 135884
rect 220136 135872 220142 135924
rect 268746 135872 268752 135924
rect 268804 135912 268810 135924
rect 289170 135912 289176 135924
rect 268804 135884 289176 135912
rect 268804 135872 268810 135884
rect 289170 135872 289176 135884
rect 289228 135872 289234 135924
rect 266354 135600 266360 135652
rect 266412 135640 266418 135652
rect 268562 135640 268568 135652
rect 266412 135612 268568 135640
rect 266412 135600 266418 135612
rect 268562 135600 268568 135612
rect 268620 135600 268626 135652
rect 235258 135328 235264 135380
rect 235316 135368 235322 135380
rect 249702 135368 249708 135380
rect 235316 135340 249708 135368
rect 235316 135328 235322 135340
rect 249702 135328 249708 135340
rect 249760 135328 249766 135380
rect 167638 135260 167644 135312
rect 167696 135300 167702 135312
rect 249150 135300 249156 135312
rect 167696 135272 249156 135300
rect 167696 135260 167702 135272
rect 249150 135260 249156 135272
rect 249208 135260 249214 135312
rect 266354 135192 266360 135244
rect 266412 135232 266418 135244
rect 276658 135232 276664 135244
rect 266412 135204 276664 135232
rect 266412 135192 266418 135204
rect 276658 135192 276664 135204
rect 276716 135192 276722 135244
rect 303706 135192 303712 135244
rect 303764 135232 303770 135244
rect 339586 135232 339592 135244
rect 303764 135204 339592 135232
rect 303764 135192 303770 135204
rect 339586 135192 339592 135204
rect 339644 135192 339650 135244
rect 197998 134512 198004 134564
rect 198056 134552 198062 134564
rect 246482 134552 246488 134564
rect 198056 134524 246488 134552
rect 198056 134512 198062 134524
rect 246482 134512 246488 134524
rect 246540 134512 246546 134564
rect 304718 134512 304724 134564
rect 304776 134552 304782 134564
rect 312170 134552 312176 134564
rect 304776 134524 312176 134552
rect 304776 134512 304782 134524
rect 312170 134512 312176 134524
rect 312228 134512 312234 134564
rect 171778 133900 171784 133952
rect 171836 133940 171842 133952
rect 249702 133940 249708 133952
rect 171836 133912 249708 133940
rect 171836 133900 171842 133912
rect 249702 133900 249708 133912
rect 249760 133900 249766 133952
rect 266354 133832 266360 133884
rect 266412 133872 266418 133884
rect 273898 133872 273904 133884
rect 266412 133844 273904 133872
rect 266412 133832 266418 133844
rect 273898 133832 273904 133844
rect 273956 133832 273962 133884
rect 303890 133832 303896 133884
rect 303948 133872 303954 133884
rect 331398 133872 331404 133884
rect 303948 133844 331404 133872
rect 303948 133832 303954 133844
rect 331398 133832 331404 133844
rect 331456 133832 331462 133884
rect 303798 133764 303804 133816
rect 303856 133804 303862 133816
rect 321646 133804 321652 133816
rect 303856 133776 321652 133804
rect 303856 133764 303862 133776
rect 321646 133764 321652 133776
rect 321704 133764 321710 133816
rect 274266 133220 274272 133272
rect 274324 133260 274330 133272
rect 287422 133260 287428 133272
rect 274324 133232 287428 133260
rect 274324 133220 274330 133232
rect 287422 133220 287428 133232
rect 287480 133220 287486 133272
rect 173342 133152 173348 133204
rect 173400 133192 173406 133204
rect 249242 133192 249248 133204
rect 173400 133164 249248 133192
rect 173400 133152 173406 133164
rect 249242 133152 249248 133164
rect 249300 133152 249306 133204
rect 269942 133152 269948 133204
rect 270000 133192 270006 133204
rect 284294 133192 284300 133204
rect 270000 133164 284300 133192
rect 270000 133152 270006 133164
rect 284294 133152 284300 133164
rect 284352 133152 284358 133204
rect 266354 132948 266360 133000
rect 266412 132988 266418 133000
rect 268654 132988 268660 133000
rect 266412 132960 268660 132988
rect 266412 132948 266418 132960
rect 268654 132948 268660 132960
rect 268712 132948 268718 133000
rect 285214 132472 285220 132524
rect 285272 132512 285278 132524
rect 288342 132512 288348 132524
rect 285272 132484 288348 132512
rect 285272 132472 285278 132484
rect 288342 132472 288348 132484
rect 288400 132472 288406 132524
rect 266446 132404 266452 132456
rect 266504 132444 266510 132456
rect 275370 132444 275376 132456
rect 266504 132416 275376 132444
rect 266504 132404 266510 132416
rect 275370 132404 275376 132416
rect 275428 132404 275434 132456
rect 303798 132404 303804 132456
rect 303856 132444 303862 132456
rect 327166 132444 327172 132456
rect 303856 132416 327172 132444
rect 303856 132404 303862 132416
rect 327166 132404 327172 132416
rect 327224 132404 327230 132456
rect 266354 132336 266360 132388
rect 266412 132376 266418 132388
rect 274082 132376 274088 132388
rect 266412 132348 274088 132376
rect 266412 132336 266418 132348
rect 274082 132336 274088 132348
rect 274140 132336 274146 132388
rect 303890 132336 303896 132388
rect 303948 132376 303954 132388
rect 317506 132376 317512 132388
rect 303948 132348 317512 132376
rect 303948 132336 303954 132348
rect 317506 132336 317512 132348
rect 317564 132336 317570 132388
rect 176010 131724 176016 131776
rect 176068 131764 176074 131776
rect 246390 131764 246396 131776
rect 176068 131736 246396 131764
rect 176068 131724 176074 131736
rect 246390 131724 246396 131736
rect 246448 131724 246454 131776
rect 173250 131112 173256 131164
rect 173308 131152 173314 131164
rect 249702 131152 249708 131164
rect 173308 131124 249708 131152
rect 173308 131112 173314 131124
rect 249702 131112 249708 131124
rect 249760 131112 249766 131164
rect 274542 131112 274548 131164
rect 274600 131152 274606 131164
rect 288342 131152 288348 131164
rect 274600 131124 288348 131152
rect 274600 131112 274606 131124
rect 288342 131112 288348 131124
rect 288400 131112 288406 131164
rect 266446 131044 266452 131096
rect 266504 131084 266510 131096
rect 271414 131084 271420 131096
rect 266504 131056 271420 131084
rect 266504 131044 266510 131056
rect 271414 131044 271420 131056
rect 271472 131044 271478 131096
rect 303798 131044 303804 131096
rect 303856 131084 303862 131096
rect 329926 131084 329932 131096
rect 303856 131056 329932 131084
rect 303856 131044 303862 131056
rect 329926 131044 329932 131056
rect 329984 131044 329990 131096
rect 266538 130908 266544 130960
rect 266596 130948 266602 130960
rect 270034 130948 270040 130960
rect 266596 130920 270040 130948
rect 266596 130908 266602 130920
rect 270034 130908 270040 130920
rect 270092 130908 270098 130960
rect 278314 130364 278320 130416
rect 278372 130404 278378 130416
rect 289262 130404 289268 130416
rect 278372 130376 289268 130404
rect 278372 130364 278378 130376
rect 289262 130364 289268 130376
rect 289320 130364 289326 130416
rect 304258 130364 304264 130416
rect 304316 130404 304322 130416
rect 318978 130404 318984 130416
rect 304316 130376 318984 130404
rect 304316 130364 304322 130376
rect 318978 130364 318984 130376
rect 319036 130364 319042 130416
rect 213270 129820 213276 129872
rect 213328 129860 213334 129872
rect 249610 129860 249616 129872
rect 213328 129832 249616 129860
rect 213328 129820 213334 129832
rect 249610 129820 249616 129832
rect 249668 129820 249674 129872
rect 211890 129752 211896 129804
rect 211948 129792 211954 129804
rect 249702 129792 249708 129804
rect 211948 129764 249708 129792
rect 211948 129752 211954 129764
rect 249702 129752 249708 129764
rect 249760 129752 249766 129804
rect 277026 129752 277032 129804
rect 277084 129792 277090 129804
rect 288342 129792 288348 129804
rect 277084 129764 288348 129792
rect 277084 129752 277090 129764
rect 288342 129752 288348 129764
rect 288400 129752 288406 129804
rect 266354 129684 266360 129736
rect 266412 129724 266418 129736
rect 276842 129724 276848 129736
rect 266412 129696 276848 129724
rect 266412 129684 266418 129696
rect 276842 129684 276848 129696
rect 276900 129684 276906 129736
rect 303798 129684 303804 129736
rect 303856 129724 303862 129736
rect 314930 129724 314936 129736
rect 303856 129696 314936 129724
rect 303856 129684 303862 129696
rect 314930 129684 314936 129696
rect 314988 129684 314994 129736
rect 267090 129616 267096 129668
rect 267148 129656 267154 129668
rect 269758 129656 269764 129668
rect 267148 129628 269764 129656
rect 267148 129616 267154 129628
rect 269758 129616 269764 129628
rect 269816 129616 269822 129668
rect 270034 129004 270040 129056
rect 270092 129044 270098 129056
rect 287698 129044 287704 129056
rect 270092 129016 287704 129044
rect 270092 129004 270098 129016
rect 287698 129004 287704 129016
rect 287756 129004 287762 129056
rect 195330 128324 195336 128376
rect 195388 128364 195394 128376
rect 249702 128364 249708 128376
rect 195388 128336 249708 128364
rect 195388 128324 195394 128336
rect 249702 128324 249708 128336
rect 249760 128324 249766 128376
rect 276750 128324 276756 128376
rect 276808 128364 276814 128376
rect 287974 128364 287980 128376
rect 276808 128336 287980 128364
rect 276808 128324 276814 128336
rect 287974 128324 287980 128336
rect 288032 128324 288038 128376
rect 303798 128256 303804 128308
rect 303856 128296 303862 128308
rect 336734 128296 336740 128308
rect 303856 128268 336740 128296
rect 303856 128256 303862 128268
rect 336734 128256 336740 128268
rect 336792 128256 336798 128308
rect 303614 128188 303620 128240
rect 303672 128228 303678 128240
rect 313366 128228 313372 128240
rect 303672 128200 313372 128228
rect 303672 128188 303678 128200
rect 313366 128188 313372 128200
rect 313424 128188 313430 128240
rect 266354 127984 266360 128036
rect 266412 128024 266418 128036
rect 268746 128024 268752 128036
rect 266412 127996 268752 128024
rect 266412 127984 266418 127996
rect 268746 127984 268752 127996
rect 268804 127984 268810 128036
rect 264790 127644 264796 127696
rect 264848 127684 264854 127696
rect 266998 127684 267004 127696
rect 264848 127656 267004 127684
rect 264848 127644 264854 127656
rect 266998 127644 267004 127656
rect 267056 127644 267062 127696
rect 266446 127576 266452 127628
rect 266504 127616 266510 127628
rect 273990 127616 273996 127628
rect 266504 127588 273996 127616
rect 266504 127576 266510 127588
rect 273990 127576 273996 127588
rect 274048 127576 274054 127628
rect 268562 127440 268568 127492
rect 268620 127480 268626 127492
rect 272794 127480 272800 127492
rect 268620 127452 272800 127480
rect 268620 127440 268626 127452
rect 272794 127440 272800 127452
rect 272852 127440 272858 127492
rect 229738 127032 229744 127084
rect 229796 127072 229802 127084
rect 249702 127072 249708 127084
rect 229796 127044 249708 127072
rect 229796 127032 229802 127044
rect 249702 127032 249708 127044
rect 249760 127032 249766 127084
rect 188522 126964 188528 127016
rect 188580 127004 188586 127016
rect 249610 127004 249616 127016
rect 188580 126976 249616 127004
rect 188580 126964 188586 126976
rect 249610 126964 249616 126976
rect 249668 126964 249674 127016
rect 283926 126964 283932 127016
rect 283984 127004 283990 127016
rect 287974 127004 287980 127016
rect 283984 126976 287980 127004
rect 283984 126964 283990 126976
rect 287974 126964 287980 126976
rect 288032 126964 288038 127016
rect 266354 126896 266360 126948
rect 266412 126936 266418 126948
rect 271322 126936 271328 126948
rect 266412 126908 271328 126936
rect 266412 126896 266418 126908
rect 271322 126896 271328 126908
rect 271380 126896 271386 126948
rect 184290 126284 184296 126336
rect 184348 126324 184354 126336
rect 196618 126324 196624 126336
rect 184348 126296 196624 126324
rect 184348 126284 184354 126296
rect 196618 126284 196624 126296
rect 196676 126284 196682 126336
rect 178770 126216 178776 126268
rect 178828 126256 178834 126268
rect 214650 126256 214656 126268
rect 178828 126228 214656 126256
rect 178828 126216 178834 126228
rect 214650 126216 214656 126228
rect 214708 126216 214714 126268
rect 266998 126216 267004 126268
rect 267056 126256 267062 126268
rect 277118 126256 277124 126268
rect 267056 126228 277124 126256
rect 267056 126216 267062 126228
rect 277118 126216 277124 126228
rect 277176 126216 277182 126268
rect 220170 125672 220176 125724
rect 220228 125712 220234 125724
rect 249610 125712 249616 125724
rect 220228 125684 249616 125712
rect 220228 125672 220234 125684
rect 249610 125672 249616 125684
rect 249668 125672 249674 125724
rect 280798 125672 280804 125724
rect 280856 125712 280862 125724
rect 288250 125712 288256 125724
rect 280856 125684 288256 125712
rect 280856 125672 280862 125684
rect 288250 125672 288256 125684
rect 288308 125672 288314 125724
rect 200850 125604 200856 125656
rect 200908 125644 200914 125656
rect 249702 125644 249708 125656
rect 200908 125616 249708 125644
rect 200908 125604 200914 125616
rect 249702 125604 249708 125616
rect 249760 125604 249766 125656
rect 272702 125604 272708 125656
rect 272760 125644 272766 125656
rect 288342 125644 288348 125656
rect 272760 125616 288348 125644
rect 272760 125604 272766 125616
rect 288342 125604 288348 125616
rect 288400 125604 288406 125656
rect 266354 125536 266360 125588
rect 266412 125576 266418 125588
rect 275278 125576 275284 125588
rect 266412 125548 275284 125576
rect 266412 125536 266418 125548
rect 275278 125536 275284 125548
rect 275336 125536 275342 125588
rect 303706 125536 303712 125588
rect 303764 125576 303770 125588
rect 328454 125576 328460 125588
rect 303764 125548 328460 125576
rect 303764 125536 303770 125548
rect 328454 125536 328460 125548
rect 328512 125536 328518 125588
rect 202322 124924 202328 124976
rect 202380 124964 202386 124976
rect 228450 124964 228456 124976
rect 202380 124936 228456 124964
rect 202380 124924 202386 124936
rect 228450 124924 228456 124936
rect 228508 124924 228514 124976
rect 184382 124856 184388 124908
rect 184440 124896 184446 124908
rect 232682 124896 232688 124908
rect 184440 124868 232688 124896
rect 184440 124856 184446 124868
rect 232682 124856 232688 124868
rect 232740 124856 232746 124908
rect 266906 124856 266912 124908
rect 266964 124896 266970 124908
rect 285122 124896 285128 124908
rect 266964 124868 285128 124896
rect 266964 124856 266970 124868
rect 285122 124856 285128 124868
rect 285180 124856 285186 124908
rect 238110 124244 238116 124296
rect 238168 124284 238174 124296
rect 249610 124284 249616 124296
rect 238168 124256 249616 124284
rect 238168 124244 238174 124256
rect 249610 124244 249616 124256
rect 249668 124244 249674 124296
rect 232590 124176 232596 124228
rect 232648 124216 232654 124228
rect 249702 124216 249708 124228
rect 232648 124188 249708 124216
rect 232648 124176 232654 124188
rect 249702 124176 249708 124188
rect 249760 124176 249766 124228
rect 282822 124176 282828 124228
rect 282880 124216 282886 124228
rect 288342 124216 288348 124228
rect 282880 124188 288348 124216
rect 282880 124176 282886 124188
rect 288342 124176 288348 124188
rect 288400 124176 288406 124228
rect 303706 124108 303712 124160
rect 303764 124148 303770 124160
rect 327258 124148 327264 124160
rect 303764 124120 327264 124148
rect 303764 124108 303770 124120
rect 327258 124108 327264 124120
rect 327316 124108 327322 124160
rect 303798 124040 303804 124092
rect 303856 124080 303862 124092
rect 325694 124080 325700 124092
rect 303856 124052 325700 124080
rect 303856 124040 303862 124052
rect 325694 124040 325700 124052
rect 325752 124040 325758 124092
rect 164878 123428 164884 123480
rect 164936 123468 164942 123480
rect 231302 123468 231308 123480
rect 164936 123440 231308 123468
rect 164936 123428 164942 123440
rect 231302 123428 231308 123440
rect 231360 123428 231366 123480
rect 272794 123428 272800 123480
rect 272852 123468 272858 123480
rect 287882 123468 287888 123480
rect 272852 123440 287888 123468
rect 272852 123428 272858 123440
rect 287882 123428 287888 123440
rect 287940 123428 287946 123480
rect 266354 123156 266360 123208
rect 266412 123196 266418 123208
rect 268470 123196 268476 123208
rect 266412 123168 268476 123196
rect 266412 123156 266418 123168
rect 268470 123156 268476 123168
rect 268528 123156 268534 123208
rect 243722 122884 243728 122936
rect 243780 122924 243786 122936
rect 249518 122924 249524 122936
rect 243780 122896 249524 122924
rect 243780 122884 243786 122896
rect 249518 122884 249524 122896
rect 249576 122884 249582 122936
rect 185670 122816 185676 122868
rect 185728 122856 185734 122868
rect 248966 122856 248972 122868
rect 185728 122828 248972 122856
rect 185728 122816 185734 122828
rect 248966 122816 248972 122828
rect 249024 122816 249030 122868
rect 275278 122816 275284 122868
rect 275336 122856 275342 122868
rect 287974 122856 287980 122868
rect 275336 122828 287980 122856
rect 275336 122816 275342 122828
rect 287974 122816 287980 122828
rect 288032 122816 288038 122868
rect 266538 122748 266544 122800
rect 266596 122788 266602 122800
rect 286318 122788 286324 122800
rect 266596 122760 286324 122788
rect 266596 122748 266602 122760
rect 286318 122748 286324 122760
rect 286376 122748 286382 122800
rect 303614 122748 303620 122800
rect 303672 122788 303678 122800
rect 324406 122788 324412 122800
rect 303672 122760 324412 122788
rect 303672 122748 303678 122760
rect 324406 122748 324412 122760
rect 324464 122748 324470 122800
rect 266354 122680 266360 122732
rect 266412 122720 266418 122732
rect 282454 122720 282460 122732
rect 266412 122692 282460 122720
rect 266412 122680 266418 122692
rect 282454 122680 282460 122692
rect 282512 122680 282518 122732
rect 191190 122068 191196 122120
rect 191248 122108 191254 122120
rect 238018 122108 238024 122120
rect 191248 122080 238024 122108
rect 191248 122068 191254 122080
rect 238018 122068 238024 122080
rect 238076 122068 238082 122120
rect 239398 121524 239404 121576
rect 239456 121564 239462 121576
rect 248782 121564 248788 121576
rect 239456 121536 248788 121564
rect 239456 121524 239462 121536
rect 248782 121524 248788 121536
rect 248840 121524 248846 121576
rect 166258 121456 166264 121508
rect 166316 121496 166322 121508
rect 249702 121496 249708 121508
rect 166316 121468 249708 121496
rect 166316 121456 166322 121468
rect 249702 121456 249708 121468
rect 249760 121456 249766 121508
rect 283742 121456 283748 121508
rect 283800 121496 283806 121508
rect 288250 121496 288256 121508
rect 283800 121468 288256 121496
rect 283800 121456 283806 121468
rect 288250 121456 288256 121468
rect 288308 121456 288314 121508
rect 303798 121388 303804 121440
rect 303856 121428 303862 121440
rect 320358 121428 320364 121440
rect 303856 121400 320364 121428
rect 303856 121388 303862 121400
rect 320358 121388 320364 121400
rect 320416 121388 320422 121440
rect 222838 120708 222844 120760
rect 222896 120748 222902 120760
rect 236730 120748 236736 120760
rect 222896 120720 236736 120748
rect 222896 120708 222902 120720
rect 236730 120708 236736 120720
rect 236788 120708 236794 120760
rect 269758 120708 269764 120760
rect 269816 120748 269822 120760
rect 287146 120748 287152 120760
rect 269816 120720 287152 120748
rect 269816 120708 269822 120720
rect 287146 120708 287152 120720
rect 287204 120708 287210 120760
rect 238018 120164 238024 120216
rect 238076 120204 238082 120216
rect 249702 120204 249708 120216
rect 238076 120176 249708 120204
rect 238076 120164 238082 120176
rect 249702 120164 249708 120176
rect 249760 120164 249766 120216
rect 264238 120164 264244 120216
rect 264296 120204 264302 120216
rect 264296 120176 267734 120204
rect 264296 120164 264302 120176
rect 225598 120096 225604 120148
rect 225656 120136 225662 120148
rect 249610 120136 249616 120148
rect 225656 120108 249616 120136
rect 225656 120096 225662 120108
rect 249610 120096 249616 120108
rect 249668 120096 249674 120148
rect 264790 120096 264796 120148
rect 264848 120136 264854 120148
rect 266630 120136 266636 120148
rect 264848 120108 266636 120136
rect 264848 120096 264854 120108
rect 266630 120096 266636 120108
rect 266688 120096 266694 120148
rect 267706 120136 267734 120176
rect 288250 120136 288256 120148
rect 267706 120108 288256 120136
rect 288250 120096 288256 120108
rect 288308 120096 288314 120148
rect 266538 120028 266544 120080
rect 266596 120068 266602 120080
rect 286502 120068 286508 120080
rect 266596 120040 286508 120068
rect 266596 120028 266602 120040
rect 286502 120028 286508 120040
rect 286560 120028 286566 120080
rect 303798 120028 303804 120080
rect 303856 120068 303862 120080
rect 318886 120068 318892 120080
rect 303856 120040 318892 120068
rect 303856 120028 303862 120040
rect 318886 120028 318892 120040
rect 318944 120028 318950 120080
rect 266354 119960 266360 120012
rect 266412 120000 266418 120012
rect 281074 120000 281080 120012
rect 266412 119972 281080 120000
rect 266412 119960 266418 119972
rect 281074 119960 281080 119972
rect 281132 119960 281138 120012
rect 184290 118736 184296 118788
rect 184348 118776 184354 118788
rect 249702 118776 249708 118788
rect 184348 118748 249708 118776
rect 184348 118736 184354 118748
rect 249702 118736 249708 118748
rect 249760 118736 249766 118788
rect 182910 118668 182916 118720
rect 182968 118708 182974 118720
rect 248782 118708 248788 118720
rect 182968 118680 248788 118708
rect 182968 118668 182974 118680
rect 248782 118668 248788 118680
rect 248840 118668 248846 118720
rect 285122 118668 285128 118720
rect 285180 118708 285186 118720
rect 287606 118708 287612 118720
rect 285180 118680 287612 118708
rect 285180 118668 285186 118680
rect 287606 118668 287612 118680
rect 287664 118668 287670 118720
rect 266354 118600 266360 118652
rect 266412 118640 266418 118652
rect 279418 118640 279424 118652
rect 266412 118612 279424 118640
rect 266412 118600 266418 118612
rect 279418 118600 279424 118612
rect 279476 118600 279482 118652
rect 303890 118600 303896 118652
rect 303948 118640 303954 118652
rect 311986 118640 311992 118652
rect 303948 118612 311992 118640
rect 303948 118600 303954 118612
rect 311986 118600 311992 118612
rect 312044 118600 312050 118652
rect 266538 118532 266544 118584
rect 266596 118572 266602 118584
rect 274174 118572 274180 118584
rect 266596 118544 274180 118572
rect 266596 118532 266602 118544
rect 274174 118532 274180 118544
rect 274232 118532 274238 118584
rect 303798 118396 303804 118448
rect 303856 118436 303862 118448
rect 307846 118436 307852 118448
rect 303856 118408 307852 118436
rect 303856 118396 303862 118408
rect 307846 118396 307852 118408
rect 307904 118396 307910 118448
rect 186958 117920 186964 117972
rect 187016 117960 187022 117972
rect 249610 117960 249616 117972
rect 187016 117932 249616 117960
rect 187016 117920 187022 117932
rect 249610 117920 249616 117932
rect 249668 117920 249674 117972
rect 278498 117444 278504 117496
rect 278556 117484 278562 117496
rect 282822 117484 282828 117496
rect 278556 117456 282828 117484
rect 278556 117444 278562 117456
rect 282822 117444 282828 117456
rect 282880 117444 282886 117496
rect 235994 117308 236000 117360
rect 236052 117348 236058 117360
rect 248782 117348 248788 117360
rect 236052 117320 248788 117348
rect 236052 117308 236058 117320
rect 248782 117308 248788 117320
rect 248840 117308 248846 117360
rect 279510 117308 279516 117360
rect 279568 117348 279574 117360
rect 288250 117348 288256 117360
rect 279568 117320 288256 117348
rect 279568 117308 279574 117320
rect 288250 117308 288256 117320
rect 288308 117308 288314 117360
rect 266354 117240 266360 117292
rect 266412 117280 266418 117292
rect 272518 117280 272524 117292
rect 266412 117252 272524 117280
rect 266412 117240 266418 117252
rect 272518 117240 272524 117252
rect 272576 117240 272582 117292
rect 303798 117240 303804 117292
rect 303856 117280 303862 117292
rect 314654 117280 314660 117292
rect 303856 117252 314660 117280
rect 303856 117240 303862 117252
rect 314654 117240 314660 117252
rect 314712 117240 314718 117292
rect 266262 117172 266268 117224
rect 266320 117212 266326 117224
rect 266630 117212 266636 117224
rect 266320 117184 266636 117212
rect 266320 117172 266326 117184
rect 266630 117172 266636 117184
rect 266688 117172 266694 117224
rect 170674 116560 170680 116612
rect 170732 116600 170738 116612
rect 235994 116600 236000 116612
rect 170732 116572 236000 116600
rect 170732 116560 170738 116572
rect 235994 116560 236000 116572
rect 236052 116560 236058 116612
rect 269022 116560 269028 116612
rect 269080 116600 269086 116612
rect 285214 116600 285220 116612
rect 269080 116572 285220 116600
rect 269080 116560 269086 116572
rect 285214 116560 285220 116572
rect 285272 116560 285278 116612
rect 266354 116152 266360 116204
rect 266412 116192 266418 116204
rect 268562 116192 268568 116204
rect 266412 116164 268568 116192
rect 266412 116152 266418 116164
rect 268562 116152 268568 116164
rect 268620 116152 268626 116204
rect 285582 116016 285588 116068
rect 285640 116056 285646 116068
rect 287422 116056 287428 116068
rect 285640 116028 287428 116056
rect 285640 116016 285646 116028
rect 287422 116016 287428 116028
rect 287480 116016 287486 116068
rect 224310 115948 224316 116000
rect 224368 115988 224374 116000
rect 248782 115988 248788 116000
rect 224368 115960 248788 115988
rect 224368 115948 224374 115960
rect 248782 115948 248788 115960
rect 248840 115948 248846 116000
rect 272610 115948 272616 116000
rect 272668 115988 272674 116000
rect 288158 115988 288164 116000
rect 272668 115960 288164 115988
rect 272668 115948 272674 115960
rect 288158 115948 288164 115960
rect 288216 115948 288222 116000
rect 266538 115880 266544 115932
rect 266596 115920 266602 115932
rect 285030 115920 285036 115932
rect 266596 115892 285036 115920
rect 266596 115880 266602 115892
rect 285030 115880 285036 115892
rect 285088 115880 285094 115932
rect 303798 115880 303804 115932
rect 303856 115920 303862 115932
rect 310514 115920 310520 115932
rect 303856 115892 310520 115920
rect 303856 115880 303862 115892
rect 310514 115880 310520 115892
rect 310572 115880 310578 115932
rect 266354 115812 266360 115864
rect 266412 115852 266418 115864
rect 271138 115852 271144 115864
rect 266412 115824 271144 115852
rect 266412 115812 266418 115824
rect 271138 115812 271144 115824
rect 271196 115812 271202 115864
rect 303614 115404 303620 115456
rect 303672 115444 303678 115456
rect 306466 115444 306472 115456
rect 303672 115416 306472 115444
rect 303672 115404 303678 115416
rect 306466 115404 306472 115416
rect 306524 115404 306530 115456
rect 238202 114520 238208 114572
rect 238260 114560 238266 114572
rect 249702 114560 249708 114572
rect 238260 114532 249708 114560
rect 238260 114520 238266 114532
rect 249702 114520 249708 114532
rect 249760 114520 249766 114572
rect 285214 114520 285220 114572
rect 285272 114560 285278 114572
rect 288250 114560 288256 114572
rect 285272 114532 288256 114560
rect 285272 114520 285278 114532
rect 288250 114520 288256 114532
rect 288308 114520 288314 114572
rect 266538 114452 266544 114504
rect 266596 114492 266602 114504
rect 275554 114492 275560 114504
rect 266596 114464 275560 114492
rect 266596 114452 266602 114464
rect 275554 114452 275560 114464
rect 275612 114452 275618 114504
rect 303798 114452 303804 114504
rect 303856 114492 303862 114504
rect 316034 114492 316040 114504
rect 303856 114464 316040 114492
rect 303856 114452 303862 114464
rect 316034 114452 316040 114464
rect 316092 114452 316098 114504
rect 273162 113772 273168 113824
rect 273220 113812 273226 113824
rect 282454 113812 282460 113824
rect 273220 113784 282460 113812
rect 273220 113772 273226 113784
rect 282454 113772 282460 113784
rect 282512 113772 282518 113824
rect 266354 113636 266360 113688
rect 266412 113676 266418 113688
rect 269850 113676 269856 113688
rect 266412 113648 269856 113676
rect 266412 113636 266418 113648
rect 269850 113636 269856 113648
rect 269908 113636 269914 113688
rect 173434 113228 173440 113280
rect 173492 113268 173498 113280
rect 230474 113268 230480 113280
rect 173492 113240 230480 113268
rect 173492 113228 173498 113240
rect 230474 113228 230480 113240
rect 230532 113228 230538 113280
rect 235350 113228 235356 113280
rect 235408 113268 235414 113280
rect 249702 113268 249708 113280
rect 235408 113240 249708 113268
rect 235408 113228 235414 113240
rect 249702 113228 249708 113240
rect 249760 113228 249766 113280
rect 284018 113228 284024 113280
rect 284076 113268 284082 113280
rect 287974 113268 287980 113280
rect 284076 113240 287980 113268
rect 284076 113228 284082 113240
rect 287974 113228 287980 113240
rect 288032 113228 288038 113280
rect 167822 113160 167828 113212
rect 167880 113200 167886 113212
rect 249610 113200 249616 113212
rect 167880 113172 249616 113200
rect 167880 113160 167886 113172
rect 249610 113160 249616 113172
rect 249668 113160 249674 113212
rect 275370 113160 275376 113212
rect 275428 113200 275434 113212
rect 287606 113200 287612 113212
rect 275428 113172 287612 113200
rect 275428 113160 275434 113172
rect 287606 113160 287612 113172
rect 287664 113160 287670 113212
rect 230474 113092 230480 113144
rect 230532 113132 230538 113144
rect 243722 113132 243728 113144
rect 230532 113104 243728 113132
rect 230532 113092 230538 113104
rect 243722 113092 243728 113104
rect 243780 113092 243786 113144
rect 266538 113092 266544 113144
rect 266596 113132 266602 113144
rect 289078 113132 289084 113144
rect 266596 113104 289084 113132
rect 266596 113092 266602 113104
rect 289078 113092 289084 113104
rect 289136 113092 289142 113144
rect 303798 113092 303804 113144
rect 303856 113132 303862 113144
rect 307754 113132 307760 113144
rect 303856 113104 307760 113132
rect 303856 113092 303862 113104
rect 307754 113092 307760 113104
rect 307812 113092 307818 113144
rect 266354 113024 266360 113076
rect 266412 113064 266418 113076
rect 278222 113064 278228 113076
rect 266412 113036 278228 113064
rect 266412 113024 266418 113036
rect 278222 113024 278228 113036
rect 278280 113024 278286 113076
rect 303706 112752 303712 112804
rect 303764 112792 303770 112804
rect 306650 112792 306656 112804
rect 303764 112764 306656 112792
rect 303764 112752 303770 112764
rect 306650 112752 306656 112764
rect 306708 112752 306714 112804
rect 174630 112412 174636 112464
rect 174688 112452 174694 112464
rect 224218 112452 224224 112464
rect 174688 112424 224224 112452
rect 174688 112412 174694 112424
rect 224218 112412 224224 112424
rect 224276 112412 224282 112464
rect 243630 111868 243636 111920
rect 243688 111908 243694 111920
rect 248966 111908 248972 111920
rect 243688 111880 248972 111908
rect 243688 111868 243694 111880
rect 248966 111868 248972 111880
rect 249024 111868 249030 111920
rect 244918 111800 244924 111852
rect 244976 111840 244982 111852
rect 249242 111840 249248 111852
rect 244976 111812 249248 111840
rect 244976 111800 244982 111812
rect 249242 111800 249248 111812
rect 249300 111800 249306 111852
rect 278406 111800 278412 111852
rect 278464 111840 278470 111852
rect 285122 111840 285128 111852
rect 278464 111812 285128 111840
rect 278464 111800 278470 111812
rect 285122 111800 285128 111812
rect 285180 111800 285186 111852
rect 168282 111732 168288 111784
rect 168340 111772 168346 111784
rect 178862 111772 178868 111784
rect 168340 111744 178868 111772
rect 168340 111732 168346 111744
rect 178862 111732 178868 111744
rect 178920 111732 178926 111784
rect 303706 111732 303712 111784
rect 303764 111772 303770 111784
rect 325786 111772 325792 111784
rect 303764 111744 325792 111772
rect 303764 111732 303770 111744
rect 325786 111732 325792 111744
rect 325844 111732 325850 111784
rect 303798 111664 303804 111716
rect 303856 111704 303862 111716
rect 313274 111704 313280 111716
rect 303856 111676 313280 111704
rect 303856 111664 303862 111676
rect 313274 111664 313280 111676
rect 313332 111664 313338 111716
rect 266998 111120 267004 111172
rect 267056 111160 267062 111172
rect 272610 111160 272616 111172
rect 267056 111132 272616 111160
rect 267056 111120 267062 111132
rect 272610 111120 272616 111132
rect 272668 111120 272674 111172
rect 268470 111052 268476 111104
rect 268528 111092 268534 111104
rect 278498 111092 278504 111104
rect 268528 111064 278504 111092
rect 268528 111052 268534 111064
rect 278498 111052 278504 111064
rect 278556 111052 278562 111104
rect 180334 110508 180340 110560
rect 180392 110548 180398 110560
rect 248966 110548 248972 110560
rect 180392 110520 248972 110548
rect 180392 110508 180398 110520
rect 248966 110508 248972 110520
rect 249024 110508 249030 110560
rect 282914 110508 282920 110560
rect 282972 110548 282978 110560
rect 287974 110548 287980 110560
rect 282972 110520 287980 110548
rect 282972 110508 282978 110520
rect 287974 110508 287980 110520
rect 288032 110508 288038 110560
rect 172054 110440 172060 110492
rect 172112 110480 172118 110492
rect 249242 110480 249248 110492
rect 172112 110452 249248 110480
rect 172112 110440 172118 110452
rect 249242 110440 249248 110452
rect 249300 110440 249306 110492
rect 278038 110440 278044 110492
rect 278096 110480 278102 110492
rect 288250 110480 288256 110492
rect 278096 110452 288256 110480
rect 278096 110440 278102 110452
rect 288250 110440 288256 110452
rect 288308 110440 288314 110492
rect 167914 110372 167920 110424
rect 167972 110412 167978 110424
rect 180150 110412 180156 110424
rect 167972 110384 180156 110412
rect 167972 110372 167978 110384
rect 180150 110372 180156 110384
rect 180208 110372 180214 110424
rect 266446 110372 266452 110424
rect 266504 110412 266510 110424
rect 278130 110412 278136 110424
rect 266504 110384 278136 110412
rect 266504 110372 266510 110384
rect 278130 110372 278136 110384
rect 278188 110372 278194 110424
rect 266354 110304 266360 110356
rect 266412 110344 266418 110356
rect 275462 110344 275468 110356
rect 266412 110316 275468 110344
rect 266412 110304 266418 110316
rect 275462 110304 275468 110316
rect 275520 110304 275526 110356
rect 211798 109080 211804 109132
rect 211856 109120 211862 109132
rect 249702 109120 249708 109132
rect 211856 109092 249708 109120
rect 211856 109080 211862 109092
rect 249702 109080 249708 109092
rect 249760 109080 249766 109132
rect 283558 109080 283564 109132
rect 283616 109120 283622 109132
rect 288250 109120 288256 109132
rect 283616 109092 288256 109120
rect 283616 109080 283622 109092
rect 288250 109080 288256 109092
rect 288308 109080 288314 109132
rect 180242 109012 180248 109064
rect 180300 109052 180306 109064
rect 249610 109052 249616 109064
rect 180300 109024 249616 109052
rect 180300 109012 180306 109024
rect 249610 109012 249616 109024
rect 249668 109012 249674 109064
rect 278222 109012 278228 109064
rect 278280 109052 278286 109064
rect 288342 109052 288348 109064
rect 278280 109024 288348 109052
rect 278280 109012 278286 109024
rect 288342 109012 288348 109024
rect 288400 109012 288406 109064
rect 266354 108944 266360 108996
rect 266412 108984 266418 108996
rect 280982 108984 280988 108996
rect 266412 108956 280988 108984
rect 266412 108944 266418 108956
rect 280982 108944 280988 108956
rect 281040 108944 281046 108996
rect 303798 108944 303804 108996
rect 303856 108984 303862 108996
rect 321554 108984 321560 108996
rect 303856 108956 321560 108984
rect 303856 108944 303862 108956
rect 321554 108944 321560 108956
rect 321612 108944 321618 108996
rect 170398 108264 170404 108316
rect 170456 108304 170462 108316
rect 229830 108304 229836 108316
rect 170456 108276 229836 108304
rect 170456 108264 170462 108276
rect 229830 108264 229836 108276
rect 229888 108264 229894 108316
rect 234154 107720 234160 107772
rect 234212 107760 234218 107772
rect 249702 107760 249708 107772
rect 234212 107732 249708 107760
rect 234212 107720 234218 107732
rect 249702 107720 249708 107732
rect 249760 107720 249766 107772
rect 231302 107652 231308 107704
rect 231360 107692 231366 107704
rect 249518 107692 249524 107704
rect 231360 107664 249524 107692
rect 231360 107652 231366 107664
rect 249518 107652 249524 107664
rect 249576 107652 249582 107704
rect 267182 107652 267188 107704
rect 267240 107692 267246 107704
rect 288342 107692 288348 107704
rect 267240 107664 288348 107692
rect 267240 107652 267246 107664
rect 288342 107652 288348 107664
rect 288400 107652 288406 107704
rect 266354 107584 266360 107636
rect 266412 107624 266418 107636
rect 279694 107624 279700 107636
rect 266412 107596 279700 107624
rect 266412 107584 266418 107596
rect 279694 107584 279700 107596
rect 279752 107584 279758 107636
rect 303798 107584 303804 107636
rect 303856 107624 303862 107636
rect 309134 107624 309140 107636
rect 303856 107596 309140 107624
rect 303856 107584 303862 107596
rect 309134 107584 309140 107596
rect 309192 107584 309198 107636
rect 266446 107516 266452 107568
rect 266504 107556 266510 107568
rect 276934 107556 276940 107568
rect 266504 107528 276940 107556
rect 266504 107516 266510 107528
rect 276934 107516 276940 107528
rect 276992 107516 276998 107568
rect 285122 106428 285128 106480
rect 285180 106468 285186 106480
rect 287974 106468 287980 106480
rect 285180 106440 287980 106468
rect 285180 106428 285186 106440
rect 287974 106428 287980 106440
rect 288032 106428 288038 106480
rect 191282 106360 191288 106412
rect 191340 106400 191346 106412
rect 249702 106400 249708 106412
rect 191340 106372 249708 106400
rect 191340 106360 191346 106372
rect 249702 106360 249708 106372
rect 249760 106360 249766 106412
rect 280982 106360 280988 106412
rect 281040 106400 281046 106412
rect 288342 106400 288348 106412
rect 281040 106372 288348 106400
rect 281040 106360 281046 106372
rect 288342 106360 288348 106372
rect 288400 106360 288406 106412
rect 166350 106292 166356 106344
rect 166408 106332 166414 106344
rect 249518 106332 249524 106344
rect 166408 106304 249524 106332
rect 166408 106292 166414 106304
rect 249518 106292 249524 106304
rect 249576 106292 249582 106344
rect 266354 106224 266360 106276
rect 266412 106264 266418 106276
rect 282270 106264 282276 106276
rect 266412 106236 282276 106264
rect 266412 106224 266418 106236
rect 282270 106224 282276 106236
rect 282328 106224 282334 106276
rect 200758 104932 200764 104984
rect 200816 104972 200822 104984
rect 249702 104972 249708 104984
rect 200816 104944 249708 104972
rect 200816 104932 200822 104944
rect 249702 104932 249708 104944
rect 249760 104932 249766 104984
rect 281074 104932 281080 104984
rect 281132 104972 281138 104984
rect 287974 104972 287980 104984
rect 281132 104944 287980 104972
rect 281132 104932 281138 104944
rect 287974 104932 287980 104944
rect 288032 104932 288038 104984
rect 167730 104864 167736 104916
rect 167788 104904 167794 104916
rect 248782 104904 248788 104916
rect 167788 104876 248788 104904
rect 167788 104864 167794 104876
rect 248782 104864 248788 104876
rect 248840 104864 248846 104916
rect 283834 104864 283840 104916
rect 283892 104904 283898 104916
rect 288342 104904 288348 104916
rect 283892 104876 288348 104904
rect 283892 104864 283898 104876
rect 288342 104864 288348 104876
rect 288400 104864 288406 104916
rect 303798 104796 303804 104848
rect 303856 104836 303862 104848
rect 314746 104836 314752 104848
rect 303856 104808 314752 104836
rect 303856 104796 303862 104808
rect 314746 104796 314752 104808
rect 314804 104796 314810 104848
rect 272886 104184 272892 104236
rect 272944 104224 272950 104236
rect 282914 104224 282920 104236
rect 272944 104196 282920 104224
rect 272944 104184 272950 104196
rect 282914 104184 282920 104196
rect 282972 104184 282978 104236
rect 169110 104116 169116 104168
rect 169168 104156 169174 104168
rect 211890 104156 211896 104168
rect 169168 104128 211896 104156
rect 169168 104116 169174 104128
rect 211890 104116 211896 104128
rect 211948 104116 211954 104168
rect 264422 104116 264428 104168
rect 264480 104156 264486 104168
rect 283742 104156 283748 104168
rect 264480 104128 283748 104156
rect 264480 104116 264486 104128
rect 283742 104116 283748 104128
rect 283800 104116 283806 104168
rect 266354 104048 266360 104100
rect 266412 104088 266418 104100
rect 269942 104088 269948 104100
rect 266412 104060 269948 104088
rect 266412 104048 266418 104060
rect 269942 104048 269948 104060
rect 270000 104048 270006 104100
rect 171962 103504 171968 103556
rect 172020 103544 172026 103556
rect 249702 103544 249708 103556
rect 172020 103516 249708 103544
rect 172020 103504 172026 103516
rect 249702 103504 249708 103516
rect 249760 103504 249766 103556
rect 266446 103436 266452 103488
rect 266504 103476 266510 103488
rect 284938 103476 284944 103488
rect 266504 103448 284944 103476
rect 266504 103436 266510 103448
rect 284938 103436 284944 103448
rect 284996 103436 285002 103488
rect 266354 103368 266360 103420
rect 266412 103408 266418 103420
rect 271230 103408 271236 103420
rect 266412 103380 271236 103408
rect 266412 103368 266418 103380
rect 271230 103368 271236 103380
rect 271288 103368 271294 103420
rect 281534 102280 281540 102332
rect 281592 102320 281598 102332
rect 285214 102320 285220 102332
rect 281592 102292 285220 102320
rect 281592 102280 281598 102292
rect 285214 102280 285220 102292
rect 285272 102280 285278 102332
rect 278130 102212 278136 102264
rect 278188 102252 278194 102264
rect 282454 102252 282460 102264
rect 278188 102224 282460 102252
rect 278188 102212 278194 102224
rect 282454 102212 282460 102224
rect 282512 102212 282518 102264
rect 285030 102212 285036 102264
rect 285088 102252 285094 102264
rect 288342 102252 288348 102264
rect 285088 102224 288348 102252
rect 285088 102212 285094 102224
rect 288342 102212 288348 102224
rect 288400 102212 288406 102264
rect 174722 102144 174728 102196
rect 174780 102184 174786 102196
rect 249702 102184 249708 102196
rect 174780 102156 249708 102184
rect 174780 102144 174786 102156
rect 249702 102144 249708 102156
rect 249760 102144 249766 102196
rect 271506 102144 271512 102196
rect 271564 102184 271570 102196
rect 278406 102184 278412 102196
rect 271564 102156 278412 102184
rect 271564 102144 271570 102156
rect 278406 102144 278412 102156
rect 278464 102144 278470 102196
rect 284294 102144 284300 102196
rect 284352 102184 284358 102196
rect 288250 102184 288256 102196
rect 284352 102156 288256 102184
rect 284352 102144 284358 102156
rect 288250 102144 288256 102156
rect 288308 102144 288314 102196
rect 303706 102076 303712 102128
rect 303764 102116 303770 102128
rect 323026 102116 323032 102128
rect 303764 102088 323032 102116
rect 303764 102076 303770 102088
rect 323026 102076 323032 102088
rect 323084 102076 323090 102128
rect 266354 102008 266360 102060
rect 266412 102048 266418 102060
rect 270034 102048 270040 102060
rect 266412 102020 270040 102048
rect 266412 102008 266418 102020
rect 270034 102008 270040 102020
rect 270092 102008 270098 102060
rect 166442 101396 166448 101448
rect 166500 101436 166506 101448
rect 200850 101436 200856 101448
rect 166500 101408 200856 101436
rect 166500 101396 166506 101408
rect 200850 101396 200856 101408
rect 200908 101396 200914 101448
rect 218790 101396 218796 101448
rect 218848 101436 218854 101448
rect 251818 101436 251824 101448
rect 218848 101408 251824 101436
rect 218848 101396 218854 101408
rect 251818 101396 251824 101408
rect 251876 101396 251882 101448
rect 284938 100784 284944 100836
rect 284996 100824 285002 100836
rect 287606 100824 287612 100836
rect 284996 100796 287612 100824
rect 284996 100784 285002 100796
rect 287606 100784 287612 100796
rect 287664 100784 287670 100836
rect 177482 100716 177488 100768
rect 177540 100756 177546 100768
rect 249150 100756 249156 100768
rect 177540 100728 249156 100756
rect 177540 100716 177546 100728
rect 249150 100716 249156 100728
rect 249208 100716 249214 100768
rect 265618 100716 265624 100768
rect 265676 100756 265682 100768
rect 272058 100756 272064 100768
rect 265676 100728 272064 100756
rect 265676 100716 265682 100728
rect 272058 100716 272064 100728
rect 272116 100716 272122 100768
rect 279694 100716 279700 100768
rect 279752 100756 279758 100768
rect 288342 100756 288348 100768
rect 279752 100728 288348 100756
rect 279752 100716 279758 100728
rect 288342 100716 288348 100728
rect 288400 100716 288406 100768
rect 266354 100648 266360 100700
rect 266412 100688 266418 100700
rect 282362 100688 282368 100700
rect 266412 100660 282368 100688
rect 266412 100648 266418 100660
rect 282362 100648 282368 100660
rect 282420 100648 282426 100700
rect 266446 100580 266452 100632
rect 266504 100620 266510 100632
rect 272794 100620 272800 100632
rect 266504 100592 272800 100620
rect 266504 100580 266510 100592
rect 272794 100580 272800 100592
rect 272852 100580 272858 100632
rect 164970 99968 164976 100020
rect 165028 100008 165034 100020
rect 249058 100008 249064 100020
rect 165028 99980 249064 100008
rect 165028 99968 165034 99980
rect 249058 99968 249064 99980
rect 249116 99968 249122 100020
rect 284110 99424 284116 99476
rect 284168 99464 284174 99476
rect 288250 99464 288256 99476
rect 284168 99436 288256 99464
rect 284168 99424 284174 99436
rect 288250 99424 288256 99436
rect 288308 99424 288314 99476
rect 214650 99356 214656 99408
rect 214708 99396 214714 99408
rect 249702 99396 249708 99408
rect 214708 99368 249708 99396
rect 214708 99356 214714 99368
rect 249702 99356 249708 99368
rect 249760 99356 249766 99408
rect 272610 99356 272616 99408
rect 272668 99396 272674 99408
rect 288342 99396 288348 99408
rect 272668 99368 288348 99396
rect 272668 99356 272674 99368
rect 288342 99356 288348 99368
rect 288400 99356 288406 99408
rect 266446 99288 266452 99340
rect 266504 99328 266510 99340
rect 274266 99328 274272 99340
rect 266504 99300 274272 99328
rect 266504 99288 266510 99300
rect 274266 99288 274272 99300
rect 274324 99288 274330 99340
rect 276934 98676 276940 98728
rect 276992 98716 276998 98728
rect 282914 98716 282920 98728
rect 276992 98688 282920 98716
rect 276992 98676 276998 98688
rect 282914 98676 282920 98688
rect 282972 98676 282978 98728
rect 273898 98608 273904 98660
rect 273956 98648 273962 98660
rect 281534 98648 281540 98660
rect 273956 98620 281540 98648
rect 273956 98608 273962 98620
rect 281534 98608 281540 98620
rect 281592 98608 281598 98660
rect 283650 98132 283656 98184
rect 283708 98172 283714 98184
rect 287882 98172 287888 98184
rect 283708 98144 287888 98172
rect 283708 98132 283714 98144
rect 287882 98132 287888 98144
rect 287940 98132 287946 98184
rect 203518 98064 203524 98116
rect 203576 98104 203582 98116
rect 249702 98104 249708 98116
rect 203576 98076 249708 98104
rect 203576 98064 203582 98076
rect 249702 98064 249708 98076
rect 249760 98064 249766 98116
rect 282362 98064 282368 98116
rect 282420 98104 282426 98116
rect 286778 98104 286784 98116
rect 282420 98076 286784 98104
rect 282420 98064 282426 98076
rect 286778 98064 286784 98076
rect 286836 98064 286842 98116
rect 171870 97996 171876 98048
rect 171928 98036 171934 98048
rect 249610 98036 249616 98048
rect 171928 98008 249616 98036
rect 171928 97996 171934 98008
rect 249610 97996 249616 98008
rect 249668 97996 249674 98048
rect 264054 97996 264060 98048
rect 264112 98036 264118 98048
rect 268286 98036 268292 98048
rect 264112 98008 268292 98036
rect 264112 97996 264118 98008
rect 268286 97996 268292 98008
rect 268344 97996 268350 98048
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 21358 97968 21364 97980
rect 3476 97940 21364 97968
rect 3476 97928 3482 97940
rect 21358 97928 21364 97940
rect 21416 97928 21422 97980
rect 210418 97928 210424 97980
rect 210476 97968 210482 97980
rect 252186 97968 252192 97980
rect 210476 97940 252192 97968
rect 210476 97928 210482 97940
rect 252186 97928 252192 97940
rect 252244 97928 252250 97980
rect 265802 97724 265808 97776
rect 265860 97764 265866 97776
rect 267274 97764 267280 97776
rect 265860 97736 267280 97764
rect 265860 97724 265866 97736
rect 267274 97724 267280 97736
rect 267332 97724 267338 97776
rect 178862 97248 178868 97300
rect 178920 97288 178926 97300
rect 209222 97288 209228 97300
rect 178920 97260 209228 97288
rect 178920 97248 178926 97260
rect 209222 97248 209228 97260
rect 209280 97248 209286 97300
rect 288342 97288 288348 97300
rect 267706 97260 288348 97288
rect 264054 96812 264060 96824
rect 259564 96784 264060 96812
rect 165522 96636 165528 96688
rect 165580 96676 165586 96688
rect 249702 96676 249708 96688
rect 165580 96648 249708 96676
rect 165580 96636 165586 96648
rect 249702 96636 249708 96648
rect 249760 96636 249766 96688
rect 252186 96636 252192 96688
rect 252244 96676 252250 96688
rect 259564 96676 259592 96784
rect 264054 96772 264060 96784
rect 264112 96772 264118 96824
rect 267706 96744 267734 97260
rect 288342 97248 288348 97260
rect 288400 97248 288406 97300
rect 252244 96648 257844 96676
rect 252244 96636 252250 96648
rect 257816 96076 257844 96648
rect 259472 96648 259592 96676
rect 261036 96716 267734 96744
rect 257798 96024 257804 96076
rect 257856 96024 257862 96076
rect 257890 96024 257896 96076
rect 257948 96064 257954 96076
rect 259472 96064 259500 96648
rect 261036 96076 261064 96716
rect 303890 96568 303896 96620
rect 303948 96608 303954 96620
rect 334066 96608 334072 96620
rect 303948 96580 334072 96608
rect 303948 96568 303954 96580
rect 334066 96568 334072 96580
rect 334124 96568 334130 96620
rect 257948 96036 259500 96064
rect 257948 96024 257954 96036
rect 261018 96024 261024 96076
rect 261076 96024 261082 96076
rect 165614 95956 165620 96008
rect 165672 95996 165678 96008
rect 214558 95996 214564 96008
rect 165672 95968 214564 95996
rect 165672 95956 165678 95968
rect 214558 95956 214564 95968
rect 214616 95956 214622 96008
rect 224862 95956 224868 96008
rect 224920 95996 224926 96008
rect 290918 95996 290924 96008
rect 224920 95968 290924 95996
rect 224920 95956 224926 95968
rect 290918 95956 290924 95968
rect 290976 95956 290982 96008
rect 168650 95888 168656 95940
rect 168708 95928 168714 95940
rect 247862 95928 247868 95940
rect 168708 95900 247868 95928
rect 168708 95888 168714 95900
rect 247862 95888 247868 95900
rect 247920 95888 247926 95940
rect 258718 95888 258724 95940
rect 258776 95928 258782 95940
rect 266262 95928 266268 95940
rect 258776 95900 266268 95928
rect 258776 95888 258782 95900
rect 266262 95888 266268 95900
rect 266320 95888 266326 95940
rect 271138 95208 271144 95260
rect 271196 95248 271202 95260
rect 278314 95248 278320 95260
rect 271196 95220 278320 95248
rect 271196 95208 271202 95220
rect 278314 95208 278320 95220
rect 278372 95208 278378 95260
rect 246390 95140 246396 95192
rect 246448 95180 246454 95192
rect 301498 95180 301504 95192
rect 246448 95152 301504 95180
rect 246448 95140 246454 95152
rect 301498 95140 301504 95152
rect 301556 95140 301562 95192
rect 289722 95072 289728 95124
rect 289780 95112 289786 95124
rect 291286 95112 291292 95124
rect 289780 95084 291292 95112
rect 289780 95072 289786 95084
rect 291286 95072 291292 95084
rect 291344 95072 291350 95124
rect 67726 94460 67732 94512
rect 67784 94500 67790 94512
rect 100018 94500 100024 94512
rect 67784 94472 100024 94500
rect 67784 94460 67790 94472
rect 100018 94460 100024 94472
rect 100076 94460 100082 94512
rect 181530 94460 181536 94512
rect 181588 94500 181594 94512
rect 248782 94500 248788 94512
rect 181588 94472 248788 94500
rect 181588 94460 181594 94472
rect 248782 94460 248788 94472
rect 248840 94460 248846 94512
rect 257338 94460 257344 94512
rect 257396 94500 257402 94512
rect 264146 94500 264152 94512
rect 257396 94472 264152 94500
rect 257396 94460 257402 94472
rect 264146 94460 264152 94472
rect 264204 94460 264210 94512
rect 162854 94392 162860 94444
rect 162912 94432 162918 94444
rect 165614 94432 165620 94444
rect 162912 94404 165620 94432
rect 162912 94392 162918 94404
rect 165614 94392 165620 94404
rect 165672 94392 165678 94444
rect 124030 93848 124036 93900
rect 124088 93888 124094 93900
rect 238110 93888 238116 93900
rect 124088 93860 238116 93888
rect 124088 93848 124094 93860
rect 238110 93848 238116 93860
rect 238168 93848 238174 93900
rect 267734 93780 267740 93832
rect 267792 93820 267798 93832
rect 295978 93820 295984 93832
rect 267792 93792 295984 93820
rect 267792 93780 267798 93792
rect 295978 93780 295984 93792
rect 296036 93780 296042 93832
rect 290918 93712 290924 93764
rect 290976 93752 290982 93764
rect 303798 93752 303804 93764
rect 290976 93724 303804 93752
rect 290976 93712 290982 93724
rect 303798 93712 303804 93724
rect 303856 93712 303862 93764
rect 67358 93168 67364 93220
rect 67416 93208 67422 93220
rect 88978 93208 88984 93220
rect 67416 93180 88984 93208
rect 67416 93168 67422 93180
rect 88978 93168 88984 93180
rect 89036 93168 89042 93220
rect 119706 93168 119712 93220
rect 119764 93208 119770 93220
rect 166258 93208 166264 93220
rect 119764 93180 166264 93208
rect 119764 93168 119770 93180
rect 166258 93168 166264 93180
rect 166316 93168 166322 93220
rect 170582 93168 170588 93220
rect 170640 93208 170646 93220
rect 177574 93208 177580 93220
rect 170640 93180 177580 93208
rect 170640 93168 170646 93180
rect 177574 93168 177580 93180
rect 177632 93168 177638 93220
rect 184382 93168 184388 93220
rect 184440 93208 184446 93220
rect 206370 93208 206376 93220
rect 184440 93180 206376 93208
rect 184440 93168 184446 93180
rect 206370 93168 206376 93180
rect 206428 93168 206434 93220
rect 246298 93168 246304 93220
rect 246356 93208 246362 93220
rect 265894 93208 265900 93220
rect 246356 93180 265900 93208
rect 246356 93168 246362 93180
rect 265894 93168 265900 93180
rect 265952 93168 265958 93220
rect 66070 93100 66076 93152
rect 66128 93140 66134 93152
rect 106182 93140 106188 93152
rect 66128 93112 106188 93140
rect 66128 93100 66134 93112
rect 106182 93100 106188 93112
rect 106240 93100 106246 93152
rect 121730 93100 121736 93152
rect 121788 93140 121794 93152
rect 185670 93140 185676 93152
rect 121788 93112 185676 93140
rect 121788 93100 121794 93112
rect 185670 93100 185676 93112
rect 185728 93100 185734 93152
rect 260098 93100 260104 93152
rect 260156 93140 260162 93152
rect 283834 93140 283840 93152
rect 260156 93112 283840 93140
rect 260156 93100 260162 93112
rect 283834 93100 283840 93112
rect 283892 93100 283898 93152
rect 136082 92420 136088 92472
rect 136140 92460 136146 92472
rect 173342 92460 173348 92472
rect 136140 92432 173348 92460
rect 136140 92420 136146 92432
rect 173342 92420 173348 92432
rect 173400 92420 173406 92472
rect 250714 92420 250720 92472
rect 250772 92460 250778 92472
rect 303614 92460 303620 92472
rect 250772 92432 303620 92460
rect 250772 92420 250778 92432
rect 303614 92420 303620 92432
rect 303672 92420 303678 92472
rect 151354 92352 151360 92404
rect 151412 92392 151418 92404
rect 162854 92392 162860 92404
rect 151412 92364 162860 92392
rect 151412 92352 151418 92364
rect 162854 92352 162860 92364
rect 162912 92352 162918 92404
rect 117222 91740 117228 91792
rect 117280 91780 117286 91792
rect 126882 91780 126888 91792
rect 117280 91752 126888 91780
rect 117280 91740 117286 91752
rect 126882 91740 126888 91752
rect 126940 91740 126946 91792
rect 164142 91740 164148 91792
rect 164200 91780 164206 91792
rect 235258 91780 235264 91792
rect 164200 91752 235264 91780
rect 164200 91740 164206 91752
rect 235258 91740 235264 91752
rect 235316 91740 235322 91792
rect 235902 91740 235908 91792
rect 235960 91780 235966 91792
rect 266446 91780 266452 91792
rect 235960 91752 266452 91780
rect 235960 91740 235966 91752
rect 266446 91740 266452 91752
rect 266504 91740 266510 91792
rect 267090 91740 267096 91792
rect 267148 91780 267154 91792
rect 274634 91780 274640 91792
rect 267148 91752 274640 91780
rect 267148 91740 267154 91752
rect 274634 91740 274640 91752
rect 274692 91740 274698 91792
rect 86862 91128 86868 91180
rect 86920 91168 86926 91180
rect 106918 91168 106924 91180
rect 86920 91140 106924 91168
rect 86920 91128 86926 91140
rect 106918 91128 106924 91140
rect 106976 91128 106982 91180
rect 114462 91128 114468 91180
rect 114520 91168 114526 91180
rect 134702 91168 134708 91180
rect 114520 91140 134708 91168
rect 114520 91128 114526 91140
rect 134702 91128 134708 91140
rect 134760 91128 134766 91180
rect 89070 91060 89076 91112
rect 89128 91100 89134 91112
rect 116578 91100 116584 91112
rect 89128 91072 116584 91100
rect 89128 91060 89134 91072
rect 116578 91060 116584 91072
rect 116636 91060 116642 91112
rect 127986 91060 127992 91112
rect 128044 91100 128050 91112
rect 128998 91100 129004 91112
rect 128044 91072 129004 91100
rect 128044 91060 128050 91072
rect 128998 91060 129004 91072
rect 129056 91060 129062 91112
rect 109954 90992 109960 91044
rect 110012 91032 110018 91044
rect 224310 91032 224316 91044
rect 110012 91004 224316 91032
rect 110012 90992 110018 91004
rect 224310 90992 224316 91004
rect 224368 90992 224374 91044
rect 236730 90992 236736 91044
rect 236788 91032 236794 91044
rect 303706 91032 303712 91044
rect 236788 91004 303712 91032
rect 236788 90992 236794 91004
rect 303706 90992 303712 91004
rect 303764 90992 303770 91044
rect 111610 90924 111616 90976
rect 111668 90964 111674 90976
rect 170674 90964 170680 90976
rect 111668 90936 170680 90964
rect 111668 90924 111674 90936
rect 170674 90924 170680 90936
rect 170732 90924 170738 90976
rect 65978 90312 65984 90364
rect 66036 90352 66042 90364
rect 111058 90352 111064 90364
rect 66036 90324 111064 90352
rect 66036 90312 66042 90324
rect 111058 90312 111064 90324
rect 111116 90312 111122 90364
rect 175918 90312 175924 90364
rect 175976 90352 175982 90364
rect 196710 90352 196716 90364
rect 175976 90324 196716 90352
rect 175976 90312 175982 90324
rect 196710 90312 196716 90324
rect 196768 90312 196774 90364
rect 198090 90312 198096 90364
rect 198148 90352 198154 90364
rect 286502 90352 286508 90364
rect 198148 90324 286508 90352
rect 198148 90312 198154 90324
rect 286502 90312 286508 90324
rect 286560 90312 286566 90364
rect 122834 89632 122840 89684
rect 122892 89672 122898 89684
rect 232590 89672 232596 89684
rect 122892 89644 232596 89672
rect 122892 89632 122898 89644
rect 232590 89632 232596 89644
rect 232648 89632 232654 89684
rect 251818 89632 251824 89684
rect 251876 89672 251882 89684
rect 301130 89672 301136 89684
rect 251876 89644 301136 89672
rect 251876 89632 251882 89644
rect 301130 89632 301136 89644
rect 301188 89632 301194 89684
rect 107470 89564 107476 89616
rect 107528 89604 107534 89616
rect 158714 89604 158720 89616
rect 107528 89576 158720 89604
rect 107528 89564 107534 89576
rect 158714 89564 158720 89576
rect 158772 89564 158778 89616
rect 98730 88952 98736 89004
rect 98788 88992 98794 89004
rect 122190 88992 122196 89004
rect 98788 88964 122196 88992
rect 98788 88952 98794 88964
rect 122190 88952 122196 88964
rect 122248 88952 122254 89004
rect 160094 88952 160100 89004
rect 160152 88992 160158 89004
rect 176010 88992 176016 89004
rect 160152 88964 176016 88992
rect 160152 88952 160158 88964
rect 176010 88952 176016 88964
rect 176068 88952 176074 89004
rect 196710 88952 196716 89004
rect 196768 88992 196774 89004
rect 264422 88992 264428 89004
rect 196768 88964 264428 88992
rect 196768 88952 196774 88964
rect 264422 88952 264428 88964
rect 264480 88952 264486 89004
rect 102594 88272 102600 88324
rect 102652 88312 102658 88324
rect 235350 88312 235356 88324
rect 102652 88284 235356 88312
rect 102652 88272 102658 88284
rect 235350 88272 235356 88284
rect 235408 88272 235414 88324
rect 134702 88204 134708 88256
rect 134760 88244 134766 88256
rect 164142 88244 164148 88256
rect 134760 88216 164148 88244
rect 134760 88204 134766 88216
rect 164142 88204 164148 88216
rect 164200 88204 164206 88256
rect 164970 87592 164976 87644
rect 165028 87632 165034 87644
rect 243630 87632 243636 87644
rect 165028 87604 243636 87632
rect 165028 87592 165034 87604
rect 243630 87592 243636 87604
rect 243688 87592 243694 87644
rect 260190 87592 260196 87644
rect 260248 87632 260254 87644
rect 272886 87632 272892 87644
rect 260248 87604 272892 87632
rect 260248 87592 260254 87604
rect 272886 87592 272892 87604
rect 272944 87592 272950 87644
rect 75914 86912 75920 86964
rect 75972 86952 75978 86964
rect 249334 86952 249340 86964
rect 75972 86924 249340 86952
rect 75972 86912 75978 86924
rect 249334 86912 249340 86924
rect 249392 86912 249398 86964
rect 113450 86844 113456 86896
rect 113508 86884 113514 86896
rect 182910 86884 182916 86896
rect 113508 86856 182916 86884
rect 113508 86844 113514 86856
rect 182910 86844 182916 86856
rect 182968 86844 182974 86896
rect 253198 86300 253204 86352
rect 253256 86340 253262 86352
rect 270126 86340 270132 86352
rect 253256 86312 270132 86340
rect 253256 86300 253262 86312
rect 270126 86300 270132 86312
rect 270184 86300 270190 86352
rect 66162 86232 66168 86284
rect 66220 86272 66226 86284
rect 107010 86272 107016 86284
rect 66220 86244 107016 86272
rect 66220 86232 66226 86244
rect 107010 86232 107016 86244
rect 107068 86232 107074 86284
rect 191098 86232 191104 86284
rect 191156 86272 191162 86284
rect 278130 86272 278136 86284
rect 191156 86244 278136 86272
rect 191156 86232 191162 86244
rect 278130 86232 278136 86244
rect 278188 86232 278194 86284
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 29638 85524 29644 85536
rect 3200 85496 29644 85524
rect 3200 85484 3206 85496
rect 29638 85484 29644 85496
rect 29696 85484 29702 85536
rect 125410 85484 125416 85536
rect 125468 85524 125474 85536
rect 166442 85524 166448 85536
rect 125468 85496 166448 85524
rect 125468 85484 125474 85496
rect 166442 85484 166448 85496
rect 166500 85484 166506 85536
rect 151630 85416 151636 85468
rect 151688 85456 151694 85468
rect 160094 85456 160100 85468
rect 151688 85428 160100 85456
rect 151688 85416 151694 85428
rect 160094 85416 160100 85428
rect 160152 85416 160158 85468
rect 206278 84872 206284 84924
rect 206336 84912 206342 84924
rect 275554 84912 275560 84924
rect 206336 84884 275560 84912
rect 206336 84872 206342 84884
rect 275554 84872 275560 84884
rect 275612 84872 275618 84924
rect 160738 84804 160744 84856
rect 160796 84844 160802 84856
rect 263042 84844 263048 84856
rect 160796 84816 263048 84844
rect 160796 84804 160802 84816
rect 263042 84804 263048 84816
rect 263100 84804 263106 84856
rect 95050 84124 95056 84176
rect 95108 84164 95114 84176
rect 231302 84164 231308 84176
rect 95108 84136 231308 84164
rect 95108 84124 95114 84136
rect 231302 84124 231308 84136
rect 231360 84124 231366 84176
rect 97902 84056 97908 84108
rect 97960 84096 97966 84108
rect 180242 84096 180248 84108
rect 97960 84068 180248 84096
rect 97960 84056 97966 84068
rect 180242 84056 180248 84068
rect 180300 84056 180306 84108
rect 255958 83512 255964 83564
rect 256016 83552 256022 83564
rect 276934 83552 276940 83564
rect 256016 83524 276940 83552
rect 256016 83512 256022 83524
rect 276934 83512 276940 83524
rect 276992 83512 276998 83564
rect 221458 83444 221464 83496
rect 221516 83484 221522 83496
rect 295978 83484 295984 83496
rect 221516 83456 295984 83484
rect 221516 83444 221522 83456
rect 295978 83444 295984 83456
rect 296036 83444 296042 83496
rect 96522 82764 96528 82816
rect 96580 82804 96586 82816
rect 211798 82804 211804 82816
rect 96580 82776 211804 82804
rect 96580 82764 96586 82776
rect 211798 82764 211804 82776
rect 211856 82764 211862 82816
rect 114278 82696 114284 82748
rect 114336 82736 114342 82748
rect 167638 82736 167644 82748
rect 114336 82708 167644 82736
rect 114336 82696 114342 82708
rect 167638 82696 167644 82708
rect 167696 82696 167702 82748
rect 95142 81336 95148 81388
rect 95200 81376 95206 81388
rect 234154 81376 234160 81388
rect 95200 81348 234160 81376
rect 95200 81336 95206 81348
rect 234154 81336 234160 81348
rect 234212 81336 234218 81388
rect 151078 81268 151084 81320
rect 151136 81308 151142 81320
rect 162210 81308 162216 81320
rect 151136 81280 162216 81308
rect 151136 81268 151142 81280
rect 162210 81268 162216 81280
rect 162268 81268 162274 81320
rect 162118 80656 162124 80708
rect 162176 80696 162182 80708
rect 264330 80696 264336 80708
rect 162176 80668 264336 80696
rect 162176 80656 162182 80668
rect 264330 80656 264336 80668
rect 264388 80656 264394 80708
rect 122190 79976 122196 80028
rect 122248 80016 122254 80028
rect 163498 80016 163504 80028
rect 122248 79988 163504 80016
rect 122248 79976 122254 79988
rect 163498 79976 163504 79988
rect 163556 79976 163562 80028
rect 151722 79908 151728 79960
rect 151780 79948 151786 79960
rect 178770 79948 178776 79960
rect 151780 79920 178776 79948
rect 151780 79908 151786 79920
rect 178770 79908 178776 79920
rect 178828 79908 178834 79960
rect 88978 78616 88984 78668
rect 89036 78656 89042 78668
rect 200758 78656 200764 78668
rect 89036 78628 200764 78656
rect 89036 78616 89042 78628
rect 200758 78616 200764 78628
rect 200816 78616 200822 78668
rect 324958 78616 324964 78668
rect 325016 78656 325022 78668
rect 325694 78656 325700 78668
rect 325016 78628 325700 78656
rect 325016 78616 325022 78628
rect 325694 78616 325700 78628
rect 325752 78616 325758 78668
rect 125502 78548 125508 78600
rect 125560 78588 125566 78600
rect 170398 78588 170404 78600
rect 125560 78560 170404 78588
rect 125560 78548 125566 78560
rect 170398 78548 170404 78560
rect 170456 78548 170462 78600
rect 229738 77936 229744 77988
rect 229796 77976 229802 77988
rect 275278 77976 275284 77988
rect 229796 77948 275284 77976
rect 229796 77936 229802 77948
rect 275278 77936 275284 77948
rect 275336 77936 275342 77988
rect 91002 77188 91008 77240
rect 91060 77228 91066 77240
rect 167730 77228 167736 77240
rect 91060 77200 167736 77228
rect 91060 77188 91066 77200
rect 167730 77188 167736 77200
rect 167788 77188 167794 77240
rect 118510 77120 118516 77172
rect 118568 77160 118574 77172
rect 181438 77160 181444 77172
rect 118568 77132 181444 77160
rect 118568 77120 118574 77132
rect 181438 77120 181444 77132
rect 181496 77120 181502 77172
rect 121362 75828 121368 75880
rect 121420 75868 121426 75880
rect 173434 75868 173440 75880
rect 121420 75840 173440 75868
rect 121420 75828 121426 75840
rect 173434 75828 173440 75840
rect 173492 75828 173498 75880
rect 97902 75148 97908 75200
rect 97960 75188 97966 75200
rect 278222 75188 278228 75200
rect 97960 75160 278228 75188
rect 97960 75148 97966 75160
rect 278222 75148 278228 75160
rect 278280 75148 278286 75200
rect 116578 74468 116584 74520
rect 116636 74508 116642 74520
rect 214650 74508 214656 74520
rect 116636 74480 214656 74508
rect 116636 74468 116642 74480
rect 214650 74468 214656 74480
rect 214708 74468 214714 74520
rect 153102 74400 153108 74452
rect 153160 74440 153166 74452
rect 233970 74440 233976 74452
rect 153160 74412 233976 74440
rect 153160 74400 153166 74412
rect 233970 74400 233976 74412
rect 234028 74400 234034 74452
rect 86770 73788 86776 73840
rect 86828 73828 86834 73840
rect 105538 73828 105544 73840
rect 86828 73800 105544 73828
rect 86828 73788 86834 73800
rect 105538 73788 105544 73800
rect 105596 73788 105602 73840
rect 100018 73108 100024 73160
rect 100076 73148 100082 73160
rect 209130 73148 209136 73160
rect 100076 73120 209136 73148
rect 100076 73108 100082 73120
rect 209130 73108 209136 73120
rect 209188 73108 209194 73160
rect 124122 73040 124128 73092
rect 124180 73080 124186 73092
rect 174630 73080 174636 73092
rect 124180 73052 174636 73080
rect 124180 73040 124186 73052
rect 174630 73040 174636 73052
rect 174688 73040 174694 73092
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 18598 71720 18604 71732
rect 3476 71692 18604 71720
rect 3476 71680 3482 71692
rect 18598 71680 18604 71692
rect 18656 71680 18662 71732
rect 119982 71680 119988 71732
rect 120040 71720 120046 71732
rect 177390 71720 177396 71732
rect 120040 71692 177396 71720
rect 120040 71680 120046 71692
rect 177390 71680 177396 71692
rect 177448 71680 177454 71732
rect 113082 71000 113088 71052
rect 113140 71040 113146 71052
rect 274082 71040 274088 71052
rect 113140 71012 274088 71040
rect 113140 71000 113146 71012
rect 274082 71000 274088 71012
rect 274140 71000 274146 71052
rect 129642 70320 129648 70372
rect 129700 70360 129706 70372
rect 175918 70360 175924 70372
rect 129700 70332 175924 70360
rect 129700 70320 129706 70332
rect 175918 70320 175924 70332
rect 175976 70320 175982 70372
rect 119982 69640 119988 69692
rect 120040 69680 120046 69692
rect 272702 69680 272708 69692
rect 120040 69652 272708 69680
rect 120040 69640 120046 69652
rect 272702 69640 272708 69652
rect 272760 69640 272766 69692
rect 108850 68960 108856 69012
rect 108908 69000 108914 69012
rect 184382 69000 184388 69012
rect 108908 68972 184388 69000
rect 108908 68960 108914 68972
rect 184382 68960 184388 68972
rect 184440 68960 184446 69012
rect 133782 68892 133788 68944
rect 133840 68932 133846 68944
rect 197998 68932 198004 68944
rect 133840 68904 198004 68932
rect 133840 68892 133846 68904
rect 197998 68892 198004 68904
rect 198056 68892 198062 68944
rect 110322 67532 110328 67584
rect 110380 67572 110386 67584
rect 170582 67572 170588 67584
rect 110380 67544 170588 67572
rect 110380 67532 110386 67544
rect 170582 67532 170588 67544
rect 170640 67532 170646 67584
rect 71038 66852 71044 66904
rect 71096 66892 71102 66904
rect 245010 66892 245016 66904
rect 71096 66864 245016 66892
rect 71096 66852 71102 66864
rect 245010 66852 245016 66864
rect 245068 66852 245074 66904
rect 112990 66172 112996 66224
rect 113048 66212 113054 66224
rect 186958 66212 186964 66224
rect 113048 66184 186964 66212
rect 113048 66172 113054 66184
rect 186958 66172 186964 66184
rect 187016 66172 187022 66224
rect 106918 66104 106924 66156
rect 106976 66144 106982 66156
rect 171870 66144 171876 66156
rect 106976 66116 171876 66144
rect 106976 66104 106982 66116
rect 171870 66104 171876 66116
rect 171928 66104 171934 66156
rect 251818 65492 251824 65544
rect 251876 65532 251882 65544
rect 268654 65532 268660 65544
rect 251876 65504 268660 65532
rect 251876 65492 251882 65504
rect 268654 65492 268660 65504
rect 268712 65492 268718 65544
rect 88150 64812 88156 64864
rect 88208 64852 88214 64864
rect 199470 64852 199476 64864
rect 88208 64824 199476 64852
rect 88208 64812 88214 64824
rect 199470 64812 199476 64824
rect 199528 64812 199534 64864
rect 103422 64744 103428 64796
rect 103480 64784 103486 64796
rect 213270 64784 213276 64796
rect 103480 64756 213276 64784
rect 103480 64744 103486 64756
rect 213270 64744 213276 64756
rect 213328 64744 213334 64796
rect 126698 63452 126704 63504
rect 126756 63492 126762 63504
rect 220170 63492 220176 63504
rect 126756 63464 220176 63492
rect 126756 63452 126762 63464
rect 220170 63452 220176 63464
rect 220228 63452 220234 63504
rect 104802 63384 104808 63436
rect 104860 63424 104866 63436
rect 178862 63424 178868 63436
rect 104860 63396 178868 63424
rect 104860 63384 104866 63396
rect 178862 63384 178868 63396
rect 178920 63384 178926 63436
rect 115842 62024 115848 62076
rect 115900 62064 115906 62076
rect 238018 62064 238024 62076
rect 115900 62036 238024 62064
rect 115900 62024 115906 62036
rect 238018 62024 238024 62036
rect 238076 62024 238082 62076
rect 59170 61344 59176 61396
rect 59228 61384 59234 61396
rect 274174 61384 274180 61396
rect 59228 61356 274180 61384
rect 59228 61344 59234 61356
rect 274174 61344 274180 61356
rect 274232 61344 274238 61396
rect 105538 60664 105544 60716
rect 105596 60704 105602 60716
rect 203518 60704 203524 60716
rect 105596 60676 203524 60704
rect 105596 60664 105602 60676
rect 203518 60664 203524 60676
rect 203576 60664 203582 60716
rect 128998 60596 129004 60648
rect 129056 60636 129062 60648
rect 191190 60636 191196 60648
rect 129056 60608 191196 60636
rect 129056 60596 129062 60608
rect 191190 60596 191196 60608
rect 191248 60596 191254 60648
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 17218 59344 17224 59356
rect 3108 59316 17224 59344
rect 3108 59304 3114 59316
rect 17218 59304 17224 59316
rect 17276 59304 17282 59356
rect 108942 59304 108948 59356
rect 109000 59344 109006 59356
rect 202322 59344 202328 59356
rect 109000 59316 202328 59344
rect 109000 59304 109006 59316
rect 202322 59304 202328 59316
rect 202380 59304 202386 59356
rect 126790 59236 126796 59288
rect 126848 59276 126854 59288
rect 188430 59276 188436 59288
rect 126848 59248 188436 59276
rect 126848 59236 126854 59248
rect 188430 59236 188436 59248
rect 188488 59236 188494 59288
rect 214650 58624 214656 58676
rect 214708 58664 214714 58676
rect 235994 58664 236000 58676
rect 214708 58636 236000 58664
rect 214708 58624 214714 58636
rect 235994 58624 236000 58636
rect 236052 58624 236058 58676
rect 101950 57876 101956 57928
rect 102008 57916 102014 57928
rect 195330 57916 195336 57928
rect 102008 57888 195336 57916
rect 102008 57876 102014 57888
rect 195330 57876 195336 57888
rect 195388 57876 195394 57928
rect 77202 57196 77208 57248
rect 77260 57236 77266 57248
rect 280982 57236 280988 57248
rect 77260 57208 280988 57236
rect 77260 57196 77266 57208
rect 280982 57196 280988 57208
rect 281040 57196 281046 57248
rect 126882 56516 126888 56568
rect 126940 56556 126946 56568
rect 242250 56556 242256 56568
rect 126940 56528 242256 56556
rect 126940 56516 126946 56528
rect 242250 56516 242256 56528
rect 242308 56516 242314 56568
rect 91002 55836 91008 55888
rect 91060 55876 91066 55888
rect 267182 55876 267188 55888
rect 91060 55848 267188 55876
rect 91060 55836 91066 55848
rect 267182 55836 267188 55848
rect 267240 55836 267246 55888
rect 102042 55156 102048 55208
rect 102100 55196 102106 55208
rect 244918 55196 244924 55208
rect 102100 55168 244924 55196
rect 102100 55156 102106 55168
rect 244918 55156 244924 55168
rect 244976 55156 244982 55208
rect 95050 54476 95056 54528
rect 95108 54516 95114 54528
rect 286318 54516 286324 54528
rect 95108 54488 286324 54516
rect 95108 54476 95114 54488
rect 286318 54476 286324 54488
rect 286376 54476 286382 54528
rect 118602 53728 118608 53780
rect 118660 53768 118666 53780
rect 239398 53768 239404 53780
rect 118660 53740 239404 53768
rect 118660 53728 118666 53740
rect 239398 53728 239404 53740
rect 239456 53728 239462 53780
rect 102042 53048 102048 53100
rect 102100 53088 102106 53100
rect 273990 53088 273996 53100
rect 102100 53060 273996 53088
rect 102100 53048 102106 53060
rect 273990 53048 273996 53060
rect 274048 53048 274054 53100
rect 117222 52368 117228 52420
rect 117280 52408 117286 52420
rect 225598 52408 225604 52420
rect 117280 52380 225604 52408
rect 117280 52368 117286 52380
rect 225598 52368 225604 52380
rect 225656 52368 225662 52420
rect 104802 51688 104808 51740
rect 104860 51728 104866 51740
rect 283558 51728 283564 51740
rect 104860 51700 283564 51728
rect 104860 51688 104866 51700
rect 283558 51688 283564 51700
rect 283616 51688 283622 51740
rect 174538 50396 174544 50448
rect 174596 50436 174602 50448
rect 273254 50436 273260 50448
rect 174596 50408 273260 50436
rect 174596 50396 174602 50408
rect 273254 50396 273260 50408
rect 273312 50396 273318 50448
rect 86862 50328 86868 50380
rect 86920 50368 86926 50380
rect 289078 50368 289084 50380
rect 86920 50340 289084 50368
rect 86920 50328 86926 50340
rect 289078 50328 289084 50340
rect 289136 50328 289142 50380
rect 107562 49036 107568 49088
rect 107620 49076 107626 49088
rect 250530 49076 250536 49088
rect 107620 49048 250536 49076
rect 107620 49036 107626 49048
rect 250530 49036 250536 49048
rect 250588 49036 250594 49088
rect 37182 48968 37188 49020
rect 37240 49008 37246 49020
rect 276750 49008 276756 49020
rect 37240 48980 276756 49008
rect 37240 48968 37246 48980
rect 276750 48968 276756 48980
rect 276808 48968 276814 49020
rect 71682 47608 71688 47660
rect 71740 47648 71746 47660
rect 265802 47648 265808 47660
rect 71740 47620 265808 47648
rect 71740 47608 71746 47620
rect 265802 47608 265808 47620
rect 265860 47608 265866 47660
rect 39942 47540 39948 47592
rect 40000 47580 40006 47592
rect 236638 47580 236644 47592
rect 40000 47552 236644 47580
rect 40000 47540 40006 47552
rect 236638 47540 236644 47552
rect 236696 47540 236702 47592
rect 238018 47540 238024 47592
rect 238076 47580 238082 47592
rect 249058 47580 249064 47592
rect 238076 47552 249064 47580
rect 238076 47540 238082 47552
rect 249058 47540 249064 47552
rect 249116 47540 249122 47592
rect 119890 46248 119896 46300
rect 119948 46288 119954 46300
rect 268562 46288 268568 46300
rect 119948 46260 268568 46288
rect 119948 46248 119954 46260
rect 268562 46248 268568 46260
rect 268620 46248 268626 46300
rect 126238 46180 126244 46232
rect 126296 46220 126302 46232
rect 282362 46220 282368 46232
rect 126296 46192 282368 46220
rect 126296 46180 126302 46192
rect 282362 46180 282368 46192
rect 282420 46180 282426 46232
rect 2774 45500 2780 45552
rect 2832 45540 2838 45552
rect 4798 45540 4804 45552
rect 2832 45512 4804 45540
rect 2832 45500 2838 45512
rect 4798 45500 4804 45512
rect 4856 45500 4862 45552
rect 115842 44820 115848 44872
rect 115900 44860 115906 44872
rect 260190 44860 260196 44872
rect 115900 44832 260196 44860
rect 115900 44820 115906 44832
rect 260190 44820 260196 44832
rect 260248 44820 260254 44872
rect 84102 43460 84108 43512
rect 84160 43500 84166 43512
rect 271322 43500 271328 43512
rect 84160 43472 271328 43500
rect 84160 43460 84166 43472
rect 271322 43460 271328 43472
rect 271380 43460 271386 43512
rect 75822 43392 75828 43444
rect 75880 43432 75886 43444
rect 283650 43432 283656 43444
rect 75880 43404 283656 43432
rect 75880 43392 75886 43404
rect 283650 43392 283656 43404
rect 283708 43392 283714 43444
rect 12250 42100 12256 42152
rect 12308 42140 12314 42152
rect 272610 42140 272616 42152
rect 12308 42112 272616 42140
rect 12308 42100 12314 42112
rect 272610 42100 272616 42112
rect 272668 42100 272674 42152
rect 5442 42032 5448 42084
rect 5500 42072 5506 42084
rect 291194 42072 291200 42084
rect 5500 42044 291200 42072
rect 5500 42032 5506 42044
rect 291194 42032 291200 42044
rect 291252 42032 291258 42084
rect 205082 40740 205088 40792
rect 205140 40780 205146 40792
rect 214650 40780 214656 40792
rect 205140 40752 214656 40780
rect 205140 40740 205146 40752
rect 214650 40740 214656 40752
rect 214708 40740 214714 40792
rect 217318 40740 217324 40792
rect 217376 40780 217382 40792
rect 291194 40780 291200 40792
rect 217376 40752 291200 40780
rect 217376 40740 217382 40752
rect 291194 40740 291200 40752
rect 291252 40740 291258 40792
rect 57238 40672 57244 40724
rect 57296 40712 57302 40724
rect 253198 40712 253204 40724
rect 57296 40684 253204 40712
rect 57296 40672 57302 40684
rect 253198 40672 253204 40684
rect 253256 40672 253262 40724
rect 74442 39380 74448 39432
rect 74500 39420 74506 39432
rect 160738 39420 160744 39432
rect 74500 39392 160744 39420
rect 74500 39380 74506 39392
rect 160738 39380 160744 39392
rect 160796 39380 160802 39432
rect 213178 39380 213184 39432
rect 213236 39420 213242 39432
rect 276014 39420 276020 39432
rect 213236 39392 276020 39420
rect 213236 39380 213242 39392
rect 276014 39380 276020 39392
rect 276072 39380 276078 39432
rect 146938 39312 146944 39364
rect 146996 39352 147002 39364
rect 260098 39352 260104 39364
rect 146996 39324 260104 39352
rect 146996 39312 147002 39324
rect 260098 39312 260104 39324
rect 260156 39312 260162 39364
rect 55030 37884 55036 37936
rect 55088 37924 55094 37936
rect 282270 37924 282276 37936
rect 55088 37896 282276 37924
rect 55088 37884 55094 37896
rect 282270 37884 282276 37896
rect 282328 37884 282334 37936
rect 79318 36592 79324 36644
rect 79376 36632 79382 36644
rect 251818 36632 251824 36644
rect 79376 36604 251824 36632
rect 79376 36592 79382 36604
rect 251818 36592 251824 36604
rect 251876 36592 251882 36644
rect 3970 36524 3976 36576
rect 4028 36564 4034 36576
rect 262858 36564 262864 36576
rect 4028 36536 262864 36564
rect 4028 36524 4034 36536
rect 262858 36524 262864 36536
rect 262916 36524 262922 36576
rect 204898 35232 204904 35284
rect 204956 35272 204962 35284
rect 287054 35272 287060 35284
rect 204956 35244 287060 35272
rect 204956 35232 204962 35244
rect 287054 35232 287060 35244
rect 287112 35232 287118 35284
rect 1394 35164 1400 35216
rect 1452 35204 1458 35216
rect 229830 35204 229836 35216
rect 1452 35176 229836 35204
rect 1452 35164 1458 35176
rect 229830 35164 229836 35176
rect 229888 35164 229894 35216
rect 142798 33804 142804 33856
rect 142856 33844 142862 33856
rect 206278 33844 206284 33856
rect 142856 33816 206284 33844
rect 142856 33804 142862 33816
rect 206278 33804 206284 33816
rect 206336 33804 206342 33856
rect 41322 33736 41328 33788
rect 41380 33776 41386 33788
rect 147030 33776 147036 33788
rect 41380 33748 147036 33776
rect 41380 33736 41386 33748
rect 147030 33736 147036 33748
rect 147088 33736 147094 33788
rect 199378 33736 199384 33788
rect 199436 33776 199442 33788
rect 269114 33776 269120 33788
rect 199436 33748 269120 33776
rect 199436 33736 199442 33748
rect 269114 33736 269120 33748
rect 269172 33736 269178 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 39298 33096 39304 33108
rect 3568 33068 39304 33096
rect 3568 33056 3574 33068
rect 39298 33056 39304 33068
rect 39356 33056 39362 33108
rect 189718 32444 189724 32496
rect 189776 32484 189782 32496
rect 271322 32484 271328 32496
rect 189776 32456 271328 32484
rect 189776 32444 189782 32456
rect 271322 32444 271328 32456
rect 271380 32444 271386 32496
rect 124122 32376 124128 32428
rect 124180 32416 124186 32428
rect 280798 32416 280804 32428
rect 124180 32388 280804 32416
rect 124180 32376 124186 32388
rect 280798 32376 280804 32388
rect 280856 32376 280862 32428
rect 196618 31084 196624 31136
rect 196676 31124 196682 31136
rect 259454 31124 259460 31136
rect 196676 31096 259460 31124
rect 196676 31084 196682 31096
rect 259454 31084 259460 31096
rect 259512 31084 259518 31136
rect 118602 31016 118608 31068
rect 118660 31056 118666 31068
rect 232590 31056 232596 31068
rect 118660 31028 232596 31056
rect 118660 31016 118666 31028
rect 232590 31016 232596 31028
rect 232648 31016 232654 31068
rect 122742 29656 122748 29708
rect 122800 29696 122806 29708
rect 198090 29696 198096 29708
rect 122800 29668 198096 29696
rect 122800 29656 122806 29668
rect 198090 29656 198096 29668
rect 198148 29656 198154 29708
rect 185578 29588 185584 29640
rect 185636 29628 185642 29640
rect 267734 29628 267740 29640
rect 185636 29600 267740 29628
rect 185636 29588 185642 29600
rect 267734 29588 267740 29600
rect 267792 29588 267798 29640
rect 130378 28296 130384 28348
rect 130436 28336 130442 28348
rect 168374 28336 168380 28348
rect 130436 28308 168380 28336
rect 130436 28296 130442 28308
rect 168374 28296 168380 28308
rect 168432 28296 168438 28348
rect 182818 28296 182824 28348
rect 182876 28336 182882 28348
rect 271414 28336 271420 28348
rect 182876 28308 271420 28336
rect 182876 28296 182882 28308
rect 271414 28296 271420 28308
rect 271472 28296 271478 28348
rect 53650 28228 53656 28280
rect 53708 28268 53714 28280
rect 279510 28268 279516 28280
rect 53708 28240 279516 28268
rect 53708 28228 53714 28240
rect 279510 28228 279516 28240
rect 279568 28228 279574 28280
rect 114554 26936 114560 26988
rect 114612 26976 114618 26988
rect 205082 26976 205088 26988
rect 114612 26948 205088 26976
rect 114612 26936 114618 26948
rect 205082 26936 205088 26948
rect 205140 26936 205146 26988
rect 44082 26868 44088 26920
rect 44140 26908 44146 26920
rect 151078 26908 151084 26920
rect 44140 26880 151084 26908
rect 44140 26868 44146 26880
rect 151078 26868 151084 26880
rect 151136 26868 151142 26920
rect 204990 26868 204996 26920
rect 205048 26908 205054 26920
rect 263594 26908 263600 26920
rect 205048 26880 263600 26908
rect 205048 26868 205054 26880
rect 263594 26868 263600 26880
rect 263652 26868 263658 26920
rect 209038 25576 209044 25628
rect 209096 25616 209102 25628
rect 295334 25616 295340 25628
rect 209096 25588 295340 25616
rect 209096 25576 209102 25588
rect 295334 25576 295340 25588
rect 295392 25576 295398 25628
rect 96522 25508 96528 25560
rect 96580 25548 96586 25560
rect 271230 25548 271236 25560
rect 96580 25520 271236 25548
rect 96580 25508 96586 25520
rect 271230 25508 271236 25520
rect 271288 25508 271294 25560
rect 117222 24148 117228 24200
rect 117280 24188 117286 24200
rect 268470 24188 268476 24200
rect 117280 24160 268476 24188
rect 117280 24148 117286 24160
rect 268470 24148 268476 24160
rect 268528 24148 268534 24200
rect 81342 24080 81348 24132
rect 81400 24120 81406 24132
rect 264238 24120 264244 24132
rect 81400 24092 264244 24120
rect 81400 24080 81406 24092
rect 264238 24080 264244 24092
rect 264296 24080 264302 24132
rect 111610 22788 111616 22840
rect 111668 22828 111674 22840
rect 278038 22828 278044 22840
rect 111668 22800 278044 22828
rect 111668 22788 111674 22800
rect 278038 22788 278044 22800
rect 278096 22788 278102 22840
rect 56502 22720 56508 22772
rect 56560 22760 56566 22772
rect 276658 22760 276664 22772
rect 56560 22732 276664 22760
rect 56560 22720 56566 22732
rect 276658 22720 276664 22732
rect 276716 22720 276722 22772
rect 125502 21428 125508 21480
rect 125560 21468 125566 21480
rect 267090 21468 267096 21480
rect 125560 21440 267096 21468
rect 125560 21428 125566 21440
rect 267090 21428 267096 21440
rect 267148 21428 267154 21480
rect 50982 21360 50988 21412
rect 51040 21400 51046 21412
rect 251266 21400 251272 21412
rect 51040 21372 251272 21400
rect 51040 21360 51046 21372
rect 251266 21360 251272 21372
rect 251324 21360 251330 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 36538 20652 36544 20664
rect 3476 20624 36544 20652
rect 3476 20612 3482 20624
rect 36538 20612 36544 20624
rect 36596 20612 36602 20664
rect 112438 20136 112444 20188
rect 112496 20176 112502 20188
rect 114554 20176 114560 20188
rect 112496 20148 114560 20176
rect 112496 20136 112502 20148
rect 114554 20136 114560 20148
rect 114612 20136 114618 20188
rect 188338 20000 188344 20052
rect 188396 20040 188402 20052
rect 242894 20040 242900 20052
rect 188396 20012 242900 20040
rect 188396 20000 188402 20012
rect 242894 20000 242900 20012
rect 242952 20000 242958 20052
rect 49602 19932 49608 19984
rect 49660 19972 49666 19984
rect 266998 19972 267004 19984
rect 49660 19944 267004 19972
rect 49660 19932 49666 19944
rect 266998 19932 267004 19944
rect 267056 19932 267062 19984
rect 178678 18640 178684 18692
rect 178736 18680 178742 18692
rect 281534 18680 281540 18692
rect 178736 18652 281540 18680
rect 178736 18640 178742 18652
rect 281534 18640 281540 18652
rect 281592 18640 281598 18692
rect 60642 18572 60648 18624
rect 60700 18612 60706 18624
rect 238018 18612 238024 18624
rect 60700 18584 238024 18612
rect 60700 18572 60706 18584
rect 238018 18572 238024 18584
rect 238076 18572 238082 18624
rect 14 17280 20 17332
rect 72 17320 78 17332
rect 116578 17320 116584 17332
rect 72 17292 116584 17320
rect 72 17280 78 17292
rect 116578 17280 116584 17292
rect 116636 17280 116642 17332
rect 236638 17280 236644 17332
rect 236696 17320 236702 17332
rect 347038 17320 347044 17332
rect 236696 17292 347044 17320
rect 236696 17280 236702 17292
rect 347038 17280 347044 17292
rect 347096 17280 347102 17332
rect 106918 17212 106924 17264
rect 106976 17252 106982 17264
rect 238018 17252 238024 17264
rect 106976 17224 238024 17252
rect 106976 17212 106982 17224
rect 238018 17212 238024 17224
rect 238076 17212 238082 17264
rect 68922 15920 68928 15972
rect 68980 15960 68986 15972
rect 104158 15960 104164 15972
rect 68980 15932 104164 15960
rect 68980 15920 68986 15932
rect 104158 15920 104164 15932
rect 104216 15920 104222 15972
rect 240778 15920 240784 15972
rect 240836 15960 240842 15972
rect 264974 15960 264980 15972
rect 240836 15932 264980 15960
rect 240836 15920 240842 15932
rect 264974 15920 264980 15932
rect 265032 15920 265038 15972
rect 35158 15852 35164 15904
rect 35216 15892 35222 15904
rect 79318 15892 79324 15904
rect 35216 15864 79324 15892
rect 35216 15852 35222 15864
rect 79318 15852 79324 15864
rect 79376 15852 79382 15904
rect 88978 15852 88984 15904
rect 89036 15892 89042 15904
rect 246298 15892 246304 15904
rect 89036 15864 246304 15892
rect 89036 15852 89042 15864
rect 246298 15852 246304 15864
rect 246356 15852 246362 15904
rect 9582 14492 9588 14544
rect 9640 14532 9646 14544
rect 224218 14532 224224 14544
rect 9640 14504 224224 14532
rect 9640 14492 9646 14504
rect 224218 14492 224224 14504
rect 224276 14492 224282 14544
rect 63402 14424 63408 14476
rect 63460 14464 63466 14476
rect 314654 14464 314660 14476
rect 63460 14436 314660 14464
rect 63460 14424 63466 14436
rect 314654 14424 314660 14436
rect 314712 14424 314718 14476
rect 92382 13132 92388 13184
rect 92440 13172 92446 13184
rect 272518 13172 272524 13184
rect 92440 13144 272524 13172
rect 92440 13132 92446 13144
rect 272518 13132 272524 13144
rect 272576 13132 272582 13184
rect 23014 13064 23020 13116
rect 23072 13104 23078 13116
rect 214558 13104 214564 13116
rect 23072 13076 214564 13104
rect 23072 13064 23078 13076
rect 214558 13064 214564 13076
rect 214616 13064 214622 13116
rect 110322 11772 110328 11824
rect 110380 11812 110386 11824
rect 269758 11812 269764 11824
rect 110380 11784 269764 11812
rect 110380 11772 110386 11784
rect 269758 11772 269764 11784
rect 269816 11772 269822 11824
rect 36998 11704 37004 11756
rect 37056 11744 37062 11756
rect 269850 11744 269856 11756
rect 37056 11716 269856 11744
rect 37056 11704 37062 11716
rect 269850 11704 269856 11716
rect 269908 11704 269914 11756
rect 108942 10344 108948 10396
rect 109000 10384 109006 10396
rect 142798 10384 142804 10396
rect 109000 10356 142804 10384
rect 109000 10344 109006 10356
rect 142798 10344 142804 10356
rect 142856 10344 142862 10396
rect 202138 10344 202144 10396
rect 202196 10384 202202 10396
rect 284938 10384 284944 10396
rect 202196 10356 284944 10384
rect 202196 10344 202202 10356
rect 284938 10344 284944 10356
rect 284996 10344 285002 10396
rect 31294 10276 31300 10328
rect 31352 10316 31358 10328
rect 255958 10316 255964 10328
rect 31352 10288 255964 10316
rect 31352 10276 31358 10288
rect 255958 10276 255964 10288
rect 256016 10276 256022 10328
rect 9950 8984 9956 9036
rect 10008 9024 10014 9036
rect 162118 9024 162124 9036
rect 10008 8996 162124 9024
rect 10008 8984 10014 8996
rect 162118 8984 162124 8996
rect 162176 8984 162182 9036
rect 66714 8916 66720 8968
rect 66772 8956 66778 8968
rect 254578 8956 254584 8968
rect 66772 8928 254584 8956
rect 66772 8916 66778 8928
rect 254578 8916 254584 8928
rect 254636 8916 254642 8968
rect 44266 7624 44272 7676
rect 44324 7664 44330 7676
rect 71038 7664 71044 7676
rect 44324 7636 71044 7664
rect 44324 7624 44330 7636
rect 71038 7624 71044 7636
rect 71096 7624 71102 7676
rect 92750 7624 92756 7676
rect 92808 7664 92814 7676
rect 271138 7664 271144 7676
rect 92808 7636 271144 7664
rect 92808 7624 92814 7636
rect 271138 7624 271144 7636
rect 271196 7624 271202 7676
rect 61930 7556 61936 7608
rect 61988 7596 61994 7608
rect 268286 7596 268292 7608
rect 61988 7568 268292 7596
rect 61988 7556 61994 7568
rect 268286 7556 268292 7568
rect 268344 7556 268350 7608
rect 3418 6604 3424 6656
rect 3476 6644 3482 6656
rect 7558 6644 7564 6656
rect 3476 6616 7564 6644
rect 3476 6604 3482 6616
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 89162 6196 89168 6248
rect 89220 6236 89226 6248
rect 112438 6236 112444 6248
rect 89220 6208 112444 6236
rect 89220 6196 89226 6208
rect 112438 6196 112444 6208
rect 112496 6196 112502 6248
rect 114002 6196 114008 6248
rect 114060 6236 114066 6248
rect 279418 6236 279424 6248
rect 114060 6208 279424 6236
rect 114060 6196 114066 6208
rect 279418 6196 279424 6208
rect 279476 6196 279482 6248
rect 30098 6128 30104 6180
rect 30156 6168 30162 6180
rect 196802 6168 196808 6180
rect 30156 6140 196808 6168
rect 30156 6128 30162 6140
rect 196802 6128 196808 6140
rect 196860 6128 196866 6180
rect 233878 6128 233884 6180
rect 233936 6168 233942 6180
rect 260650 6168 260656 6180
rect 233936 6140 260656 6168
rect 233936 6128 233942 6140
rect 260650 6128 260656 6140
rect 260708 6128 260714 6180
rect 304258 6128 304264 6180
rect 304316 6168 304322 6180
rect 342162 6168 342168 6180
rect 304316 6140 342168 6168
rect 304316 6128 304322 6140
rect 342162 6128 342168 6140
rect 342220 6128 342226 6180
rect 69106 4836 69112 4888
rect 69164 4876 69170 4888
rect 146938 4876 146944 4888
rect 69164 4848 146944 4876
rect 69164 4836 69170 4848
rect 146938 4836 146944 4848
rect 146996 4836 147002 4888
rect 184198 4836 184204 4888
rect 184256 4876 184262 4888
rect 303154 4876 303160 4888
rect 184256 4848 303160 4876
rect 184256 4836 184262 4848
rect 303154 4836 303160 4848
rect 303212 4836 303218 4888
rect 11146 4768 11152 4820
rect 11204 4808 11210 4820
rect 35158 4808 35164 4820
rect 11204 4780 35164 4808
rect 11204 4768 11210 4780
rect 35158 4768 35164 4780
rect 35216 4768 35222 4820
rect 45462 4768 45468 4820
rect 45520 4808 45526 4820
rect 291286 4808 291292 4820
rect 45520 4780 291292 4808
rect 45520 4768 45526 4780
rect 291286 4768 291292 4780
rect 291344 4768 291350 4820
rect 338666 4768 338672 4820
rect 338724 4808 338730 4820
rect 360194 4808 360200 4820
rect 338724 4780 360200 4808
rect 338724 4768 338730 4780
rect 360194 4768 360200 4780
rect 360252 4768 360258 4820
rect 27706 3612 27712 3664
rect 27764 3652 27770 3664
rect 28902 3652 28908 3664
rect 27764 3624 28908 3652
rect 27764 3612 27770 3624
rect 28902 3612 28908 3624
rect 28960 3612 28966 3664
rect 35986 3544 35992 3596
rect 36044 3584 36050 3596
rect 37090 3584 37096 3596
rect 36044 3556 37096 3584
rect 36044 3544 36050 3556
rect 37090 3544 37096 3556
rect 37148 3544 37154 3596
rect 51350 3544 51356 3596
rect 51408 3584 51414 3596
rect 57146 3584 57152 3596
rect 51408 3556 57152 3584
rect 51408 3544 51414 3556
rect 57146 3544 57152 3556
rect 57204 3544 57210 3596
rect 60826 3544 60832 3596
rect 60884 3584 60890 3596
rect 62022 3584 62028 3596
rect 60884 3556 62028 3584
rect 60884 3544 60890 3556
rect 62022 3544 62028 3556
rect 62080 3544 62086 3596
rect 102226 3544 102232 3596
rect 102284 3584 102290 3596
rect 122098 3584 122104 3596
rect 102284 3556 122104 3584
rect 102284 3544 102290 3556
rect 122098 3544 122104 3556
rect 122156 3544 122162 3596
rect 228358 3544 228364 3596
rect 228416 3584 228422 3596
rect 239306 3584 239312 3596
rect 228416 3556 239312 3584
rect 228416 3544 228422 3556
rect 239306 3544 239312 3556
rect 239364 3544 239370 3596
rect 251174 3544 251180 3596
rect 251232 3584 251238 3596
rect 252370 3584 252376 3596
rect 251232 3556 252376 3584
rect 251232 3544 251238 3556
rect 252370 3544 252376 3556
rect 252428 3544 252434 3596
rect 299566 3544 299572 3596
rect 299624 3584 299630 3596
rect 300762 3584 300768 3596
rect 299624 3556 300768 3584
rect 299624 3544 299630 3556
rect 300762 3544 300768 3556
rect 300820 3544 300826 3596
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3970 3516 3976 3528
rect 2924 3488 3976 3516
rect 2924 3476 2930 3488
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 9582 3516 9588 3528
rect 8812 3488 9588 3516
rect 8812 3476 8818 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 16482 3516 16488 3528
rect 15988 3488 16488 3516
rect 15988 3476 15994 3488
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 19242 3516 19248 3528
rect 18288 3488 19248 3516
rect 18288 3476 18294 3488
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 20622 3476 20628 3528
rect 20680 3516 20686 3528
rect 22738 3516 22744 3528
rect 20680 3488 22744 3516
rect 20680 3476 20686 3488
rect 22738 3476 22744 3488
rect 22796 3476 22802 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 24762 3516 24768 3528
rect 24268 3488 24768 3516
rect 24268 3476 24274 3488
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 25314 3476 25320 3528
rect 25372 3516 25378 3528
rect 26142 3516 26148 3528
rect 25372 3488 26148 3516
rect 25372 3476 25378 3488
rect 26142 3476 26148 3488
rect 26200 3476 26206 3528
rect 28902 3476 28908 3528
rect 28960 3516 28966 3528
rect 29638 3516 29644 3528
rect 28960 3488 29644 3516
rect 28960 3476 28966 3488
rect 29638 3476 29644 3488
rect 29696 3476 29702 3528
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 33042 3516 33048 3528
rect 32456 3488 33048 3516
rect 32456 3476 32462 3488
rect 33042 3476 33048 3488
rect 33100 3476 33106 3528
rect 33594 3476 33600 3528
rect 33652 3516 33658 3528
rect 34422 3516 34428 3528
rect 33652 3488 34428 3516
rect 33652 3476 33658 3488
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 34790 3476 34796 3528
rect 34848 3516 34854 3528
rect 35802 3516 35808 3528
rect 34848 3488 35808 3516
rect 34848 3476 34854 3488
rect 35802 3476 35808 3488
rect 35860 3476 35866 3528
rect 40678 3476 40684 3528
rect 40736 3516 40742 3528
rect 41322 3516 41328 3528
rect 40736 3488 41328 3516
rect 40736 3476 40742 3488
rect 41322 3476 41328 3488
rect 41380 3476 41386 3528
rect 41874 3476 41880 3528
rect 41932 3516 41938 3528
rect 42702 3516 42708 3528
rect 41932 3488 42708 3516
rect 41932 3476 41938 3488
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 43070 3476 43076 3528
rect 43128 3516 43134 3528
rect 44082 3516 44088 3528
rect 43128 3488 44088 3516
rect 43128 3476 43134 3488
rect 44082 3476 44088 3488
rect 44140 3476 44146 3528
rect 48958 3476 48964 3528
rect 49016 3516 49022 3528
rect 49602 3516 49608 3528
rect 49016 3488 49608 3516
rect 49016 3476 49022 3488
rect 49602 3476 49608 3488
rect 49660 3476 49666 3528
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50890 3516 50896 3528
rect 50212 3488 50896 3516
rect 50212 3476 50218 3488
rect 50890 3476 50896 3488
rect 50948 3476 50954 3528
rect 52546 3476 52552 3528
rect 52604 3516 52610 3528
rect 53650 3516 53656 3528
rect 52604 3488 53656 3516
rect 52604 3476 52610 3488
rect 53650 3476 53656 3488
rect 53708 3476 53714 3528
rect 56042 3476 56048 3528
rect 56100 3516 56106 3528
rect 56502 3516 56508 3528
rect 56100 3488 56508 3516
rect 56100 3476 56106 3488
rect 56502 3476 56508 3488
rect 56560 3476 56566 3528
rect 57238 3476 57244 3528
rect 57296 3516 57302 3528
rect 57790 3516 57796 3528
rect 57296 3488 57796 3516
rect 57296 3476 57302 3488
rect 57790 3476 57796 3488
rect 57848 3476 57854 3528
rect 58434 3476 58440 3528
rect 58492 3516 58498 3528
rect 59170 3516 59176 3528
rect 58492 3488 59176 3516
rect 58492 3476 58498 3488
rect 59170 3476 59176 3488
rect 59228 3476 59234 3528
rect 59630 3476 59636 3528
rect 59688 3516 59694 3528
rect 60642 3516 60648 3528
rect 59688 3488 60648 3516
rect 59688 3476 59694 3488
rect 60642 3476 60648 3488
rect 60700 3476 60706 3528
rect 63218 3476 63224 3528
rect 63276 3516 63282 3528
rect 63276 3488 93854 3516
rect 63276 3476 63282 3488
rect 7650 3408 7656 3460
rect 7708 3448 7714 3460
rect 33778 3448 33784 3460
rect 7708 3420 33784 3448
rect 7708 3408 7714 3420
rect 33778 3408 33784 3420
rect 33836 3408 33842 3460
rect 64322 3408 64328 3460
rect 64380 3448 64386 3460
rect 64782 3448 64788 3460
rect 64380 3420 64788 3448
rect 64380 3408 64386 3420
rect 64782 3408 64788 3420
rect 64840 3408 64846 3460
rect 65518 3408 65524 3460
rect 65576 3448 65582 3460
rect 66162 3448 66168 3460
rect 65576 3420 66168 3448
rect 65576 3408 65582 3420
rect 66162 3408 66168 3420
rect 66220 3408 66226 3460
rect 67910 3408 67916 3460
rect 67968 3448 67974 3460
rect 68922 3448 68928 3460
rect 67968 3420 68928 3448
rect 67968 3408 67974 3420
rect 68922 3408 68928 3420
rect 68980 3408 68986 3460
rect 72602 3408 72608 3460
rect 72660 3448 72666 3460
rect 73062 3448 73068 3460
rect 72660 3420 73068 3448
rect 72660 3408 72666 3420
rect 73062 3408 73068 3420
rect 73120 3408 73126 3460
rect 73798 3408 73804 3460
rect 73856 3448 73862 3460
rect 74442 3448 74448 3460
rect 73856 3420 74448 3448
rect 73856 3408 73862 3420
rect 74442 3408 74448 3420
rect 74500 3408 74506 3460
rect 74994 3408 75000 3460
rect 75052 3448 75058 3460
rect 75822 3448 75828 3460
rect 75052 3420 75828 3448
rect 75052 3408 75058 3420
rect 75822 3408 75828 3420
rect 75880 3408 75886 3460
rect 76190 3408 76196 3460
rect 76248 3448 76254 3460
rect 77202 3448 77208 3460
rect 76248 3420 77208 3448
rect 76248 3408 76254 3420
rect 77202 3408 77208 3420
rect 77260 3408 77266 3460
rect 80882 3408 80888 3460
rect 80940 3448 80946 3460
rect 81342 3448 81348 3460
rect 80940 3420 81348 3448
rect 80940 3408 80946 3420
rect 81342 3408 81348 3420
rect 81400 3408 81406 3460
rect 83274 3408 83280 3460
rect 83332 3448 83338 3460
rect 84102 3448 84108 3460
rect 83332 3420 84108 3448
rect 83332 3408 83338 3420
rect 84102 3408 84108 3420
rect 84160 3408 84166 3460
rect 85666 3408 85672 3460
rect 85724 3448 85730 3460
rect 86770 3448 86776 3460
rect 85724 3420 86776 3448
rect 85724 3408 85730 3420
rect 86770 3408 86776 3420
rect 86828 3408 86834 3460
rect 91554 3408 91560 3460
rect 91612 3448 91618 3460
rect 92382 3448 92388 3460
rect 91612 3420 92388 3448
rect 91612 3408 91618 3420
rect 92382 3408 92388 3420
rect 92440 3408 92446 3460
rect 93826 3448 93854 3488
rect 97442 3476 97448 3528
rect 97500 3516 97506 3528
rect 97902 3516 97908 3528
rect 97500 3488 97908 3516
rect 97500 3476 97506 3488
rect 97902 3476 97908 3488
rect 97960 3476 97966 3528
rect 98638 3476 98644 3528
rect 98696 3516 98702 3528
rect 99282 3516 99288 3528
rect 98696 3488 99288 3516
rect 98696 3476 98702 3488
rect 99282 3476 99288 3488
rect 99340 3476 99346 3528
rect 99834 3476 99840 3528
rect 99892 3516 99898 3528
rect 100662 3516 100668 3528
rect 99892 3488 100668 3516
rect 99892 3476 99898 3488
rect 100662 3476 100668 3488
rect 100720 3476 100726 3528
rect 101030 3476 101036 3528
rect 101088 3516 101094 3528
rect 102042 3516 102048 3528
rect 101088 3488 102048 3516
rect 101088 3476 101094 3488
rect 102042 3476 102048 3488
rect 102100 3476 102106 3528
rect 106918 3476 106924 3528
rect 106976 3516 106982 3528
rect 107562 3516 107568 3528
rect 106976 3488 107568 3516
rect 106976 3476 106982 3488
rect 107562 3476 107568 3488
rect 107620 3476 107626 3528
rect 108114 3476 108120 3528
rect 108172 3516 108178 3528
rect 108942 3516 108948 3528
rect 108172 3488 108948 3516
rect 108172 3476 108178 3488
rect 108942 3476 108948 3488
rect 109000 3476 109006 3528
rect 109310 3476 109316 3528
rect 109368 3516 109374 3528
rect 110322 3516 110328 3528
rect 109368 3488 110328 3516
rect 109368 3476 109374 3488
rect 110322 3476 110328 3488
rect 110380 3476 110386 3528
rect 110506 3476 110512 3528
rect 110564 3516 110570 3528
rect 111702 3516 111708 3528
rect 110564 3488 111708 3516
rect 110564 3476 110570 3488
rect 111702 3476 111708 3488
rect 111760 3476 111766 3528
rect 115198 3476 115204 3528
rect 115256 3516 115262 3528
rect 115842 3516 115848 3528
rect 115256 3488 115848 3516
rect 115256 3476 115262 3488
rect 115842 3476 115848 3488
rect 115900 3476 115906 3528
rect 116394 3476 116400 3528
rect 116452 3516 116458 3528
rect 117222 3516 117228 3528
rect 116452 3488 117228 3516
rect 116452 3476 116458 3488
rect 117222 3476 117228 3488
rect 117280 3476 117286 3528
rect 117590 3476 117596 3528
rect 117648 3516 117654 3528
rect 118602 3516 118608 3528
rect 117648 3488 118608 3516
rect 117648 3476 117654 3488
rect 118602 3476 118608 3488
rect 118660 3476 118666 3528
rect 118786 3476 118792 3528
rect 118844 3516 118850 3528
rect 119798 3516 119804 3528
rect 118844 3488 119804 3516
rect 118844 3476 118850 3488
rect 119798 3476 119804 3488
rect 119856 3476 119862 3528
rect 122282 3476 122288 3528
rect 122340 3516 122346 3528
rect 122742 3516 122748 3528
rect 122340 3488 122748 3516
rect 122340 3476 122346 3488
rect 122742 3476 122748 3488
rect 122800 3476 122806 3528
rect 123478 3476 123484 3528
rect 123536 3516 123542 3528
rect 124122 3516 124128 3528
rect 123536 3488 124128 3516
rect 123536 3476 123542 3488
rect 124122 3476 124128 3488
rect 124180 3476 124186 3528
rect 124674 3476 124680 3528
rect 124732 3516 124738 3528
rect 125502 3516 125508 3528
rect 124732 3488 125508 3516
rect 124732 3476 124738 3488
rect 125502 3476 125508 3488
rect 125560 3476 125566 3528
rect 129366 3476 129372 3528
rect 129424 3516 129430 3528
rect 130378 3516 130384 3528
rect 129424 3488 130384 3516
rect 129424 3476 129430 3488
rect 130378 3476 130384 3488
rect 130436 3476 130442 3528
rect 231118 3476 231124 3528
rect 231176 3516 231182 3528
rect 247586 3516 247592 3528
rect 231176 3488 247592 3516
rect 231176 3476 231182 3488
rect 247586 3476 247592 3488
rect 247644 3476 247650 3528
rect 250438 3476 250444 3528
rect 250496 3516 250502 3528
rect 271230 3516 271236 3528
rect 250496 3488 271236 3516
rect 250496 3476 250502 3488
rect 271230 3476 271236 3488
rect 271288 3476 271294 3528
rect 271414 3476 271420 3528
rect 271472 3516 271478 3528
rect 272426 3516 272432 3528
rect 271472 3488 272432 3516
rect 271472 3476 271478 3488
rect 272426 3476 272432 3488
rect 272484 3476 272490 3528
rect 307754 3476 307760 3528
rect 307812 3516 307818 3528
rect 309042 3516 309048 3528
rect 307812 3488 309048 3516
rect 307812 3476 307818 3488
rect 309042 3476 309048 3488
rect 309100 3476 309106 3528
rect 322198 3476 322204 3528
rect 322256 3516 322262 3528
rect 323302 3516 323308 3528
rect 322256 3488 323308 3516
rect 322256 3476 322262 3488
rect 323302 3476 323308 3488
rect 323360 3476 323366 3528
rect 324314 3476 324320 3528
rect 324372 3516 324378 3528
rect 325602 3516 325608 3528
rect 324372 3488 325608 3516
rect 324372 3476 324378 3488
rect 325602 3476 325608 3488
rect 325660 3476 325666 3528
rect 332594 3476 332600 3528
rect 332652 3516 332658 3528
rect 333882 3516 333888 3528
rect 332652 3488 333888 3516
rect 332652 3476 332658 3488
rect 333882 3476 333888 3488
rect 333940 3476 333946 3528
rect 337470 3476 337476 3528
rect 337528 3516 337534 3528
rect 338114 3516 338120 3528
rect 337528 3488 338120 3516
rect 337528 3476 337534 3488
rect 338114 3476 338120 3488
rect 338172 3476 338178 3528
rect 350442 3476 350448 3528
rect 350500 3516 350506 3528
rect 353294 3516 353300 3528
rect 350500 3488 353300 3516
rect 350500 3476 350506 3488
rect 353294 3476 353300 3488
rect 353352 3476 353358 3528
rect 582190 3476 582196 3528
rect 582248 3516 582254 3528
rect 583478 3516 583484 3528
rect 582248 3488 583484 3516
rect 582248 3476 582254 3488
rect 583478 3476 583484 3488
rect 583536 3476 583542 3528
rect 105538 3448 105544 3460
rect 93826 3420 105544 3448
rect 105538 3408 105544 3420
rect 105596 3408 105602 3460
rect 105722 3408 105728 3460
rect 105780 3448 105786 3460
rect 229738 3448 229744 3460
rect 105780 3420 229744 3448
rect 105780 3408 105786 3420
rect 229738 3408 229744 3420
rect 229796 3408 229802 3460
rect 242158 3408 242164 3460
rect 242216 3448 242222 3460
rect 293678 3448 293684 3460
rect 242216 3420 293684 3448
rect 242216 3408 242222 3420
rect 293678 3408 293684 3420
rect 293736 3408 293742 3460
rect 295978 3408 295984 3460
rect 296036 3448 296042 3460
rect 304350 3448 304356 3460
rect 296036 3420 304356 3448
rect 296036 3408 296042 3420
rect 304350 3408 304356 3420
rect 304408 3408 304414 3460
rect 306742 3408 306748 3460
rect 306800 3448 306806 3460
rect 317414 3448 317420 3460
rect 306800 3420 317420 3448
rect 306800 3408 306806 3420
rect 317414 3408 317420 3420
rect 317472 3408 317478 3460
rect 77386 3340 77392 3392
rect 77444 3380 77450 3392
rect 88978 3380 88984 3392
rect 77444 3352 88984 3380
rect 77444 3340 77450 3352
rect 88978 3340 88984 3352
rect 89036 3340 89042 3392
rect 298738 3272 298744 3324
rect 298796 3312 298802 3324
rect 301958 3312 301964 3324
rect 298796 3284 301964 3312
rect 298796 3272 298802 3284
rect 301958 3272 301964 3284
rect 302016 3272 302022 3324
rect 316218 3272 316224 3324
rect 316276 3312 316282 3324
rect 320174 3312 320180 3324
rect 316276 3284 320180 3312
rect 316276 3272 316282 3284
rect 320174 3272 320180 3284
rect 320232 3272 320238 3324
rect 346946 3272 346952 3324
rect 347004 3312 347010 3324
rect 351914 3312 351920 3324
rect 347004 3284 351920 3312
rect 347004 3272 347010 3284
rect 351914 3272 351920 3284
rect 351972 3272 351978 3324
rect 17034 3204 17040 3256
rect 17092 3244 17098 3256
rect 17862 3244 17868 3256
rect 17092 3216 17868 3244
rect 17092 3204 17098 3216
rect 17862 3204 17868 3216
rect 17920 3204 17926 3256
rect 280798 3068 280804 3120
rect 280856 3108 280862 3120
rect 283098 3108 283104 3120
rect 280856 3080 283104 3108
rect 280856 3068 280862 3080
rect 283098 3068 283104 3080
rect 283156 3068 283162 3120
rect 347038 3068 347044 3120
rect 347096 3108 347102 3120
rect 349246 3108 349252 3120
rect 347096 3080 349252 3108
rect 347096 3068 347102 3080
rect 349246 3068 349252 3080
rect 349304 3068 349310 3120
rect 90358 3000 90364 3052
rect 90416 3040 90422 3052
rect 91002 3040 91008 3052
rect 90416 3012 91008 3040
rect 90416 3000 90422 3012
rect 91002 3000 91008 3012
rect 91060 3000 91066 3052
rect 93946 3000 93952 3052
rect 94004 3040 94010 3052
rect 95050 3040 95056 3052
rect 94004 3012 95056 3040
rect 94004 3000 94010 3012
rect 95050 3000 95056 3012
rect 95108 3000 95114 3052
rect 580994 3000 581000 3052
rect 581052 3040 581058 3052
rect 583570 3040 583576 3052
rect 581052 3012 583576 3040
rect 581052 3000 581058 3012
rect 583570 3000 583576 3012
rect 583628 3000 583634 3052
rect 332686 2932 332692 2984
rect 332744 2972 332750 2984
rect 335354 2972 335360 2984
rect 332744 2944 335360 2972
rect 332744 2932 332750 2944
rect 335354 2932 335360 2944
rect 335412 2932 335418 2984
rect 84470 2116 84476 2168
rect 84528 2156 84534 2168
rect 196710 2156 196716 2168
rect 84528 2128 196716 2156
rect 84528 2116 84534 2128
rect 196710 2116 196716 2128
rect 196768 2116 196774 2168
rect 238018 2116 238024 2168
rect 238076 2156 238082 2168
rect 305546 2156 305552 2168
rect 238076 2128 305552 2156
rect 238076 2116 238082 2128
rect 305546 2116 305552 2128
rect 305604 2116 305610 2168
rect 26510 2048 26516 2100
rect 26568 2088 26574 2100
rect 265618 2088 265624 2100
rect 26568 2060 265624 2088
rect 26568 2048 26574 2060
rect 265618 2048 265624 2060
rect 265676 2048 265682 2100
<< via1 >>
rect 75828 703604 75880 703656
rect 202604 703604 202656 703656
rect 86868 703536 86920 703588
rect 234988 703536 235040 703588
rect 67640 703468 67692 703520
rect 267464 703468 267516 703520
rect 93768 703400 93820 703452
rect 300124 703400 300176 703452
rect 59268 703332 59320 703384
rect 283840 703332 283892 703384
rect 73068 703264 73120 703316
rect 332508 703264 332560 703316
rect 130384 703196 130436 703248
rect 413652 703196 413704 703248
rect 62028 703128 62080 703180
rect 348792 703128 348844 703180
rect 98736 703060 98788 703112
rect 397460 703060 397512 703112
rect 124864 702992 124916 703044
rect 429844 702992 429896 703044
rect 57888 702924 57940 702976
rect 364984 702924 365036 702976
rect 126244 702856 126296 702908
rect 462320 702856 462372 702908
rect 71044 702788 71096 702840
rect 494796 702788 494848 702840
rect 97908 702720 97960 702772
rect 478512 702720 478564 702772
rect 129004 702652 129056 702704
rect 543464 702652 543516 702704
rect 8116 702584 8168 702636
rect 89812 702584 89864 702636
rect 94504 702584 94556 702636
rect 527180 702584 527232 702636
rect 55128 702516 55180 702568
rect 580264 702516 580316 702568
rect 66168 702448 66220 702500
rect 559656 702448 559708 702500
rect 83464 700272 83516 700324
rect 89168 700272 89220 700324
rect 88984 700204 89036 700256
rect 105452 700272 105504 700324
rect 133144 700272 133196 700324
rect 218980 700272 219032 700324
rect 24308 698912 24360 698964
rect 79324 698912 79376 698964
rect 3516 670692 3568 670744
rect 22744 670692 22796 670744
rect 2780 656956 2832 657008
rect 4804 656956 4856 657008
rect 3516 632068 3568 632120
rect 25504 632068 25556 632120
rect 3516 618264 3568 618316
rect 36544 618264 36596 618316
rect 3516 605820 3568 605872
rect 87604 605820 87656 605872
rect 79324 600244 79376 600296
rect 79968 600244 80020 600296
rect 67456 599564 67508 599616
rect 88984 599564 89036 599616
rect 79968 598952 80020 599004
rect 114560 598952 114612 599004
rect 40040 598204 40092 598256
rect 88892 598204 88944 598256
rect 67548 596776 67600 596828
rect 169760 596776 169812 596828
rect 88984 595416 89036 595468
rect 108304 595416 108356 595468
rect 582748 595416 582800 595468
rect 79784 594804 79836 594856
rect 105544 594804 105596 594856
rect 87604 594396 87656 594448
rect 91192 594396 91244 594448
rect 86224 593376 86276 593428
rect 128544 593376 128596 593428
rect 582748 593376 582800 593428
rect 4804 592628 4856 592680
rect 69020 592628 69072 592680
rect 75644 592084 75696 592136
rect 96620 592084 96672 592136
rect 77944 592016 77996 592068
rect 102140 592016 102192 592068
rect 70308 590724 70360 590776
rect 75184 590724 75236 590776
rect 84108 590724 84160 590776
rect 95884 590724 95936 590776
rect 78404 590656 78456 590708
rect 100760 590656 100812 590708
rect 75184 589908 75236 589960
rect 89720 589908 89772 589960
rect 72884 589364 72936 589416
rect 93860 589364 93912 589416
rect 4804 589296 4856 589348
rect 74862 589296 74914 589348
rect 75644 589296 75696 589348
rect 82636 589228 82688 589280
rect 86960 589228 87012 589280
rect 69480 588616 69532 588668
rect 85304 588548 85356 588600
rect 87052 588548 87104 588600
rect 113180 588548 113232 588600
rect 83740 588412 83792 588464
rect 52368 587868 52420 587920
rect 66812 587868 66864 587920
rect 88892 588276 88944 588328
rect 100760 588140 100812 588192
rect 103520 588140 103572 588192
rect 92480 587800 92532 587852
rect 59176 586508 59228 586560
rect 66260 586508 66312 586560
rect 48228 585148 48280 585200
rect 67732 585148 67784 585200
rect 91928 584400 91980 584452
rect 93768 584400 93820 584452
rect 124220 584400 124272 584452
rect 91836 583652 91888 583704
rect 93768 583652 93820 583704
rect 94504 583652 94556 583704
rect 50896 582360 50948 582412
rect 66812 582360 66864 582412
rect 91100 581000 91152 581052
rect 104164 581000 104216 581052
rect 2780 580456 2832 580508
rect 4804 580456 4856 580508
rect 64788 579640 64840 579692
rect 66812 579640 66864 579692
rect 91100 578212 91152 578264
rect 121644 578212 121696 578264
rect 143448 577464 143500 577516
rect 582472 577464 582524 577516
rect 91100 576852 91152 576904
rect 142160 576852 142212 576904
rect 143448 576852 143500 576904
rect 25504 576104 25556 576156
rect 47860 576104 47912 576156
rect 91192 576104 91244 576156
rect 105636 576104 105688 576156
rect 47860 575492 47912 575544
rect 48136 575492 48188 575544
rect 66904 575492 66956 575544
rect 55036 574744 55088 574796
rect 67456 574744 67508 574796
rect 91100 574744 91152 574796
rect 95148 574744 95200 574796
rect 98736 574744 98788 574796
rect 91100 572704 91152 572756
rect 120632 572704 120684 572756
rect 91192 571412 91244 571464
rect 108396 571412 108448 571464
rect 63316 571344 63368 571396
rect 66444 571344 66496 571396
rect 91100 571344 91152 571396
rect 129740 571344 129792 571396
rect 91100 569916 91152 569968
rect 116584 569916 116636 569968
rect 60556 568556 60608 568608
rect 66904 568556 66956 568608
rect 57796 567196 57848 567248
rect 66904 567196 66956 567248
rect 88892 567196 88944 567248
rect 133880 567196 133932 567248
rect 53748 566448 53800 566500
rect 67548 566448 67600 566500
rect 3240 565836 3292 565888
rect 43444 565836 43496 565888
rect 91100 565836 91152 565888
rect 126980 565836 127032 565888
rect 95884 565088 95936 565140
rect 111800 565088 111852 565140
rect 51724 564340 51776 564392
rect 55128 564340 55180 564392
rect 66812 564340 66864 564392
rect 91100 563048 91152 563100
rect 133236 563048 133288 563100
rect 92204 562300 92256 562352
rect 120724 562300 120776 562352
rect 35808 561688 35860 561740
rect 66812 561688 66864 561740
rect 39948 560260 40000 560312
rect 66536 560260 66588 560312
rect 56508 558900 56560 558952
rect 66536 558900 66588 558952
rect 95148 558152 95200 558204
rect 123208 558152 123260 558204
rect 50988 557540 51040 557592
rect 67640 557540 67692 557592
rect 91192 557540 91244 557592
rect 125600 557540 125652 557592
rect 91192 556180 91244 556232
rect 121460 556180 121512 556232
rect 58900 554752 58952 554804
rect 66628 554752 66680 554804
rect 91192 554752 91244 554804
rect 100668 554752 100720 554804
rect 582472 554752 582524 554804
rect 3516 553800 3568 553852
rect 7564 553800 7616 553852
rect 59268 553460 59320 553512
rect 64144 553460 64196 553512
rect 66536 553460 66588 553512
rect 107016 553052 107068 553104
rect 109040 553052 109092 553104
rect 91192 552304 91244 552356
rect 95240 552304 95292 552356
rect 91192 552032 91244 552084
rect 106924 552032 106976 552084
rect 60648 549244 60700 549296
rect 66444 549244 66496 549296
rect 91192 549244 91244 549296
rect 98736 549244 98788 549296
rect 91836 548496 91888 548548
rect 121552 548496 121604 548548
rect 63408 547884 63460 547936
rect 66536 547884 66588 547936
rect 62028 547748 62080 547800
rect 66628 547748 66680 547800
rect 3424 547136 3476 547188
rect 41236 547136 41288 547188
rect 41328 547136 41380 547188
rect 62028 547136 62080 547188
rect 89996 546388 90048 546440
rect 91008 546388 91060 546440
rect 126244 546388 126296 546440
rect 57520 545708 57572 545760
rect 66168 545708 66220 545760
rect 91192 544348 91244 544400
rect 95148 544348 95200 544400
rect 129004 544348 129056 544400
rect 57888 543736 57940 543788
rect 62028 543736 62080 543788
rect 66812 543736 66864 543788
rect 41236 542376 41288 542428
rect 44088 542376 44140 542428
rect 66812 542376 66864 542428
rect 91192 542376 91244 542428
rect 104256 542376 104308 542428
rect 22744 541628 22796 541680
rect 67088 541628 67140 541680
rect 91192 541628 91244 541680
rect 136640 541628 136692 541680
rect 67548 540880 67600 540932
rect 68652 540880 68704 540932
rect 582656 540880 582708 540932
rect 65984 539656 66036 539708
rect 91192 539656 91244 539708
rect 93124 539656 93176 539708
rect 55128 539588 55180 539640
rect 67548 539588 67600 539640
rect 69848 539588 69900 539640
rect 89536 539520 89588 539572
rect 89904 539520 89956 539572
rect 67088 539452 67140 539504
rect 67548 539452 67600 539504
rect 67824 538908 67876 538960
rect 74724 538908 74776 538960
rect 3424 538296 3476 538348
rect 89536 538296 89588 538348
rect 80336 538228 80388 538280
rect 80796 538228 80848 538280
rect 582564 538228 582616 538280
rect 7564 538160 7616 538212
rect 70676 538160 70728 538212
rect 86868 538160 86920 538212
rect 133144 538160 133196 538212
rect 72424 537480 72476 537532
rect 579804 537480 579856 537532
rect 43444 536732 43496 536784
rect 69664 536732 69716 536784
rect 82728 536732 82780 536784
rect 130384 536732 130436 536784
rect 85488 536188 85540 536240
rect 86224 536188 86276 536240
rect 36544 536052 36596 536104
rect 49608 536052 49660 536104
rect 73160 536052 73212 536104
rect 73160 535440 73212 535492
rect 73988 535440 74040 535492
rect 88616 535440 88668 535492
rect 89628 535440 89680 535492
rect 8208 534692 8260 534744
rect 91284 534692 91336 534744
rect 56508 534012 56560 534064
rect 580264 534012 580316 534064
rect 67640 533400 67692 533452
rect 68468 533400 68520 533452
rect 78680 533400 78732 533452
rect 79508 533400 79560 533452
rect 4804 533332 4856 533384
rect 91376 533332 91428 533384
rect 64788 531972 64840 532024
rect 77944 531972 77996 532024
rect 23388 530544 23440 530596
rect 91100 530544 91152 530596
rect 66168 529184 66220 529236
rect 76472 529184 76524 529236
rect 3424 514768 3476 514820
rect 11704 514768 11756 514820
rect 39948 511232 40000 511284
rect 580172 511232 580224 511284
rect 2780 501848 2832 501900
rect 4804 501848 4856 501900
rect 67732 476008 67784 476060
rect 76564 476008 76616 476060
rect 63316 475464 63368 475516
rect 67824 475464 67876 475516
rect 3332 475328 3384 475380
rect 8208 475328 8260 475380
rect 17224 475328 17276 475380
rect 57612 471248 57664 471300
rect 78680 471248 78732 471300
rect 59084 468460 59136 468512
rect 75920 468460 75972 468512
rect 89536 465740 89588 465792
rect 125692 465740 125744 465792
rect 53656 465672 53708 465724
rect 95884 465672 95936 465724
rect 66076 464312 66128 464364
rect 78680 464312 78732 464364
rect 59176 462952 59228 463004
rect 85580 462952 85632 463004
rect 2780 462544 2832 462596
rect 4804 462544 4856 462596
rect 69020 462272 69072 462324
rect 69848 462272 69900 462324
rect 52276 461592 52328 461644
rect 73160 461592 73212 461644
rect 69020 460912 69072 460964
rect 178040 460912 178092 460964
rect 48228 460164 48280 460216
rect 82820 460164 82872 460216
rect 112444 458872 112496 458924
rect 117320 458872 117372 458924
rect 106280 458804 106332 458856
rect 114560 458804 114612 458856
rect 152464 458804 152516 458856
rect 52368 458192 52420 458244
rect 53564 458192 53616 458244
rect 86960 458192 87012 458244
rect 63316 457444 63368 457496
rect 80060 457444 80112 457496
rect 61844 456016 61896 456068
rect 70492 456016 70544 456068
rect 77392 455336 77444 455388
rect 77944 455336 77996 455388
rect 48136 454656 48188 454708
rect 73160 454656 73212 454708
rect 77392 454112 77444 454164
rect 128452 454112 128504 454164
rect 73160 454044 73212 454096
rect 144184 454044 144236 454096
rect 22744 453976 22796 454028
rect 23388 453976 23440 454028
rect 61752 453296 61804 453348
rect 78772 453296 78824 453348
rect 82820 452684 82872 452736
rect 83464 452684 83516 452736
rect 161480 452684 161532 452736
rect 22744 452616 22796 452668
rect 124956 452616 125008 452668
rect 61936 451868 61988 451920
rect 91560 451868 91612 451920
rect 50804 451256 50856 451308
rect 74724 451256 74776 451308
rect 98644 451256 98696 451308
rect 179420 451256 179472 451308
rect 4804 451188 4856 451240
rect 103520 451188 103572 451240
rect 104624 451188 104676 451240
rect 173808 451188 173860 451240
rect 582472 451188 582524 451240
rect 55036 450508 55088 450560
rect 71780 450508 71832 450560
rect 104072 449964 104124 450016
rect 104624 449964 104676 450016
rect 167000 449964 167052 450016
rect 50896 449828 50948 449880
rect 80888 449828 80940 449880
rect 172520 449896 172572 449948
rect 173808 449896 173860 449948
rect 64696 449148 64748 449200
rect 74632 449148 74684 449200
rect 116584 449148 116636 449200
rect 128360 449148 128412 449200
rect 3148 448536 3200 448588
rect 40684 448536 40736 448588
rect 108304 448536 108356 448588
rect 130384 448536 130436 448588
rect 11704 448468 11756 448520
rect 111800 448468 111852 448520
rect 105636 447788 105688 447840
rect 122932 447788 122984 447840
rect 68376 447108 68428 447160
rect 88800 447108 88852 447160
rect 60464 446360 60516 446412
rect 77300 446360 77352 446412
rect 111800 445816 111852 445868
rect 112996 445816 113048 445868
rect 142804 445816 142856 445868
rect 76564 445748 76616 445800
rect 124864 445748 124916 445800
rect 59176 444456 59228 444508
rect 92480 444456 92532 444508
rect 93078 444456 93130 444508
rect 101404 444456 101456 444508
rect 126244 444456 126296 444508
rect 4804 444388 4856 444440
rect 118700 444388 118752 444440
rect 67364 442892 67416 442944
rect 67732 442892 67784 442944
rect 60372 442212 60424 442264
rect 68376 442212 68428 442264
rect 124128 439492 124180 439544
rect 125692 439492 125744 439544
rect 157340 439492 157392 439544
rect 60556 439016 60608 439068
rect 66996 439016 67048 439068
rect 67364 439016 67416 439068
rect 57796 438132 57848 438184
rect 66076 438132 66128 438184
rect 66536 438132 66588 438184
rect 123668 438132 123720 438184
rect 124220 438132 124272 438184
rect 157984 438132 158036 438184
rect 52460 436024 52512 436076
rect 53748 436024 53800 436076
rect 66812 436024 66864 436076
rect 39856 435344 39908 435396
rect 52460 435344 52512 435396
rect 52184 433304 52236 433356
rect 65524 433304 65576 433356
rect 66444 433236 66496 433288
rect 123852 432556 123904 432608
rect 171140 432556 171192 432608
rect 582380 432556 582432 432608
rect 48136 431944 48188 431996
rect 51724 431876 51776 431928
rect 66812 431876 66864 431928
rect 34520 429088 34572 429140
rect 35808 429088 35860 429140
rect 66812 429088 66864 429140
rect 15844 428408 15896 428460
rect 34520 428408 34572 428460
rect 39948 425688 40000 425740
rect 58992 425688 59044 425740
rect 58992 425076 59044 425128
rect 66812 425076 66864 425128
rect 56508 424328 56560 424380
rect 63224 424328 63276 424380
rect 66812 424328 66864 424380
rect 3424 423580 3476 423632
rect 22744 423580 22796 423632
rect 50988 421540 51040 421592
rect 64788 421540 64840 421592
rect 66812 421540 66864 421592
rect 123208 421540 123260 421592
rect 134524 421540 134576 421592
rect 56508 419500 56560 419552
rect 66904 419500 66956 419552
rect 58900 418072 58952 418124
rect 65524 418072 65576 418124
rect 66444 418072 66496 418124
rect 124128 415148 124180 415200
rect 129740 415148 129792 415200
rect 57796 414672 57848 414724
rect 64144 414672 64196 414724
rect 66812 414672 66864 414724
rect 129740 414672 129792 414724
rect 131120 414672 131172 414724
rect 123024 412564 123076 412616
rect 128360 412564 128412 412616
rect 123024 411272 123076 411324
rect 123484 411272 123536 411324
rect 121184 409844 121236 409896
rect 135904 409844 135956 409896
rect 60648 408416 60700 408468
rect 68376 408416 68428 408468
rect 124128 407736 124180 407788
rect 133880 407736 133932 407788
rect 134616 407736 134668 407788
rect 63408 406580 63460 406632
rect 64604 406580 64656 406632
rect 64604 406104 64656 406156
rect 66260 406104 66312 406156
rect 124128 406104 124180 406156
rect 126888 406104 126940 406156
rect 41328 404948 41380 405000
rect 57704 404948 57756 405000
rect 57704 403588 57756 403640
rect 66260 403588 66312 403640
rect 163504 403588 163556 403640
rect 582380 403588 582432 403640
rect 124036 402976 124088 403028
rect 163504 402976 163556 403028
rect 50896 401548 50948 401600
rect 57520 401548 57572 401600
rect 66260 401548 66312 401600
rect 124128 401548 124180 401600
rect 133236 401548 133288 401600
rect 133788 401548 133840 401600
rect 124956 400188 125008 400240
rect 169760 400188 169812 400240
rect 123668 400120 123720 400172
rect 2780 398692 2832 398744
rect 4804 398692 4856 398744
rect 43996 398080 44048 398132
rect 62028 398080 62080 398132
rect 66444 398080 66496 398132
rect 44088 396720 44140 396772
rect 66996 396720 67048 396772
rect 67272 396720 67324 396772
rect 121552 396040 121604 396092
rect 171232 396040 171284 396092
rect 123668 395972 123720 396024
rect 125600 395972 125652 396024
rect 55128 393252 55180 393304
rect 61936 393252 61988 393304
rect 66812 393252 66864 393304
rect 59084 391212 59136 391264
rect 81440 390940 81492 390992
rect 82084 390940 82136 390992
rect 115848 390532 115900 390584
rect 120816 390532 120868 390584
rect 3424 389784 3476 389836
rect 85488 389784 85540 389836
rect 57612 389172 57664 389224
rect 86960 389172 87012 389224
rect 117780 389172 117832 389224
rect 165620 389172 165672 389224
rect 49608 389104 49660 389156
rect 76656 389104 76708 389156
rect 104072 389104 104124 389156
rect 136640 389104 136692 389156
rect 61844 389036 61896 389088
rect 67640 389036 67692 389088
rect 68468 389036 68520 389088
rect 119436 389036 119488 389088
rect 120172 389036 120224 389088
rect 73160 388968 73212 389020
rect 73344 388968 73396 389020
rect 93400 388424 93452 388476
rect 112444 388424 112496 388476
rect 93676 388016 93728 388068
rect 94228 388016 94280 388068
rect 79968 387812 80020 387864
rect 80612 387812 80664 387864
rect 64696 387744 64748 387796
rect 79324 387744 79376 387796
rect 111708 387064 111760 387116
rect 120632 387064 120684 387116
rect 52276 386316 52328 386368
rect 77944 386316 77996 386368
rect 61752 386248 61804 386300
rect 85580 386248 85632 386300
rect 63316 384956 63368 385008
rect 88984 384956 89036 385008
rect 52276 384276 52328 384328
rect 122932 384276 122984 384328
rect 60464 383596 60516 383648
rect 82820 383596 82872 383648
rect 108764 382916 108816 382968
rect 160100 382916 160152 382968
rect 4804 381488 4856 381540
rect 123484 381488 123536 381540
rect 110420 380196 110472 380248
rect 158720 380196 158772 380248
rect 67732 380128 67784 380180
rect 124956 380128 125008 380180
rect 53564 378768 53616 378820
rect 75920 378768 75972 378820
rect 104900 376728 104952 376780
rect 228364 376728 228416 376780
rect 52184 375980 52236 376032
rect 163596 375980 163648 376032
rect 39856 375368 39908 375420
rect 188344 375368 188396 375420
rect 118700 374688 118752 374740
rect 165712 374688 165764 374740
rect 70308 374620 70360 374672
rect 164332 374620 164384 374672
rect 71688 374212 71740 374264
rect 73160 374212 73212 374264
rect 3424 373260 3476 373312
rect 118608 373260 118660 373312
rect 67548 372648 67600 372700
rect 201500 372648 201552 372700
rect 142068 372580 142120 372632
rect 331220 372580 331272 372632
rect 129740 371288 129792 371340
rect 232504 371288 232556 371340
rect 81440 371220 81492 371272
rect 240508 371220 240560 371272
rect 3148 370472 3200 370524
rect 7564 370472 7616 370524
rect 11704 370472 11756 370524
rect 60372 370472 60424 370524
rect 78680 370472 78732 370524
rect 79968 370472 80020 370524
rect 161572 370472 161624 370524
rect 73160 369860 73212 369912
rect 188436 369860 188488 369912
rect 107476 369180 107528 369232
rect 151084 369180 151136 369232
rect 62028 369112 62080 369164
rect 111800 369112 111852 369164
rect 125600 368908 125652 368960
rect 126244 368908 126296 368960
rect 126244 368500 126296 368552
rect 231124 368500 231176 368552
rect 99288 367752 99340 367804
rect 170404 367752 170456 367804
rect 132500 367072 132552 367124
rect 251272 367072 251324 367124
rect 137284 367004 137336 367056
rect 137836 367004 137888 367056
rect 137836 365780 137888 365832
rect 162124 365780 162176 365832
rect 78680 365712 78732 365764
rect 243176 365712 243228 365764
rect 93124 365644 93176 365696
rect 93676 365644 93728 365696
rect 128360 365644 128412 365696
rect 129004 365644 129056 365696
rect 79324 364964 79376 365016
rect 122932 364964 122984 365016
rect 128360 364964 128412 365016
rect 212908 364964 212960 365016
rect 98736 362992 98788 363044
rect 181536 362992 181588 363044
rect 80060 362924 80112 362976
rect 81348 362924 81400 362976
rect 251180 362924 251232 362976
rect 78772 361564 78824 361616
rect 79968 361564 80020 361616
rect 198004 361632 198056 361684
rect 117228 361564 117280 361616
rect 241520 361564 241572 361616
rect 115204 360204 115256 360256
rect 115848 360204 115900 360256
rect 214564 360204 214616 360256
rect 71596 359456 71648 359508
rect 123116 359456 123168 359508
rect 122932 358844 122984 358896
rect 186964 358844 187016 358896
rect 124956 358776 125008 358828
rect 224224 358776 224276 358828
rect 105636 358028 105688 358080
rect 155316 358028 155368 358080
rect 155868 357484 155920 357536
rect 176016 357484 176068 357536
rect 140688 357416 140740 357468
rect 207664 357416 207716 357468
rect 70400 356736 70452 356788
rect 71688 356736 71740 356788
rect 102140 356124 102192 356176
rect 193864 356124 193916 356176
rect 71688 356056 71740 356108
rect 238024 356056 238076 356108
rect 90364 354764 90416 354816
rect 191104 354764 191156 354816
rect 128360 354696 128412 354748
rect 230480 354696 230532 354748
rect 134616 353336 134668 353388
rect 138020 353336 138072 353388
rect 169024 353336 169076 353388
rect 65616 353268 65668 353320
rect 67640 353268 67692 353320
rect 69848 353268 69900 353320
rect 184296 353268 184348 353320
rect 202144 352724 202196 352776
rect 202788 352724 202840 352776
rect 97816 352520 97868 352572
rect 154672 352520 154724 352572
rect 202788 352520 202840 352572
rect 580172 352520 580224 352572
rect 144184 351908 144236 351960
rect 146300 351908 146352 351960
rect 195428 351908 195480 351960
rect 104808 351228 104860 351280
rect 120724 351228 120776 351280
rect 110328 351160 110380 351212
rect 155224 351160 155276 351212
rect 85488 350548 85540 350600
rect 90364 350548 90416 350600
rect 123484 350548 123536 350600
rect 177396 350548 177448 350600
rect 63316 349800 63368 349852
rect 71596 349800 71648 349852
rect 222844 349800 222896 349852
rect 118700 349120 118752 349172
rect 119344 349120 119396 349172
rect 249800 349120 249852 349172
rect 92296 349052 92348 349104
rect 118792 349052 118844 349104
rect 119436 349052 119488 349104
rect 122748 348440 122800 348492
rect 130476 348440 130528 348492
rect 96528 348372 96580 348424
rect 128452 348372 128504 348424
rect 142804 348372 142856 348424
rect 156052 348372 156104 348424
rect 133144 347760 133196 347812
rect 222936 347760 222988 347812
rect 78588 347012 78640 347064
rect 93124 347012 93176 347064
rect 96436 347012 96488 347064
rect 116584 347012 116636 347064
rect 135168 346468 135220 346520
rect 198096 346468 198148 346520
rect 66076 346400 66128 346452
rect 196716 346400 196768 346452
rect 3148 346332 3200 346384
rect 33784 346332 33836 346384
rect 92388 345652 92440 345704
rect 121460 345652 121512 345704
rect 143540 345108 143592 345160
rect 183008 345108 183060 345160
rect 67272 345040 67324 345092
rect 224316 345040 224368 345092
rect 49608 344292 49660 344344
rect 82820 344292 82872 344344
rect 99380 343680 99432 343732
rect 100116 343680 100168 343732
rect 167644 343680 167696 343732
rect 97264 343612 97316 343664
rect 246304 343612 246356 343664
rect 134248 342320 134300 342372
rect 173348 342320 173400 342372
rect 67640 342252 67692 342304
rect 167736 342252 167788 342304
rect 61752 340960 61804 341012
rect 141424 341028 141476 341080
rect 140780 340960 140832 341012
rect 225604 340960 225656 341012
rect 60556 340892 60608 340944
rect 145380 340892 145432 340944
rect 146208 340892 146260 340944
rect 357440 340892 357492 340944
rect 74356 340144 74408 340196
rect 93216 340144 93268 340196
rect 63224 339532 63276 339584
rect 159456 339532 159508 339584
rect 115940 339464 115992 339516
rect 244280 339464 244332 339516
rect 137008 338172 137060 338224
rect 164884 338172 164936 338224
rect 71780 338104 71832 338156
rect 216036 338104 216088 338156
rect 66168 337424 66220 337476
rect 74540 337424 74592 337476
rect 54852 337356 54904 337408
rect 86960 337356 87012 337408
rect 120080 337356 120132 337408
rect 140780 337356 140832 337408
rect 92848 336812 92900 336864
rect 178776 336812 178828 336864
rect 146944 336744 146996 336796
rect 252652 336744 252704 336796
rect 113180 335996 113232 336048
rect 139400 335996 139452 336048
rect 140780 335996 140832 336048
rect 146944 335996 146996 336048
rect 61844 335384 61896 335436
rect 203524 335384 203576 335436
rect 149152 335316 149204 335368
rect 335360 335316 335412 335368
rect 60464 334568 60516 334620
rect 113180 334568 113232 334620
rect 115664 334024 115716 334076
rect 173256 334024 173308 334076
rect 59268 333956 59320 334008
rect 89904 333956 89956 334008
rect 104256 333956 104308 334008
rect 220176 333956 220228 334008
rect 91560 333072 91612 333124
rect 94504 333072 94556 333124
rect 113640 332664 113692 332716
rect 160836 332664 160888 332716
rect 71872 332596 71924 332648
rect 73068 332596 73120 332648
rect 133328 332596 133380 332648
rect 133420 332596 133472 332648
rect 170496 332596 170548 332648
rect 91008 332528 91060 332580
rect 93860 332528 93912 332580
rect 207664 331848 207716 331900
rect 239404 331848 239456 331900
rect 129740 331440 129792 331492
rect 130108 331440 130160 331492
rect 53748 331304 53800 331356
rect 129740 331304 129792 331356
rect 141240 331304 141292 331356
rect 157432 331304 157484 331356
rect 107200 331236 107252 331288
rect 189724 331236 189776 331288
rect 56508 331168 56560 331220
rect 123484 331168 123536 331220
rect 78680 331100 78732 331152
rect 79324 331100 79376 331152
rect 82728 331100 82780 331152
rect 83464 331100 83516 331152
rect 95792 331100 95844 331152
rect 96436 331100 96488 331152
rect 117780 331100 117832 331152
rect 118608 331100 118660 331152
rect 118700 331100 118752 331152
rect 119436 331100 119488 331152
rect 137836 331100 137888 331152
rect 139400 331100 139452 331152
rect 144184 331100 144236 331152
rect 144828 331100 144880 331152
rect 198096 330556 198148 330608
rect 247132 330556 247184 330608
rect 25504 330488 25556 330540
rect 56508 330488 56560 330540
rect 85856 330488 85908 330540
rect 97264 330488 97316 330540
rect 101496 330488 101548 330540
rect 132592 330488 132644 330540
rect 157432 330488 157484 330540
rect 213828 330488 213880 330540
rect 107752 330352 107804 330404
rect 108028 330352 108080 330404
rect 127716 330352 127768 330404
rect 133420 330352 133472 330404
rect 139216 330352 139268 330404
rect 143448 330352 143500 330404
rect 97264 330080 97316 330132
rect 98736 330080 98788 330132
rect 100024 330080 100076 330132
rect 101404 330080 101456 330132
rect 110604 330080 110656 330132
rect 111708 330080 111760 330132
rect 88616 329944 88668 329996
rect 89628 329944 89680 329996
rect 63408 329808 63460 329860
rect 74540 329808 74592 329860
rect 136916 329808 136968 329860
rect 137928 329808 137980 329860
rect 149060 329808 149112 329860
rect 154304 329808 154356 329860
rect 154580 329808 154632 329860
rect 159364 329808 159416 329860
rect 50528 329740 50580 329792
rect 50804 329740 50856 329792
rect 135168 329740 135220 329792
rect 36544 329060 36596 329112
rect 50528 329060 50580 329112
rect 133420 329060 133472 329112
rect 184204 329060 184256 329112
rect 32404 328448 32456 328500
rect 124956 328448 125008 328500
rect 143448 328448 143500 328500
rect 147404 328448 147456 328500
rect 148968 328448 149020 328500
rect 177488 328448 177540 328500
rect 67824 328380 67876 328432
rect 71872 328380 71924 328432
rect 151728 327768 151780 327820
rect 162216 327768 162268 327820
rect 153936 327700 153988 327752
rect 164976 327700 165028 327752
rect 76472 327156 76524 327208
rect 154396 327156 154448 327208
rect 22744 327088 22796 327140
rect 122932 327088 122984 327140
rect 123668 327088 123720 327140
rect 154304 327088 154356 327140
rect 154856 327088 154908 327140
rect 68652 327020 68704 327072
rect 99380 327020 99432 327072
rect 100116 327020 100168 327072
rect 133328 327020 133380 327072
rect 141240 327020 141292 327072
rect 141424 327020 141476 327072
rect 68560 326952 68612 327004
rect 69388 326952 69440 327004
rect 70032 326952 70084 327004
rect 76564 326952 76616 327004
rect 67732 326884 67784 326936
rect 69572 326884 69624 326936
rect 152096 327020 152148 327072
rect 154396 327020 154448 327072
rect 147404 326952 147456 327004
rect 153108 326884 153160 326936
rect 154304 326884 154356 326936
rect 155868 326884 155920 326936
rect 242164 326340 242216 326392
rect 59084 325660 59136 325712
rect 67180 325660 67232 325712
rect 156420 325660 156472 325712
rect 360200 325660 360252 325712
rect 67364 325592 67416 325644
rect 67732 325592 67784 325644
rect 157156 325320 157208 325372
rect 158720 325320 158772 325372
rect 157248 324912 157300 324964
rect 203616 324912 203668 324964
rect 52368 324300 52420 324352
rect 66904 324300 66956 324352
rect 60648 322940 60700 322992
rect 66812 322940 66864 322992
rect 156880 322940 156932 322992
rect 204996 322940 205048 322992
rect 176016 322260 176068 322312
rect 189816 322260 189868 322312
rect 158720 322192 158772 322244
rect 248420 322192 248472 322244
rect 61936 321580 61988 321632
rect 157248 321580 157300 321632
rect 163688 321580 163740 321632
rect 65616 321512 65668 321564
rect 66444 321512 66496 321564
rect 155868 320900 155920 320952
rect 196624 320900 196676 320952
rect 67364 320832 67416 320884
rect 68284 320832 68336 320884
rect 178684 320832 178736 320884
rect 236644 320832 236696 320884
rect 218704 320152 218756 320204
rect 219348 320152 219400 320204
rect 295984 320152 296036 320204
rect 4068 320084 4120 320136
rect 4804 320084 4856 320136
rect 167736 319472 167788 319524
rect 206376 319472 206428 319524
rect 164884 319404 164936 319456
rect 238116 319404 238168 319456
rect 64420 318792 64472 318844
rect 66812 318792 66864 318844
rect 157248 318792 157300 318844
rect 160928 318792 160980 318844
rect 208492 318792 208544 318844
rect 209136 318792 209188 318844
rect 284944 318792 284996 318844
rect 219716 318384 219768 318436
rect 220176 318384 220228 318436
rect 11704 318044 11756 318096
rect 53840 318044 53892 318096
rect 164976 318044 165028 318096
rect 224868 318044 224920 318096
rect 56508 317500 56560 317552
rect 66812 317500 66864 317552
rect 53840 317432 53892 317484
rect 54944 317432 54996 317484
rect 66904 317432 66956 317484
rect 219716 317432 219768 317484
rect 305000 317432 305052 317484
rect 157248 317364 157300 317416
rect 161572 317364 161624 317416
rect 162768 317364 162820 317416
rect 162768 316752 162820 316804
rect 173164 316752 173216 316804
rect 178776 316752 178828 316804
rect 249064 316752 249116 316804
rect 163780 316684 163832 316736
rect 242256 316684 242308 316736
rect 63316 315936 63368 315988
rect 66812 315936 66864 315988
rect 157248 315324 157300 315376
rect 164332 315324 164384 315376
rect 35164 315256 35216 315308
rect 63316 315256 63368 315308
rect 160928 315256 160980 315308
rect 246028 315256 246080 315308
rect 156788 314644 156840 314696
rect 160744 314644 160796 314696
rect 164332 314644 164384 314696
rect 165068 314644 165120 314696
rect 224868 314644 224920 314696
rect 269764 314644 269816 314696
rect 158076 313896 158128 313948
rect 199476 313896 199528 313948
rect 226340 313352 226392 313404
rect 288440 313352 288492 313404
rect 53564 313284 53616 313336
rect 61660 313284 61712 313336
rect 66904 313284 66956 313336
rect 187056 313284 187108 313336
rect 187608 313284 187660 313336
rect 268384 313284 268436 313336
rect 64788 313216 64840 313268
rect 66812 313216 66864 313268
rect 189816 312536 189868 312588
rect 239220 312536 239272 312588
rect 246304 312536 246356 312588
rect 255412 312536 255464 312588
rect 156420 311856 156472 311908
rect 218704 311856 218756 311908
rect 220084 311856 220136 311908
rect 220728 311856 220780 311908
rect 304264 311856 304316 311908
rect 64604 311788 64656 311840
rect 66444 311788 66496 311840
rect 184296 311176 184348 311228
rect 230020 311176 230072 311228
rect 173348 311108 173400 311160
rect 236000 311108 236052 311160
rect 157248 310496 157300 310548
rect 180156 310496 180208 310548
rect 204996 310428 205048 310480
rect 209964 310428 210016 310480
rect 170496 309748 170548 309800
rect 191196 309748 191248 309800
rect 156144 309272 156196 309324
rect 158076 309272 158128 309324
rect 157248 309204 157300 309256
rect 199384 309204 199436 309256
rect 53656 309136 53708 309188
rect 66812 309136 66864 309188
rect 191288 309136 191340 309188
rect 254032 309136 254084 309188
rect 167828 309068 167880 309120
rect 168288 309068 168340 309120
rect 226340 309068 226392 309120
rect 156696 308456 156748 308508
rect 159548 308456 159600 308508
rect 14464 308388 14516 308440
rect 67640 308388 67692 308440
rect 193128 307844 193180 307896
rect 280160 307844 280212 307896
rect 228456 307776 228508 307828
rect 228916 307776 228968 307828
rect 324412 307776 324464 307828
rect 154764 307708 154816 307760
rect 155316 307708 155368 307760
rect 239220 307708 239272 307760
rect 242532 307708 242584 307760
rect 18604 307028 18656 307080
rect 66720 307028 66772 307080
rect 207756 306416 207808 306468
rect 286416 306416 286468 306468
rect 61752 306348 61804 306400
rect 66996 306348 67048 306400
rect 154764 306348 154816 306400
rect 239496 306348 239548 306400
rect 3424 306280 3476 306332
rect 36544 306280 36596 306332
rect 63224 306280 63276 306332
rect 66904 306280 66956 306332
rect 157248 306280 157300 306332
rect 160192 306280 160244 306332
rect 160192 305668 160244 305720
rect 174728 305668 174780 305720
rect 163688 305600 163740 305652
rect 245752 305600 245804 305652
rect 184388 304988 184440 305040
rect 258080 304988 258132 305040
rect 157248 304240 157300 304292
rect 183468 304240 183520 304292
rect 224316 304240 224368 304292
rect 247040 304240 247092 304292
rect 157248 303696 157300 303748
rect 215944 303696 215996 303748
rect 57888 303628 57940 303680
rect 66260 303628 66312 303680
rect 197176 303628 197228 303680
rect 198188 303628 198240 303680
rect 262956 303628 263008 303680
rect 60464 303560 60516 303612
rect 66812 303560 66864 303612
rect 183468 302268 183520 302320
rect 261484 302268 261536 302320
rect 157248 302200 157300 302252
rect 243912 302200 243964 302252
rect 64696 302132 64748 302184
rect 66812 302132 66864 302184
rect 197268 301520 197320 301572
rect 198096 301520 198148 301572
rect 193864 301316 193916 301368
rect 194508 301316 194560 301368
rect 215300 300908 215352 300960
rect 216036 300908 216088 300960
rect 267004 300908 267056 300960
rect 194508 300840 194560 300892
rect 246304 300840 246356 300892
rect 60556 300772 60608 300824
rect 66812 300772 66864 300824
rect 63316 299548 63368 299600
rect 66260 299548 66312 299600
rect 157248 299548 157300 299600
rect 244464 299548 244516 299600
rect 162400 299480 162452 299532
rect 256700 299480 256752 299532
rect 157248 299412 157300 299464
rect 165712 299412 165764 299464
rect 166080 299412 166132 299464
rect 231124 299412 231176 299464
rect 233148 299412 233200 299464
rect 214564 298800 214616 298852
rect 227444 298800 227496 298852
rect 50804 298732 50856 298784
rect 66904 298732 66956 298784
rect 166080 298732 166132 298784
rect 216588 298732 216640 298784
rect 233148 298120 233200 298172
rect 583760 298120 583812 298172
rect 238208 298052 238260 298104
rect 238668 298052 238720 298104
rect 156788 296760 156840 296812
rect 252744 296760 252796 296812
rect 238668 296692 238720 296744
rect 582564 296692 582616 296744
rect 39948 296624 40000 296676
rect 66444 296624 66496 296676
rect 157248 295944 157300 295996
rect 161480 295944 161532 295996
rect 162768 295944 162820 295996
rect 203708 295400 203760 295452
rect 277400 295400 277452 295452
rect 200580 295332 200632 295384
rect 216680 295332 216732 295384
rect 233976 295332 234028 295384
rect 582472 295332 582524 295384
rect 156420 295264 156472 295316
rect 169760 295264 169812 295316
rect 216588 294652 216640 294704
rect 228364 294652 228416 294704
rect 169760 294584 169812 294636
rect 204352 294584 204404 294636
rect 218704 294584 218756 294636
rect 245844 294584 245896 294636
rect 246304 294584 246356 294636
rect 297364 294584 297416 294636
rect 46848 294040 46900 294092
rect 66260 294040 66312 294092
rect 33784 293972 33836 294024
rect 67548 293972 67600 294024
rect 199476 293972 199528 294024
rect 218060 293972 218112 294024
rect 240876 293972 240928 294024
rect 583208 293972 583260 294024
rect 215944 293292 215996 293344
rect 236736 293292 236788 293344
rect 170404 293224 170456 293276
rect 202788 293224 202840 293276
rect 209964 293224 210016 293276
rect 235172 293224 235224 293276
rect 241520 293224 241572 293276
rect 291844 293224 291896 293276
rect 2780 292816 2832 292868
rect 4804 292816 4856 292868
rect 157248 292544 157300 292596
rect 215484 292544 215536 292596
rect 40684 292476 40736 292528
rect 66812 292476 66864 292528
rect 218060 291796 218112 291848
rect 244372 291796 244424 291848
rect 204352 291592 204404 291644
rect 208584 291592 208636 291644
rect 157248 291252 157300 291304
rect 193956 291252 194008 291304
rect 193864 291184 193916 291236
rect 223028 291184 223080 291236
rect 223580 291184 223632 291236
rect 265624 291184 265676 291236
rect 64696 291116 64748 291168
rect 65524 291116 65576 291168
rect 158076 291116 158128 291168
rect 160744 291116 160796 291168
rect 64696 289892 64748 289944
rect 66812 289892 66864 289944
rect 174544 289892 174596 289944
rect 247224 289892 247276 289944
rect 157248 289824 157300 289876
rect 244556 289824 244608 289876
rect 233884 289756 233936 289808
rect 235540 289756 235592 289808
rect 61844 289212 61896 289264
rect 66260 289212 66312 289264
rect 157248 288464 157300 288516
rect 208400 288464 208452 288516
rect 218060 288464 218112 288516
rect 220636 288464 220688 288516
rect 264244 288464 264296 288516
rect 163688 288396 163740 288448
rect 223580 288396 223632 288448
rect 236736 288396 236788 288448
rect 262864 288396 262916 288448
rect 215484 288328 215536 288380
rect 218060 288328 218112 288380
rect 208400 287648 208452 287700
rect 224684 287648 224736 287700
rect 208400 287512 208452 287564
rect 208584 287512 208636 287564
rect 224684 287104 224736 287156
rect 253204 287104 253256 287156
rect 60556 287036 60608 287088
rect 66812 287036 66864 287088
rect 164884 287036 164936 287088
rect 210884 287036 210936 287088
rect 219440 287036 219492 287088
rect 267740 287036 267792 287088
rect 159456 286288 159508 286340
rect 187056 286288 187108 286340
rect 187608 286288 187660 286340
rect 200764 286288 200816 286340
rect 218704 286288 218756 286340
rect 236460 286288 236512 286340
rect 156144 285880 156196 285932
rect 158076 285880 158128 285932
rect 219348 285880 219400 285932
rect 221188 285880 221240 285932
rect 55128 285744 55180 285796
rect 66996 285744 67048 285796
rect 48228 285676 48280 285728
rect 66812 285676 66864 285728
rect 162308 285676 162360 285728
rect 164240 285676 164292 285728
rect 195520 285676 195572 285728
rect 205548 285744 205600 285796
rect 250444 285744 250496 285796
rect 203156 285676 203208 285728
rect 204168 285676 204220 285728
rect 204904 285676 204956 285728
rect 208124 285676 208176 285728
rect 232596 285676 232648 285728
rect 234252 285676 234304 285728
rect 237564 285676 237616 285728
rect 237932 285676 237984 285728
rect 300124 285676 300176 285728
rect 156788 285608 156840 285660
rect 174544 285608 174596 285660
rect 201500 285268 201552 285320
rect 202420 285268 202472 285320
rect 208400 285268 208452 285320
rect 208676 285268 208728 285320
rect 177488 284996 177540 285048
rect 184296 284996 184348 285048
rect 159548 284928 159600 284980
rect 196716 284928 196768 284980
rect 216680 284928 216732 284980
rect 240048 284928 240100 284980
rect 216772 284724 216824 284776
rect 219440 284724 219492 284776
rect 200120 284384 200172 284436
rect 216772 284384 216824 284436
rect 230756 284384 230808 284436
rect 231124 284384 231176 284436
rect 243912 284384 243964 284436
rect 199568 284316 199620 284368
rect 217324 284316 217376 284368
rect 241980 284316 242032 284368
rect 313924 284316 313976 284368
rect 157248 284248 157300 284300
rect 191288 284248 191340 284300
rect 195980 283908 196032 283960
rect 204352 283908 204404 283960
rect 178776 283840 178828 283892
rect 200120 283840 200172 283892
rect 243912 283840 243964 283892
rect 282920 283840 282972 283892
rect 50988 282888 51040 282940
rect 66628 282888 66680 282940
rect 245384 282888 245436 282940
rect 273260 282888 273312 282940
rect 246120 282820 246172 282872
rect 251364 282820 251416 282872
rect 582840 282820 582892 282872
rect 157248 282616 157300 282668
rect 162400 282616 162452 282668
rect 173348 282208 173400 282260
rect 198740 282208 198792 282260
rect 157156 282140 157208 282192
rect 185768 282140 185820 282192
rect 56416 281528 56468 281580
rect 66352 281528 66404 281580
rect 185768 281528 185820 281580
rect 186228 281528 186280 281580
rect 197360 281528 197412 281580
rect 245660 281528 245712 281580
rect 249708 281528 249760 281580
rect 157248 281460 157300 281512
rect 184388 281460 184440 281512
rect 246120 281460 246172 281512
rect 258172 281460 258224 281512
rect 259368 281460 259420 281512
rect 174728 281392 174780 281444
rect 197360 281392 197412 281444
rect 259368 280780 259420 280832
rect 286324 280780 286376 280832
rect 63132 280168 63184 280220
rect 66812 280168 66864 280220
rect 245660 280168 245712 280220
rect 298744 280168 298796 280220
rect 183468 280100 183520 280152
rect 197360 280100 197412 280152
rect 156972 279624 157024 279676
rect 160928 279624 160980 279676
rect 173440 279420 173492 279472
rect 197452 279420 197504 279472
rect 249708 279420 249760 279472
rect 266360 279420 266412 279472
rect 29644 278740 29696 278792
rect 60464 278740 60516 278792
rect 66628 278740 66680 278792
rect 157064 278740 157116 278792
rect 175188 278740 175240 278792
rect 246120 278740 246172 278792
rect 251364 278740 251416 278792
rect 583576 278740 583628 278792
rect 173256 277992 173308 278044
rect 197268 277992 197320 278044
rect 246120 277992 246172 278044
rect 249984 277992 250036 278044
rect 583392 277992 583444 278044
rect 156512 277380 156564 277432
rect 187056 277380 187108 277432
rect 175188 277312 175240 277364
rect 193128 277312 193180 277364
rect 193128 277108 193180 277160
rect 197360 277108 197412 277160
rect 155316 276632 155368 276684
rect 198004 276632 198056 276684
rect 246028 276632 246080 276684
rect 282184 276632 282236 276684
rect 245844 276224 245896 276276
rect 246028 276224 246080 276276
rect 244280 276088 244332 276140
rect 245660 276088 245712 276140
rect 157248 275952 157300 276004
rect 198280 275952 198332 276004
rect 245936 275952 245988 276004
rect 249892 275952 249944 276004
rect 582656 275952 582708 276004
rect 157248 274660 157300 274712
rect 169208 274660 169260 274712
rect 183100 274660 183152 274712
rect 197452 274660 197504 274712
rect 168288 274592 168340 274644
rect 197360 274592 197412 274644
rect 57612 273912 57664 273964
rect 66260 273912 66312 273964
rect 245936 273912 245988 273964
rect 327172 273912 327224 273964
rect 157248 273232 157300 273284
rect 166448 273232 166500 273284
rect 180248 273232 180300 273284
rect 197360 273232 197412 273284
rect 245844 273232 245896 273284
rect 249892 273232 249944 273284
rect 245936 272552 245988 272604
rect 251272 272552 251324 272604
rect 251824 272552 251876 272604
rect 169116 272484 169168 272536
rect 195888 272484 195940 272536
rect 245844 272484 245896 272536
rect 325700 272484 325752 272536
rect 61752 271940 61804 271992
rect 66996 271940 67048 271992
rect 52184 271872 52236 271924
rect 66812 271872 66864 271924
rect 157248 271872 157300 271924
rect 192484 271872 192536 271924
rect 195888 271872 195940 271924
rect 197360 271872 197412 271924
rect 162492 271124 162544 271176
rect 178776 271124 178828 271176
rect 245752 271124 245804 271176
rect 248604 271124 248656 271176
rect 253204 271124 253256 271176
rect 274640 271124 274692 271176
rect 193036 270580 193088 270632
rect 197452 270580 197504 270632
rect 53748 270512 53800 270564
rect 66812 270512 66864 270564
rect 157248 270512 157300 270564
rect 174544 270512 174596 270564
rect 183008 270512 183060 270564
rect 197360 270512 197412 270564
rect 245660 270444 245712 270496
rect 249064 270512 249116 270564
rect 280252 270512 280304 270564
rect 4068 269764 4120 269816
rect 35900 269764 35952 269816
rect 245936 269764 245988 269816
rect 312176 269764 312228 269816
rect 157248 269152 157300 269204
rect 166264 269152 166316 269204
rect 178868 269152 178920 269204
rect 197360 269152 197412 269204
rect 64512 269084 64564 269136
rect 66444 269084 66496 269136
rect 156788 269084 156840 269136
rect 199660 269084 199712 269136
rect 156512 269016 156564 269068
rect 163688 269016 163740 269068
rect 165068 269016 165120 269068
rect 197360 269016 197412 269068
rect 158168 268336 158220 268388
rect 171232 268336 171284 268388
rect 172428 268336 172480 268388
rect 185584 268336 185636 268388
rect 199568 268336 199620 268388
rect 245936 268336 245988 268388
rect 256792 268336 256844 268388
rect 244464 267724 244516 267776
rect 331312 267724 331364 267776
rect 62028 267656 62080 267708
rect 66444 267656 66496 267708
rect 157248 267656 157300 267708
rect 199476 267656 199528 267708
rect 195428 267452 195480 267504
rect 197360 267452 197412 267504
rect 3424 266976 3476 267028
rect 15844 266976 15896 267028
rect 52092 266976 52144 267028
rect 66904 266976 66956 267028
rect 177396 266976 177448 267028
rect 195060 266976 195112 267028
rect 245936 266976 245988 267028
rect 262220 266976 262272 267028
rect 246028 266364 246080 266416
rect 250076 266364 250128 266416
rect 186964 266296 187016 266348
rect 197360 266296 197412 266348
rect 245752 266296 245804 266348
rect 254124 266296 254176 266348
rect 583116 266296 583168 266348
rect 245844 266228 245896 266280
rect 255412 266228 255464 266280
rect 162400 265616 162452 265668
rect 192576 265616 192628 265668
rect 255412 265616 255464 265668
rect 274732 265616 274784 265668
rect 177856 265140 177908 265192
rect 183100 265140 183152 265192
rect 41328 264936 41380 264988
rect 66812 264936 66864 264988
rect 157248 264936 157300 264988
rect 171876 264936 171928 264988
rect 184204 264868 184256 264920
rect 197360 264868 197412 264920
rect 245936 264868 245988 264920
rect 251180 264868 251232 264920
rect 55036 264188 55088 264240
rect 65984 264188 66036 264240
rect 66444 264188 66496 264240
rect 159548 264188 159600 264240
rect 178684 264188 178736 264240
rect 55036 263644 55088 263696
rect 66812 263644 66864 263696
rect 163688 263576 163740 263628
rect 193128 263576 193180 263628
rect 197360 263576 197412 263628
rect 245844 263576 245896 263628
rect 262220 263576 262272 263628
rect 194048 262896 194100 262948
rect 195520 262896 195572 262948
rect 52276 262828 52328 262880
rect 62120 262828 62172 262880
rect 256792 262828 256844 262880
rect 582656 262828 582708 262880
rect 178684 262284 178736 262336
rect 197360 262284 197412 262336
rect 62120 262216 62172 262268
rect 63224 262216 63276 262268
rect 66812 262216 66864 262268
rect 157248 262216 157300 262268
rect 184204 262216 184256 262268
rect 245936 262216 245988 262268
rect 251180 262216 251232 262268
rect 156788 262148 156840 262200
rect 165620 262148 165672 262200
rect 35900 261468 35952 261520
rect 58992 261468 59044 261520
rect 250444 261468 250496 261520
rect 303620 261468 303672 261520
rect 185676 260924 185728 260976
rect 197360 260924 197412 260976
rect 58992 260856 59044 260908
rect 66812 260856 66864 260908
rect 173256 260856 173308 260908
rect 197452 260856 197504 260908
rect 244924 260856 244976 260908
rect 288532 260856 288584 260908
rect 245936 260788 245988 260840
rect 252744 260788 252796 260840
rect 253020 260788 253072 260840
rect 245844 260176 245896 260228
rect 276020 260176 276072 260228
rect 162216 260108 162268 260160
rect 189908 260108 189960 260160
rect 253020 260108 253072 260160
rect 306656 260108 306708 260160
rect 155408 259428 155460 259480
rect 182088 259428 182140 259480
rect 197360 259428 197412 259480
rect 195060 259360 195112 259412
rect 197452 259360 197504 259412
rect 245844 259360 245896 259412
rect 258080 259360 258132 259412
rect 259368 259360 259420 259412
rect 245936 258680 245988 258732
rect 254032 258680 254084 258732
rect 259368 258680 259420 258732
rect 293224 258680 293276 258732
rect 191748 258476 191800 258528
rect 197360 258476 197412 258528
rect 56324 258136 56376 258188
rect 66352 258136 66404 258188
rect 43904 258068 43956 258120
rect 66812 258068 66864 258120
rect 156604 258068 156656 258120
rect 162124 258068 162176 258120
rect 189724 258068 189776 258120
rect 191748 258068 191800 258120
rect 66352 258000 66404 258052
rect 68100 258000 68152 258052
rect 157248 257932 157300 257984
rect 162492 257932 162544 257984
rect 247224 257320 247276 257372
rect 322940 257320 322992 257372
rect 61844 256708 61896 256760
rect 66444 256708 66496 256760
rect 157248 256708 157300 256760
rect 171048 256708 171100 256760
rect 173440 256708 173492 256760
rect 175832 256708 175884 256760
rect 183468 256708 183520 256760
rect 197360 256708 197412 256760
rect 178776 256028 178828 256080
rect 183008 256028 183060 256080
rect 159640 255960 159692 256012
rect 181628 255960 181680 256012
rect 157248 255280 157300 255332
rect 165528 255280 165580 255332
rect 187240 255280 187292 255332
rect 197360 255280 197412 255332
rect 3424 255212 3476 255264
rect 14464 255212 14516 255264
rect 157248 254532 157300 254584
rect 189724 254532 189776 254584
rect 254032 254532 254084 254584
rect 305092 254532 305144 254584
rect 52276 253920 52328 253972
rect 66444 253920 66496 253972
rect 188528 253920 188580 253972
rect 197360 253920 197412 253972
rect 246028 253920 246080 253972
rect 249984 253920 250036 253972
rect 157248 253852 157300 253904
rect 175832 253852 175884 253904
rect 194508 253852 194560 253904
rect 197452 253852 197504 253904
rect 245936 253852 245988 253904
rect 256700 253852 256752 253904
rect 256884 253852 256936 253904
rect 167644 253172 167696 253224
rect 177396 253172 177448 253224
rect 256884 253172 256936 253224
rect 327264 253172 327316 253224
rect 245936 252832 245988 252884
rect 248512 252832 248564 252884
rect 249064 252832 249116 252884
rect 59176 252628 59228 252680
rect 64604 252628 64656 252680
rect 66628 252628 66680 252680
rect 245752 252424 245804 252476
rect 255320 252424 255372 252476
rect 165528 251812 165580 251864
rect 184848 251812 184900 251864
rect 255320 251812 255372 251864
rect 522304 251812 522356 251864
rect 192576 251268 192628 251320
rect 197452 251268 197504 251320
rect 157248 251200 157300 251252
rect 168380 251200 168432 251252
rect 184848 251200 184900 251252
rect 197360 251200 197412 251252
rect 156144 250452 156196 250504
rect 174728 250452 174780 250504
rect 287704 250452 287756 250504
rect 317512 250452 317564 250504
rect 195336 249908 195388 249960
rect 197452 249908 197504 249960
rect 157248 249772 157300 249824
rect 176108 249772 176160 249824
rect 178960 249772 179012 249824
rect 197360 249772 197412 249824
rect 245752 249772 245804 249824
rect 255320 249772 255372 249824
rect 192484 249704 192536 249756
rect 193036 249704 193088 249756
rect 197452 249704 197504 249756
rect 245936 249500 245988 249552
rect 249800 249500 249852 249552
rect 157248 249432 157300 249484
rect 163688 249432 163740 249484
rect 181996 249024 182048 249076
rect 195336 249024 195388 249076
rect 268384 249024 268436 249076
rect 334072 249024 334124 249076
rect 173164 248888 173216 248940
rect 178868 248888 178920 248940
rect 62028 248412 62080 248464
rect 66812 248412 66864 248464
rect 157156 248412 157208 248464
rect 174176 248412 174228 248464
rect 157248 247732 157300 247784
rect 165528 247732 165580 247784
rect 169208 247732 169260 247784
rect 191288 247732 191340 247784
rect 158076 247664 158128 247716
rect 192576 247664 192628 247716
rect 245936 247664 245988 247716
rect 246120 247664 246172 247716
rect 583300 247664 583352 247716
rect 59176 247052 59228 247104
rect 66812 247052 66864 247104
rect 166356 247052 166408 247104
rect 167736 247052 167788 247104
rect 194140 247052 194192 247104
rect 197360 247052 197412 247104
rect 191104 246984 191156 247036
rect 197452 246984 197504 247036
rect 244924 246304 244976 246356
rect 269120 246304 269172 246356
rect 166540 245692 166592 245744
rect 188988 245692 189040 245744
rect 197360 245692 197412 245744
rect 157248 245624 157300 245676
rect 180064 245624 180116 245676
rect 246396 245624 246448 245676
rect 247040 245624 247092 245676
rect 302240 245624 302292 245676
rect 57704 244876 57756 244928
rect 67180 244876 67232 244928
rect 280804 244876 280856 244928
rect 310520 244876 310572 244928
rect 188436 244332 188488 244384
rect 157984 244264 158036 244316
rect 189080 244264 189132 244316
rect 189908 244332 189960 244384
rect 191656 244332 191708 244384
rect 197452 244332 197504 244384
rect 190368 244264 190420 244316
rect 197360 244264 197412 244316
rect 245936 244264 245988 244316
rect 258080 244264 258132 244316
rect 174176 243516 174228 243568
rect 199568 243516 199620 243568
rect 286416 243516 286468 243568
rect 321652 243516 321704 243568
rect 156144 242972 156196 243024
rect 158076 242972 158128 243024
rect 157248 242904 157300 242956
rect 189908 242904 189960 242956
rect 246396 242904 246448 242956
rect 247224 242904 247276 242956
rect 286508 242904 286560 242956
rect 166448 242156 166500 242208
rect 184388 242156 184440 242208
rect 244280 242156 244332 242208
rect 329932 242156 329984 242208
rect 65984 242020 66036 242072
rect 71044 242020 71096 242072
rect 152464 242020 152516 242072
rect 155224 242020 155276 242072
rect 69756 241816 69808 241868
rect 72424 241816 72476 241868
rect 153844 241476 153896 241528
rect 192944 241476 192996 241528
rect 195796 241476 195848 241528
rect 197912 241476 197964 241528
rect 246304 241476 246356 241528
rect 247132 241476 247184 241528
rect 320272 241476 320324 241528
rect 3424 241408 3476 241460
rect 32404 241408 32456 241460
rect 105038 241408 105090 241460
rect 155408 241408 155460 241460
rect 67456 240796 67508 240848
rect 81256 240796 81308 240848
rect 258724 240796 258776 240848
rect 278044 240796 278096 240848
rect 64512 240728 64564 240780
rect 103612 240728 103664 240780
rect 121000 240728 121052 240780
rect 200120 240728 200172 240780
rect 244096 240728 244148 240780
rect 580264 240728 580316 240780
rect 199936 240456 199988 240508
rect 196624 240388 196676 240440
rect 200120 240320 200172 240372
rect 200304 240116 200356 240168
rect 201040 240116 201092 240168
rect 201408 240116 201460 240168
rect 231952 240116 232004 240168
rect 235816 240116 235868 240168
rect 245752 240116 245804 240168
rect 256700 240116 256752 240168
rect 86040 240048 86092 240100
rect 86868 240048 86920 240100
rect 91928 240048 91980 240100
rect 92388 240048 92440 240100
rect 101128 240048 101180 240100
rect 101956 240048 102008 240100
rect 115296 240048 115348 240100
rect 115848 240048 115900 240100
rect 118792 240048 118844 240100
rect 119988 240048 120040 240100
rect 121736 240048 121788 240100
rect 122748 240048 122800 240100
rect 124680 240048 124732 240100
rect 125508 240048 125560 240100
rect 128912 240048 128964 240100
rect 129648 240048 129700 240100
rect 130384 240048 130436 240100
rect 130936 240048 130988 240100
rect 249708 240048 249760 240100
rect 250076 240048 250128 240100
rect 96896 239980 96948 240032
rect 101496 239980 101548 240032
rect 114652 239980 114704 240032
rect 115388 239980 115440 240032
rect 116768 239980 116820 240032
rect 124312 239980 124364 240032
rect 75368 239912 75420 239964
rect 75828 239912 75880 239964
rect 88984 239912 89036 239964
rect 89536 239912 89588 239964
rect 90456 239912 90508 239964
rect 90916 239912 90968 239964
rect 147772 239912 147824 239964
rect 148324 239912 148376 239964
rect 106832 239776 106884 239828
rect 107568 239776 107620 239828
rect 109592 239776 109644 239828
rect 110328 239776 110380 239828
rect 68928 239504 68980 239556
rect 70308 239504 70360 239556
rect 81532 239504 81584 239556
rect 82728 239504 82780 239556
rect 99380 239504 99432 239556
rect 100668 239504 100720 239556
rect 70216 239436 70268 239488
rect 108304 239436 108356 239488
rect 110236 239436 110288 239488
rect 115204 239436 115256 239488
rect 149704 239436 149756 239488
rect 240324 239436 240376 239488
rect 79048 239368 79100 239420
rect 79968 239368 80020 239420
rect 80520 239368 80572 239420
rect 88984 239368 89036 239420
rect 108212 239368 108264 239420
rect 208400 239368 208452 239420
rect 102600 239232 102652 239284
rect 103336 239232 103388 239284
rect 107752 239232 107804 239284
rect 108396 239232 108448 239284
rect 111064 239232 111116 239284
rect 111708 239232 111760 239284
rect 131856 239232 131908 239284
rect 132316 239232 132368 239284
rect 144000 239232 144052 239284
rect 144736 239232 144788 239284
rect 153936 239232 153988 239284
rect 154488 239232 154540 239284
rect 145288 239096 145340 239148
rect 145932 239096 145984 239148
rect 148232 239096 148284 239148
rect 148968 239096 149020 239148
rect 133144 238960 133196 239012
rect 133696 238960 133748 239012
rect 134616 238960 134668 239012
rect 135168 238960 135220 239012
rect 74448 238756 74500 238808
rect 75460 238756 75512 238808
rect 83096 238688 83148 238740
rect 207664 238688 207716 238740
rect 208400 238688 208452 238740
rect 219900 238688 219952 238740
rect 220820 238688 220872 238740
rect 222292 238688 222344 238740
rect 101496 238620 101548 238672
rect 214196 238620 214248 238672
rect 216588 238348 216640 238400
rect 218060 238348 218112 238400
rect 67916 238076 67968 238128
rect 79324 238076 79376 238128
rect 224776 238076 224828 238128
rect 226708 238076 226760 238128
rect 67364 238008 67416 238060
rect 98552 238008 98604 238060
rect 226984 238008 227036 238060
rect 238852 238008 238904 238060
rect 240324 238008 240376 238060
rect 301504 238008 301556 238060
rect 218152 237464 218204 237516
rect 218704 237464 218756 237516
rect 220084 237464 220136 237516
rect 221924 237464 221976 237516
rect 222292 237464 222344 237516
rect 222844 237464 222896 237516
rect 222936 237464 222988 237516
rect 223764 237464 223816 237516
rect 233884 237396 233936 237448
rect 237380 237396 237432 237448
rect 240784 237396 240836 237448
rect 243268 237396 243320 237448
rect 244280 237396 244332 237448
rect 4804 237328 4856 237380
rect 54852 237328 54904 237380
rect 136640 237328 136692 237380
rect 138112 237328 138164 237380
rect 160928 237328 160980 237380
rect 189724 237328 189776 237380
rect 242716 237328 242768 237380
rect 81256 236648 81308 236700
rect 248328 236648 248380 236700
rect 136640 235968 136692 236020
rect 137284 235968 137336 236020
rect 103612 235900 103664 235952
rect 180248 235900 180300 235952
rect 199568 235900 199620 235952
rect 243636 235900 243688 235952
rect 146024 235424 146076 235476
rect 153844 235424 153896 235476
rect 61936 235288 61988 235340
rect 75184 235288 75236 235340
rect 61752 235220 61804 235272
rect 124588 235220 124640 235272
rect 126796 235220 126848 235272
rect 135260 235220 135312 235272
rect 176108 235220 176160 235272
rect 198740 235220 198792 235272
rect 243636 235220 243688 235272
rect 260104 235220 260156 235272
rect 284944 235220 284996 235272
rect 301596 235220 301648 235272
rect 234068 234608 234120 234660
rect 321560 234608 321612 234660
rect 153016 234540 153068 234592
rect 159364 234540 159416 234592
rect 198740 234540 198792 234592
rect 247224 234540 247276 234592
rect 191196 234472 191248 234524
rect 204168 234472 204220 234524
rect 114652 233928 114704 233980
rect 139216 233928 139268 233980
rect 139400 233928 139452 233980
rect 147680 233928 147732 233980
rect 63132 233860 63184 233912
rect 104164 233860 104216 233912
rect 107752 233860 107804 233912
rect 146944 233860 146996 233912
rect 147772 233860 147824 233912
rect 177948 233860 178000 233912
rect 178776 233860 178828 233912
rect 204168 233860 204220 233912
rect 214656 233860 214708 233912
rect 215944 233792 215996 233844
rect 221004 233792 221056 233844
rect 222108 233792 222160 233844
rect 159456 233248 159508 233300
rect 185676 233248 185728 233300
rect 240784 233248 240836 233300
rect 331404 233248 331456 233300
rect 98552 233180 98604 233232
rect 155592 233180 155644 233232
rect 187056 233180 187108 233232
rect 220452 233180 220504 233232
rect 220728 233180 220780 233232
rect 124588 233112 124640 233164
rect 139400 233112 139452 233164
rect 146944 233112 146996 233164
rect 159548 233112 159600 233164
rect 199384 233112 199436 233164
rect 214564 233112 214616 233164
rect 215116 233112 215168 233164
rect 58992 232500 59044 232552
rect 123484 232500 123536 232552
rect 214196 232500 214248 232552
rect 258816 232500 258868 232552
rect 232044 231888 232096 231940
rect 233148 231888 233200 231940
rect 314660 231820 314712 231872
rect 15844 231752 15896 231804
rect 92480 231752 92532 231804
rect 93860 231752 93912 231804
rect 94504 231752 94556 231804
rect 135996 231752 136048 231804
rect 147588 231752 147640 231804
rect 155316 231752 155368 231804
rect 155868 231752 155920 231804
rect 216680 231752 216732 231804
rect 136548 231684 136600 231736
rect 176660 231684 176712 231736
rect 189908 231684 189960 231736
rect 241244 231684 241296 231736
rect 241428 231684 241480 231736
rect 128360 231616 128412 231668
rect 146024 231616 146076 231668
rect 220728 231140 220780 231192
rect 253296 231140 253348 231192
rect 92480 231072 92532 231124
rect 93124 231072 93176 231124
rect 176660 231072 176712 231124
rect 177856 231072 177908 231124
rect 188436 231072 188488 231124
rect 241428 231072 241480 231124
rect 318892 231072 318944 231124
rect 71044 230392 71096 230444
rect 176016 230392 176068 230444
rect 200304 230392 200356 230444
rect 202144 230392 202196 230444
rect 137928 230324 137980 230376
rect 233148 230324 233200 230376
rect 66076 229712 66128 229764
rect 97264 229712 97316 229764
rect 184388 229712 184440 229764
rect 200120 229712 200172 229764
rect 221464 229712 221516 229764
rect 229652 229712 229704 229764
rect 249064 229712 249116 229764
rect 328552 229712 328604 229764
rect 57612 229032 57664 229084
rect 178684 229032 178736 229084
rect 180156 229032 180208 229084
rect 206836 229032 206888 229084
rect 79876 228964 79928 229016
rect 173348 228964 173400 229016
rect 211068 228420 211120 228472
rect 247132 228420 247184 228472
rect 220176 228352 220228 228404
rect 316224 228352 316276 228404
rect 206928 227876 206980 227928
rect 208308 227876 208360 227928
rect 106924 227672 106976 227724
rect 206284 227740 206336 227792
rect 206836 227740 206888 227792
rect 48136 227604 48188 227656
rect 118884 227604 118936 227656
rect 142068 227604 142120 227656
rect 155500 227604 155552 227656
rect 192576 227604 192628 227656
rect 222936 227604 222988 227656
rect 211804 226312 211856 226364
rect 582656 226312 582708 226364
rect 123024 226244 123076 226296
rect 173164 226244 173216 226296
rect 173348 226244 173400 226296
rect 184296 226244 184348 226296
rect 222384 226244 222436 226296
rect 174728 226176 174780 226228
rect 211068 226176 211120 226228
rect 146116 225564 146168 225616
rect 178684 225564 178736 225616
rect 222384 225020 222436 225072
rect 223028 225020 223080 225072
rect 229100 225020 229152 225072
rect 229744 225020 229796 225072
rect 313372 225020 313424 225072
rect 580908 225020 580960 225072
rect 583576 225020 583628 225072
rect 209872 224952 209924 225004
rect 583024 224952 583076 225004
rect 130936 224884 130988 224936
rect 185584 224884 185636 224936
rect 194508 224272 194560 224324
rect 307760 224272 307812 224324
rect 82728 224204 82780 224256
rect 195152 224204 195204 224256
rect 204996 224204 205048 224256
rect 582748 224204 582800 224256
rect 86960 223524 87012 223576
rect 164884 223524 164936 223576
rect 195152 223524 195204 223576
rect 276020 223524 276072 223576
rect 119988 223456 120040 223508
rect 187240 223456 187292 223508
rect 193036 222912 193088 222964
rect 218704 222912 218756 222964
rect 169024 222844 169076 222896
rect 195152 222844 195204 222896
rect 97264 222096 97316 222148
rect 195060 222096 195112 222148
rect 195152 222096 195204 222148
rect 219624 222096 219676 222148
rect 214656 221484 214708 221536
rect 233976 221484 234028 221536
rect 238668 221484 238720 221536
rect 267832 221484 267884 221536
rect 133880 221416 133932 221468
rect 215208 221416 215260 221468
rect 232688 221416 232740 221468
rect 282092 221416 282144 221468
rect 75828 220736 75880 220788
rect 172428 220736 172480 220788
rect 191288 220736 191340 220788
rect 249984 220736 250036 220788
rect 251088 220736 251140 220788
rect 49608 220668 49660 220720
rect 94504 220668 94556 220720
rect 251088 220124 251140 220176
rect 281540 220124 281592 220176
rect 14464 220056 14516 220108
rect 49608 220056 49660 220108
rect 104164 220056 104216 220108
rect 191840 220056 191892 220108
rect 200028 220056 200080 220108
rect 266544 220056 266596 220108
rect 282092 220056 282144 220108
rect 298836 220056 298888 220108
rect 195796 219444 195848 219496
rect 198096 219444 198148 219496
rect 99472 219376 99524 219428
rect 212632 219376 212684 219428
rect 215208 218832 215260 218884
rect 245568 218832 245620 218884
rect 224224 218764 224276 218816
rect 270776 218764 270828 218816
rect 122656 218696 122708 218748
rect 224868 218696 224920 218748
rect 52184 217948 52236 218000
rect 159456 217948 159508 218000
rect 122840 217880 122892 217932
rect 217324 217880 217376 217932
rect 258816 217268 258868 217320
rect 335544 217268 335596 217320
rect 81624 216588 81676 216640
rect 181996 216656 182048 216708
rect 191196 216656 191248 216708
rect 192576 216656 192628 216708
rect 249892 216656 249944 216708
rect 250628 216656 250680 216708
rect 178684 216520 178736 216572
rect 262220 216520 262272 216572
rect 103428 216452 103480 216504
rect 178040 216452 178092 216504
rect 204996 215908 205048 215960
rect 240784 215908 240836 215960
rect 286324 215908 286376 215960
rect 316132 215908 316184 215960
rect 262220 215296 262272 215348
rect 262956 215296 263008 215348
rect 3332 215228 3384 215280
rect 22744 215228 22796 215280
rect 132316 215228 132368 215280
rect 256700 215228 256752 215280
rect 144736 215160 144788 215212
rect 236000 215160 236052 215212
rect 256700 214752 256752 214804
rect 257344 214752 257396 214804
rect 158076 213868 158128 213920
rect 269120 213868 269172 213920
rect 171876 213800 171928 213852
rect 247040 213800 247092 213852
rect 46848 213188 46900 213240
rect 171968 213188 172020 213240
rect 113088 211828 113140 211880
rect 194784 211828 194836 211880
rect 39304 211760 39356 211812
rect 164240 211760 164292 211812
rect 193128 211760 193180 211812
rect 242164 211760 242216 211812
rect 191656 211080 191708 211132
rect 288624 211148 288676 211200
rect 193128 211012 193180 211064
rect 194140 211012 194192 211064
rect 151084 210536 151136 210588
rect 191104 210536 191156 210588
rect 131028 210468 131080 210520
rect 193128 210468 193180 210520
rect 70400 210400 70452 210452
rect 150440 210400 150492 210452
rect 212632 210400 212684 210452
rect 258816 210400 258868 210452
rect 278044 210400 278096 210452
rect 294696 210400 294748 210452
rect 69020 209720 69072 209772
rect 231124 209720 231176 209772
rect 92388 209652 92440 209704
rect 209044 209652 209096 209704
rect 231124 209040 231176 209092
rect 277492 209040 277544 209092
rect 208400 208360 208452 208412
rect 209688 208360 209740 208412
rect 281632 208360 281684 208412
rect 53656 208292 53708 208344
rect 244280 208292 244332 208344
rect 85580 207612 85632 207664
rect 214656 207612 214708 207664
rect 218980 207612 219032 207664
rect 311992 207612 312044 207664
rect 244280 207000 244332 207052
rect 244924 207000 244976 207052
rect 89536 206932 89588 206984
rect 192576 206932 192628 206984
rect 194784 206932 194836 206984
rect 258080 206932 258132 206984
rect 259368 206932 259420 206984
rect 110328 206864 110380 206916
rect 184296 206864 184348 206916
rect 259368 206320 259420 206372
rect 278780 206320 278832 206372
rect 222844 206252 222896 206304
rect 308404 206252 308456 206304
rect 125416 205572 125468 205624
rect 251180 205572 251232 205624
rect 252468 205572 252520 205624
rect 72424 204892 72476 204944
rect 233148 204892 233200 204944
rect 234436 204892 234488 204944
rect 252468 204892 252520 204944
rect 273352 204892 273404 204944
rect 67180 204212 67232 204264
rect 213736 204212 213788 204264
rect 150440 204144 150492 204196
rect 215668 204144 215720 204196
rect 214564 203532 214616 203584
rect 264060 203532 264112 203584
rect 3424 202784 3476 202836
rect 126796 202784 126848 202836
rect 97816 202716 97868 202768
rect 157984 202716 158036 202768
rect 154488 202172 154540 202224
rect 173256 202172 173308 202224
rect 201316 202172 201368 202224
rect 276020 202172 276072 202224
rect 171048 202104 171100 202156
rect 292028 202104 292080 202156
rect 77208 201424 77260 201476
rect 221372 201424 221424 201476
rect 144828 201356 144880 201408
rect 204996 201356 205048 201408
rect 226156 200812 226208 200864
rect 314752 200812 314804 200864
rect 206376 200744 206428 200796
rect 304264 200744 304316 200796
rect 139308 200064 139360 200116
rect 166264 200064 166316 200116
rect 203524 199452 203576 199504
rect 320364 199452 320416 199504
rect 111616 199384 111668 199436
rect 233884 199384 233936 199436
rect 115204 198636 115256 198688
rect 186964 198636 187016 198688
rect 207664 198024 207716 198076
rect 297456 198024 297508 198076
rect 183468 197956 183520 198008
rect 306472 197956 306524 198008
rect 74448 197276 74500 197328
rect 200764 197276 200816 197328
rect 201408 196664 201460 196716
rect 300216 196664 300268 196716
rect 148968 196596 149020 196648
rect 182824 196596 182876 196648
rect 186964 196596 187016 196648
rect 314844 196596 314896 196648
rect 52276 195916 52328 195968
rect 207756 195916 207808 195968
rect 122748 195236 122800 195288
rect 185584 195236 185636 195288
rect 186228 195236 186280 195288
rect 264336 195236 264388 195288
rect 247776 194556 247828 194608
rect 284300 194556 284352 194608
rect 93124 194488 93176 194540
rect 212724 194488 212776 194540
rect 233976 193876 234028 193928
rect 285680 193876 285732 193928
rect 100668 193808 100720 193860
rect 236644 193808 236696 193860
rect 156604 192516 156656 192568
rect 202328 192516 202380 192568
rect 242256 192516 242308 192568
rect 325884 192516 325936 192568
rect 132408 192448 132460 192500
rect 178776 192448 178828 192500
rect 201500 192448 201552 192500
rect 310612 192448 310664 192500
rect 97908 191088 97960 191140
rect 251180 191088 251232 191140
rect 106188 190476 106240 190528
rect 217324 190476 217376 190528
rect 242164 189796 242216 189848
rect 269396 189796 269448 189848
rect 217416 189728 217468 189780
rect 305184 189728 305236 189780
rect 3516 188980 3568 189032
rect 35164 188980 35216 189032
rect 67548 188980 67600 189032
rect 218428 188980 218480 189032
rect 178868 188300 178920 188352
rect 232596 188300 232648 188352
rect 233148 188300 233200 188352
rect 265072 188300 265124 188352
rect 294696 188300 294748 188352
rect 302332 188300 302384 188352
rect 251824 187688 251876 187740
rect 283104 187688 283156 187740
rect 298836 187076 298888 187128
rect 302424 187076 302476 187128
rect 202144 187008 202196 187060
rect 309416 187008 309468 187060
rect 115848 186940 115900 186992
rect 242164 186940 242216 186992
rect 254584 186940 254636 186992
rect 276112 186940 276164 186992
rect 119988 186328 120040 186380
rect 164884 186328 164936 186380
rect 302332 185784 302384 185836
rect 304448 185784 304500 185836
rect 190368 185648 190420 185700
rect 310796 185648 310848 185700
rect 91008 185580 91060 185632
rect 231124 185580 231176 185632
rect 121368 184900 121420 184952
rect 167920 184900 167972 184952
rect 245568 184220 245620 184272
rect 265256 184220 265308 184272
rect 301596 184220 301648 184272
rect 313464 184220 313516 184272
rect 177948 184152 178000 184204
rect 277584 184152 277636 184204
rect 286508 184152 286560 184204
rect 312084 184152 312136 184204
rect 148968 183608 149020 183660
rect 167644 183608 167696 183660
rect 129648 183540 129700 183592
rect 233976 183540 234028 183592
rect 304356 183472 304408 183524
rect 305276 183472 305328 183524
rect 261576 182860 261628 182912
rect 276204 182860 276256 182912
rect 276664 182860 276716 182912
rect 303804 182860 303856 182912
rect 184848 182792 184900 182844
rect 323124 182792 323176 182844
rect 103336 182248 103388 182300
rect 170496 182248 170548 182300
rect 113732 182180 113784 182232
rect 231216 182180 231268 182232
rect 302424 182112 302476 182164
rect 303712 182112 303764 182164
rect 238024 181500 238076 181552
rect 270592 181500 270644 181552
rect 296076 181500 296128 181552
rect 308036 181500 308088 181552
rect 167828 181432 167880 181484
rect 203524 181432 203576 181484
rect 203616 181432 203668 181484
rect 301044 181432 301096 181484
rect 308404 181432 308456 181484
rect 321744 181432 321796 181484
rect 132500 180888 132552 180940
rect 169116 180888 169168 180940
rect 126060 180820 126112 180872
rect 166448 180820 166500 180872
rect 262864 180140 262916 180192
rect 272064 180140 272116 180192
rect 293224 180140 293276 180192
rect 310704 180140 310756 180192
rect 253296 180072 253348 180124
rect 269304 180072 269356 180124
rect 290464 180072 290516 180124
rect 313556 180072 313608 180124
rect 313924 179868 313976 179920
rect 317696 179868 317748 179920
rect 118516 179460 118568 179512
rect 184388 179460 184440 179512
rect 132408 179392 132460 179444
rect 231584 179392 231636 179444
rect 180248 179324 180300 179376
rect 258080 179324 258132 179376
rect 574744 179324 574796 179376
rect 580172 179324 580224 179376
rect 292028 178712 292080 178764
rect 301412 178712 301464 178764
rect 253204 178644 253256 178696
rect 273444 178644 273496 178696
rect 301504 178644 301556 178696
rect 319076 178644 319128 178696
rect 124496 178100 124548 178152
rect 164976 178100 165028 178152
rect 115848 178032 115900 178084
rect 173440 178032 173492 178084
rect 259736 178032 259788 178084
rect 270500 178032 270552 178084
rect 227720 177964 227772 178016
rect 237380 177964 237432 178016
rect 127624 177692 127676 177744
rect 132500 177692 132552 177744
rect 257344 177352 257396 177404
rect 264980 177352 265032 177404
rect 305276 177352 305328 177404
rect 311900 177352 311952 177404
rect 250628 177284 250680 177336
rect 264244 177284 264296 177336
rect 264336 177284 264388 177336
rect 272156 177284 272208 177336
rect 282184 177284 282236 177336
rect 302424 177284 302476 177336
rect 307024 177284 307076 177336
rect 316316 177284 316368 177336
rect 102048 176876 102100 176928
rect 105452 176876 105504 176928
rect 298744 176876 298796 176928
rect 305276 176876 305328 176928
rect 134432 176740 134484 176792
rect 143448 176740 143500 176792
rect 158996 176740 159048 176792
rect 178868 176740 178920 176792
rect 136088 176672 136140 176724
rect 249524 176604 249576 176656
rect 264428 176604 264480 176656
rect 269212 176604 269264 176656
rect 262956 176536 263008 176588
rect 269120 176536 269172 176588
rect 300216 176536 300268 176588
rect 306564 176536 306616 176588
rect 255964 176196 256016 176248
rect 262220 176196 262272 176248
rect 300124 176196 300176 176248
rect 301136 176196 301188 176248
rect 130752 175992 130804 176044
rect 165528 175992 165580 176044
rect 187056 175992 187108 176044
rect 204904 175992 204956 176044
rect 123116 175924 123168 175976
rect 249248 175924 249300 175976
rect 298192 175788 298244 175840
rect 249708 175312 249760 175364
rect 264428 175312 264480 175364
rect 143448 175176 143500 175228
rect 249708 175176 249760 175228
rect 185676 175108 185728 175160
rect 264336 175108 264388 175160
rect 301412 175108 301464 175160
rect 283748 174020 283800 174072
rect 287796 174020 287848 174072
rect 276664 173884 276716 173936
rect 288348 173884 288400 173936
rect 165528 173816 165580 173868
rect 248604 173816 248656 173868
rect 266636 173816 266688 173868
rect 280252 173816 280304 173868
rect 231584 173748 231636 173800
rect 249708 173748 249760 173800
rect 266360 173748 266412 173800
rect 271972 173748 272024 173800
rect 287796 173340 287848 173392
rect 287980 173340 288032 173392
rect 282276 172592 282328 172644
rect 287612 172592 287664 172644
rect 273904 172524 273956 172576
rect 288348 172524 288400 172576
rect 168472 172456 168524 172508
rect 248604 172456 248656 172508
rect 266636 172456 266688 172508
rect 273352 172456 273404 172508
rect 303896 172456 303948 172508
rect 316224 172456 316276 172508
rect 233976 172388 234028 172440
rect 249340 172388 249392 172440
rect 266360 172388 266412 172440
rect 269120 172388 269172 172440
rect 280896 171164 280948 171216
rect 288348 171164 288400 171216
rect 278320 171096 278372 171148
rect 288256 171096 288308 171148
rect 166448 171028 166500 171080
rect 249616 171028 249668 171080
rect 266728 171028 266780 171080
rect 280160 171028 280212 171080
rect 169116 170960 169168 171012
rect 249708 170960 249760 171012
rect 266360 170960 266412 171012
rect 270500 170960 270552 171012
rect 279608 169736 279660 169788
rect 288348 169736 288400 169788
rect 164976 169668 165028 169720
rect 249708 169668 249760 169720
rect 266360 169668 266412 169720
rect 270776 169668 270828 169720
rect 303896 169668 303948 169720
rect 311900 169668 311952 169720
rect 217324 168988 217376 169040
rect 249156 168988 249208 169040
rect 266360 168988 266412 169040
rect 269304 168988 269356 169040
rect 269948 168988 270000 169040
rect 287244 168988 287296 169040
rect 271420 168376 271472 168428
rect 288164 168376 288216 168428
rect 167920 168308 167972 168360
rect 249616 168308 249668 168360
rect 303896 168308 303948 168360
rect 320456 168308 320508 168360
rect 185768 168240 185820 168292
rect 249708 168240 249760 168292
rect 266360 167968 266412 168020
rect 268016 167968 268068 168020
rect 268660 167084 268712 167136
rect 276020 167084 276072 167136
rect 280804 167084 280856 167136
rect 287980 167084 288032 167136
rect 272616 167016 272668 167068
rect 288348 167016 288400 167068
rect 164884 166948 164936 167000
rect 248420 166948 248472 167000
rect 303896 166948 303948 167000
rect 310796 166948 310848 167000
rect 522304 166948 522356 167000
rect 580172 166948 580224 167000
rect 184388 166880 184440 166932
rect 248512 166880 248564 166932
rect 266360 166336 266412 166388
rect 269396 166336 269448 166388
rect 268568 166268 268620 166320
rect 287888 166268 287940 166320
rect 304264 166268 304316 166320
rect 323216 166268 323268 166320
rect 283656 165588 283708 165640
rect 288348 165588 288400 165640
rect 173440 165520 173492 165572
rect 248420 165520 248472 165572
rect 264152 165520 264204 165572
rect 264980 165520 265032 165572
rect 266360 165520 266412 165572
rect 272064 165520 272116 165572
rect 303896 165520 303948 165572
rect 309416 165520 309468 165572
rect 278136 165112 278188 165164
rect 281632 165112 281684 165164
rect 271328 164840 271380 164892
rect 288256 164840 288308 164892
rect 282552 164432 282604 164484
rect 288716 164432 288768 164484
rect 3240 164160 3292 164212
rect 33784 164160 33836 164212
rect 182916 164160 182968 164212
rect 248512 164160 248564 164212
rect 266360 164160 266412 164212
rect 277400 164160 277452 164212
rect 303896 164160 303948 164212
rect 325884 164160 325936 164212
rect 231216 164092 231268 164144
rect 248420 164092 248472 164144
rect 271236 164092 271288 164144
rect 273352 164092 273404 164144
rect 170404 163480 170456 163532
rect 221464 163480 221516 163532
rect 303896 163276 303948 163328
rect 307944 163276 307996 163328
rect 276756 162868 276808 162920
rect 288164 162868 288216 162920
rect 171876 162800 171928 162852
rect 248420 162800 248472 162852
rect 266544 162800 266596 162852
rect 270592 162800 270644 162852
rect 303896 162800 303948 162852
rect 317604 162800 317656 162852
rect 181444 162732 181496 162784
rect 248512 162732 248564 162784
rect 266360 162528 266412 162580
rect 269212 162528 269264 162580
rect 269212 162120 269264 162172
rect 283104 162120 283156 162172
rect 282460 161508 282512 161560
rect 288256 161508 288308 161560
rect 285128 161440 285180 161492
rect 288348 161440 288400 161492
rect 167736 161372 167788 161424
rect 248512 161372 248564 161424
rect 266360 161372 266412 161424
rect 274824 161372 274876 161424
rect 303896 161372 303948 161424
rect 319076 161372 319128 161424
rect 238024 161304 238076 161356
rect 248420 161304 248472 161356
rect 269764 160080 269816 160132
rect 287520 160080 287572 160132
rect 177488 160012 177540 160064
rect 248420 160012 248472 160064
rect 303804 159876 303856 159928
rect 306564 159876 306616 159928
rect 265072 159332 265124 159384
rect 271880 159332 271932 159384
rect 281080 158788 281132 158840
rect 288348 158788 288400 158840
rect 279424 158720 279476 158772
rect 287428 158720 287480 158772
rect 170496 158652 170548 158704
rect 248420 158652 248472 158704
rect 266360 158652 266412 158704
rect 274640 158652 274692 158704
rect 303620 158652 303672 158704
rect 310704 158652 310756 158704
rect 275376 158244 275428 158296
rect 279608 158244 279660 158296
rect 178868 157972 178920 158024
rect 249432 157972 249484 158024
rect 266728 157972 266780 158024
rect 276112 157972 276164 158024
rect 277032 157972 277084 158024
rect 280896 157972 280948 158024
rect 283840 157904 283892 157956
rect 287152 157904 287204 157956
rect 176016 157292 176068 157344
rect 249616 157292 249668 157344
rect 266360 157292 266412 157344
rect 270592 157292 270644 157344
rect 303804 157292 303856 157344
rect 313556 157292 313608 157344
rect 188436 157224 188488 157276
rect 249708 157224 249760 157276
rect 283564 156000 283616 156052
rect 288348 156000 288400 156052
rect 279608 155932 279660 155984
rect 288164 155932 288216 155984
rect 166356 155864 166408 155916
rect 249708 155864 249760 155916
rect 266360 155864 266412 155916
rect 280344 155864 280396 155916
rect 303620 155864 303672 155916
rect 331312 155864 331364 155916
rect 220084 155796 220136 155848
rect 249616 155796 249668 155848
rect 303804 155796 303856 155848
rect 321744 155796 321796 155848
rect 266360 155320 266412 155372
rect 270040 155320 270092 155372
rect 177396 155184 177448 155236
rect 213184 155184 213236 155236
rect 287704 155184 287756 155236
rect 288532 155184 288584 155236
rect 281172 155116 281224 155168
rect 287980 155116 288032 155168
rect 269856 154572 269908 154624
rect 288348 154572 288400 154624
rect 303804 154504 303856 154556
rect 335544 154504 335596 154556
rect 303620 154436 303672 154488
rect 332692 154436 332744 154488
rect 265716 153892 265768 153944
rect 283656 153892 283708 153944
rect 268476 153824 268528 153876
rect 287888 153824 287940 153876
rect 266360 153348 266412 153400
rect 268660 153348 268712 153400
rect 246396 153280 246448 153332
rect 249708 153280 249760 153332
rect 214564 153212 214616 153264
rect 249156 153212 249208 153264
rect 303804 153144 303856 153196
rect 324504 153144 324556 153196
rect 303896 153076 303948 153128
rect 312084 153076 312136 153128
rect 174636 152464 174688 152516
rect 217324 152464 217376 152516
rect 267096 152464 267148 152516
rect 282276 152464 282328 152516
rect 222936 151852 222988 151904
rect 249708 151852 249760 151904
rect 283656 151852 283708 151904
rect 288348 151852 288400 151904
rect 214656 151784 214708 151836
rect 248972 151784 249024 151836
rect 266268 151784 266320 151836
rect 288256 151784 288308 151836
rect 266360 151580 266412 151632
rect 269120 151580 269172 151632
rect 169024 151036 169076 151088
rect 248972 151036 249024 151088
rect 278136 150492 278188 150544
rect 288348 150492 288400 150544
rect 178868 150424 178920 150476
rect 249708 150424 249760 150476
rect 275468 150424 275520 150476
rect 287980 150424 288032 150476
rect 3516 150356 3568 150408
rect 14464 150356 14516 150408
rect 167644 150356 167696 150408
rect 249616 150356 249668 150408
rect 266360 150356 266412 150408
rect 278780 150356 278832 150408
rect 303804 150356 303856 150408
rect 316316 150356 316368 150408
rect 180156 149676 180208 149728
rect 249248 149676 249300 149728
rect 280988 149064 281040 149116
rect 288348 149064 288400 149116
rect 303804 148996 303856 149048
rect 320272 148996 320324 149048
rect 267188 148384 267240 148436
rect 279516 148384 279568 148436
rect 181536 148316 181588 148368
rect 226984 148316 227036 148368
rect 270040 148316 270092 148368
rect 284944 148316 284996 148368
rect 279700 147636 279752 147688
rect 288348 147636 288400 147688
rect 266360 147568 266412 147620
rect 275560 147568 275612 147620
rect 303712 147568 303764 147620
rect 327356 147568 327408 147620
rect 276940 146888 276992 146940
rect 287244 146888 287296 146940
rect 246488 146344 246540 146396
rect 249708 146344 249760 146396
rect 177396 146276 177448 146328
rect 249156 146276 249208 146328
rect 264244 146276 264296 146328
rect 288348 146276 288400 146328
rect 303804 146208 303856 146260
rect 317696 146208 317748 146260
rect 303712 145800 303764 145852
rect 308036 145800 308088 145852
rect 274088 145664 274140 145716
rect 277032 145664 277084 145716
rect 198004 145596 198056 145648
rect 218796 145596 218848 145648
rect 171784 145528 171836 145580
rect 204996 145528 205048 145580
rect 231216 144916 231268 144968
rect 249708 144916 249760 144968
rect 284944 144916 284996 144968
rect 287428 144916 287480 144968
rect 266360 144848 266412 144900
rect 271236 144848 271288 144900
rect 303804 144848 303856 144900
rect 323124 144848 323176 144900
rect 275560 144168 275612 144220
rect 287796 144168 287848 144220
rect 303988 144168 304040 144220
rect 316132 144168 316184 144220
rect 238024 143624 238076 143676
rect 249708 143624 249760 143676
rect 196716 143556 196768 143608
rect 249156 143556 249208 143608
rect 265624 143556 265676 143608
rect 288164 143556 288216 143608
rect 266360 143488 266412 143540
rect 273260 143488 273312 143540
rect 175924 142808 175976 142860
rect 249616 142808 249668 142860
rect 274180 142808 274232 142860
rect 287888 142808 287940 142860
rect 242256 142128 242308 142180
rect 249708 142128 249760 142180
rect 272800 142128 272852 142180
rect 279608 142128 279660 142180
rect 282368 142128 282420 142180
rect 287980 142128 288032 142180
rect 303804 142060 303856 142112
rect 322940 142060 322992 142112
rect 191104 141448 191156 141500
rect 209044 141448 209096 141500
rect 271236 141448 271288 141500
rect 288256 141448 288308 141500
rect 178776 141380 178828 141432
rect 199384 141380 199436 141432
rect 266452 141380 266504 141432
rect 285220 141380 285272 141432
rect 229836 140836 229888 140888
rect 249616 140836 249668 140888
rect 224224 140768 224276 140820
rect 249708 140768 249760 140820
rect 284300 139816 284352 139868
rect 288072 139816 288124 139868
rect 303620 139816 303672 139868
rect 305276 139816 305328 139868
rect 232688 139408 232740 139460
rect 249156 139408 249208 139460
rect 266360 139340 266412 139392
rect 267740 139340 267792 139392
rect 303804 139340 303856 139392
rect 314844 139340 314896 139392
rect 264060 138864 264112 138916
rect 173256 138660 173308 138712
rect 198096 138660 198148 138712
rect 233976 138660 234028 138712
rect 249340 138660 249392 138712
rect 280804 138660 280856 138712
rect 280896 138048 280948 138100
rect 288256 138048 288308 138100
rect 181444 137980 181496 138032
rect 249708 137980 249760 138032
rect 268660 137980 268712 138032
rect 269948 137980 270000 138032
rect 279608 137980 279660 138032
rect 288348 137980 288400 138032
rect 3516 137912 3568 137964
rect 25504 137912 25556 137964
rect 303804 137912 303856 137964
rect 328552 137912 328604 137964
rect 186964 137300 187016 137352
rect 202144 137300 202196 137352
rect 277124 137300 277176 137352
rect 281172 137300 281224 137352
rect 167736 137232 167788 137284
rect 222936 137232 222988 137284
rect 266360 137232 266412 137284
rect 283748 137232 283800 137284
rect 245016 136688 245068 136740
rect 249156 136688 249208 136740
rect 203616 136620 203668 136672
rect 249708 136620 249760 136672
rect 283840 136620 283892 136672
rect 288348 136620 288400 136672
rect 303620 136552 303672 136604
rect 310612 136552 310664 136604
rect 195336 135872 195388 135924
rect 220084 135872 220136 135924
rect 268752 135872 268804 135924
rect 289176 135872 289228 135924
rect 266360 135600 266412 135652
rect 268568 135600 268620 135652
rect 235264 135328 235316 135380
rect 249708 135328 249760 135380
rect 167644 135260 167696 135312
rect 249156 135260 249208 135312
rect 266360 135192 266412 135244
rect 276664 135192 276716 135244
rect 303712 135192 303764 135244
rect 339592 135192 339644 135244
rect 198004 134512 198056 134564
rect 246488 134512 246540 134564
rect 304724 134512 304776 134564
rect 312176 134512 312228 134564
rect 171784 133900 171836 133952
rect 249708 133900 249760 133952
rect 266360 133832 266412 133884
rect 273904 133832 273956 133884
rect 303896 133832 303948 133884
rect 331404 133832 331456 133884
rect 303804 133764 303856 133816
rect 321652 133764 321704 133816
rect 274272 133220 274324 133272
rect 287428 133220 287480 133272
rect 173348 133152 173400 133204
rect 249248 133152 249300 133204
rect 269948 133152 270000 133204
rect 284300 133152 284352 133204
rect 266360 132948 266412 133000
rect 268660 132948 268712 133000
rect 285220 132472 285272 132524
rect 288348 132472 288400 132524
rect 266452 132404 266504 132456
rect 275376 132404 275428 132456
rect 303804 132404 303856 132456
rect 327172 132404 327224 132456
rect 266360 132336 266412 132388
rect 274088 132336 274140 132388
rect 303896 132336 303948 132388
rect 317512 132336 317564 132388
rect 176016 131724 176068 131776
rect 246396 131724 246448 131776
rect 173256 131112 173308 131164
rect 249708 131112 249760 131164
rect 274548 131112 274600 131164
rect 288348 131112 288400 131164
rect 266452 131044 266504 131096
rect 271420 131044 271472 131096
rect 303804 131044 303856 131096
rect 329932 131044 329984 131096
rect 266544 130908 266596 130960
rect 270040 130908 270092 130960
rect 278320 130364 278372 130416
rect 289268 130364 289320 130416
rect 304264 130364 304316 130416
rect 318984 130364 319036 130416
rect 213276 129820 213328 129872
rect 249616 129820 249668 129872
rect 211896 129752 211948 129804
rect 249708 129752 249760 129804
rect 277032 129752 277084 129804
rect 288348 129752 288400 129804
rect 266360 129684 266412 129736
rect 276848 129684 276900 129736
rect 303804 129684 303856 129736
rect 314936 129684 314988 129736
rect 267096 129616 267148 129668
rect 269764 129616 269816 129668
rect 270040 129004 270092 129056
rect 287704 129004 287756 129056
rect 195336 128324 195388 128376
rect 249708 128324 249760 128376
rect 276756 128324 276808 128376
rect 287980 128324 288032 128376
rect 303804 128256 303856 128308
rect 336740 128256 336792 128308
rect 303620 128188 303672 128240
rect 313372 128188 313424 128240
rect 266360 127984 266412 128036
rect 268752 127984 268804 128036
rect 264796 127644 264848 127696
rect 267004 127644 267056 127696
rect 266452 127576 266504 127628
rect 273996 127576 274048 127628
rect 268568 127440 268620 127492
rect 272800 127440 272852 127492
rect 229744 127032 229796 127084
rect 249708 127032 249760 127084
rect 188528 126964 188580 127016
rect 249616 126964 249668 127016
rect 283932 126964 283984 127016
rect 287980 126964 288032 127016
rect 266360 126896 266412 126948
rect 271328 126896 271380 126948
rect 184296 126284 184348 126336
rect 196624 126284 196676 126336
rect 178776 126216 178828 126268
rect 214656 126216 214708 126268
rect 267004 126216 267056 126268
rect 277124 126216 277176 126268
rect 220176 125672 220228 125724
rect 249616 125672 249668 125724
rect 280804 125672 280856 125724
rect 288256 125672 288308 125724
rect 200856 125604 200908 125656
rect 249708 125604 249760 125656
rect 272708 125604 272760 125656
rect 288348 125604 288400 125656
rect 266360 125536 266412 125588
rect 275284 125536 275336 125588
rect 303712 125536 303764 125588
rect 328460 125536 328512 125588
rect 202328 124924 202380 124976
rect 228456 124924 228508 124976
rect 184388 124856 184440 124908
rect 232688 124856 232740 124908
rect 266912 124856 266964 124908
rect 285128 124856 285180 124908
rect 238116 124244 238168 124296
rect 249616 124244 249668 124296
rect 232596 124176 232648 124228
rect 249708 124176 249760 124228
rect 282828 124176 282880 124228
rect 288348 124176 288400 124228
rect 303712 124108 303764 124160
rect 327264 124108 327316 124160
rect 303804 124040 303856 124092
rect 325700 124040 325752 124092
rect 164884 123428 164936 123480
rect 231308 123428 231360 123480
rect 272800 123428 272852 123480
rect 287888 123428 287940 123480
rect 266360 123156 266412 123208
rect 268476 123156 268528 123208
rect 243728 122884 243780 122936
rect 249524 122884 249576 122936
rect 185676 122816 185728 122868
rect 248972 122816 249024 122868
rect 275284 122816 275336 122868
rect 287980 122816 288032 122868
rect 266544 122748 266596 122800
rect 286324 122748 286376 122800
rect 303620 122748 303672 122800
rect 324412 122748 324464 122800
rect 266360 122680 266412 122732
rect 282460 122680 282512 122732
rect 191196 122068 191248 122120
rect 238024 122068 238076 122120
rect 239404 121524 239456 121576
rect 248788 121524 248840 121576
rect 166264 121456 166316 121508
rect 249708 121456 249760 121508
rect 283748 121456 283800 121508
rect 288256 121456 288308 121508
rect 303804 121388 303856 121440
rect 320364 121388 320416 121440
rect 222844 120708 222896 120760
rect 236736 120708 236788 120760
rect 269764 120708 269816 120760
rect 287152 120708 287204 120760
rect 238024 120164 238076 120216
rect 249708 120164 249760 120216
rect 264244 120164 264296 120216
rect 225604 120096 225656 120148
rect 249616 120096 249668 120148
rect 264796 120096 264848 120148
rect 266636 120096 266688 120148
rect 288256 120096 288308 120148
rect 266544 120028 266596 120080
rect 286508 120028 286560 120080
rect 303804 120028 303856 120080
rect 318892 120028 318944 120080
rect 266360 119960 266412 120012
rect 281080 119960 281132 120012
rect 184296 118736 184348 118788
rect 249708 118736 249760 118788
rect 182916 118668 182968 118720
rect 248788 118668 248840 118720
rect 285128 118668 285180 118720
rect 287612 118668 287664 118720
rect 266360 118600 266412 118652
rect 279424 118600 279476 118652
rect 303896 118600 303948 118652
rect 311992 118600 312044 118652
rect 266544 118532 266596 118584
rect 274180 118532 274232 118584
rect 303804 118396 303856 118448
rect 307852 118396 307904 118448
rect 186964 117920 187016 117972
rect 249616 117920 249668 117972
rect 278504 117444 278556 117496
rect 282828 117444 282880 117496
rect 236000 117308 236052 117360
rect 248788 117308 248840 117360
rect 279516 117308 279568 117360
rect 288256 117308 288308 117360
rect 266360 117240 266412 117292
rect 272524 117240 272576 117292
rect 303804 117240 303856 117292
rect 314660 117240 314712 117292
rect 266268 117172 266320 117224
rect 266636 117172 266688 117224
rect 170680 116560 170732 116612
rect 236000 116560 236052 116612
rect 269028 116560 269080 116612
rect 285220 116560 285272 116612
rect 266360 116152 266412 116204
rect 268568 116152 268620 116204
rect 285588 116016 285640 116068
rect 287428 116016 287480 116068
rect 224316 115948 224368 116000
rect 248788 115948 248840 116000
rect 272616 115948 272668 116000
rect 288164 115948 288216 116000
rect 266544 115880 266596 115932
rect 285036 115880 285088 115932
rect 303804 115880 303856 115932
rect 310520 115880 310572 115932
rect 266360 115812 266412 115864
rect 271144 115812 271196 115864
rect 303620 115404 303672 115456
rect 306472 115404 306524 115456
rect 238208 114520 238260 114572
rect 249708 114520 249760 114572
rect 285220 114520 285272 114572
rect 288256 114520 288308 114572
rect 266544 114452 266596 114504
rect 275560 114452 275612 114504
rect 303804 114452 303856 114504
rect 316040 114452 316092 114504
rect 273168 113772 273220 113824
rect 282460 113772 282512 113824
rect 266360 113636 266412 113688
rect 269856 113636 269908 113688
rect 173440 113228 173492 113280
rect 230480 113228 230532 113280
rect 235356 113228 235408 113280
rect 249708 113228 249760 113280
rect 284024 113228 284076 113280
rect 287980 113228 288032 113280
rect 167828 113160 167880 113212
rect 249616 113160 249668 113212
rect 275376 113160 275428 113212
rect 287612 113160 287664 113212
rect 230480 113092 230532 113144
rect 243728 113092 243780 113144
rect 266544 113092 266596 113144
rect 289084 113092 289136 113144
rect 303804 113092 303856 113144
rect 307760 113092 307812 113144
rect 266360 113024 266412 113076
rect 278228 113024 278280 113076
rect 303712 112752 303764 112804
rect 306656 112752 306708 112804
rect 174636 112412 174688 112464
rect 224224 112412 224276 112464
rect 243636 111868 243688 111920
rect 248972 111868 249024 111920
rect 244924 111800 244976 111852
rect 249248 111800 249300 111852
rect 278412 111800 278464 111852
rect 285128 111800 285180 111852
rect 168288 111732 168340 111784
rect 178868 111732 178920 111784
rect 303712 111732 303764 111784
rect 325792 111732 325844 111784
rect 303804 111664 303856 111716
rect 313280 111664 313332 111716
rect 267004 111120 267056 111172
rect 272616 111120 272668 111172
rect 268476 111052 268528 111104
rect 278504 111052 278556 111104
rect 180340 110508 180392 110560
rect 248972 110508 249024 110560
rect 282920 110508 282972 110560
rect 287980 110508 288032 110560
rect 172060 110440 172112 110492
rect 249248 110440 249300 110492
rect 278044 110440 278096 110492
rect 288256 110440 288308 110492
rect 167920 110372 167972 110424
rect 180156 110372 180208 110424
rect 266452 110372 266504 110424
rect 278136 110372 278188 110424
rect 266360 110304 266412 110356
rect 275468 110304 275520 110356
rect 211804 109080 211856 109132
rect 249708 109080 249760 109132
rect 283564 109080 283616 109132
rect 288256 109080 288308 109132
rect 180248 109012 180300 109064
rect 249616 109012 249668 109064
rect 278228 109012 278280 109064
rect 288348 109012 288400 109064
rect 266360 108944 266412 108996
rect 280988 108944 281040 108996
rect 303804 108944 303856 108996
rect 321560 108944 321612 108996
rect 170404 108264 170456 108316
rect 229836 108264 229888 108316
rect 234160 107720 234212 107772
rect 249708 107720 249760 107772
rect 231308 107652 231360 107704
rect 249524 107652 249576 107704
rect 267188 107652 267240 107704
rect 288348 107652 288400 107704
rect 266360 107584 266412 107636
rect 279700 107584 279752 107636
rect 303804 107584 303856 107636
rect 309140 107584 309192 107636
rect 266452 107516 266504 107568
rect 276940 107516 276992 107568
rect 285128 106428 285180 106480
rect 287980 106428 288032 106480
rect 191288 106360 191340 106412
rect 249708 106360 249760 106412
rect 280988 106360 281040 106412
rect 288348 106360 288400 106412
rect 166356 106292 166408 106344
rect 249524 106292 249576 106344
rect 266360 106224 266412 106276
rect 282276 106224 282328 106276
rect 200764 104932 200816 104984
rect 249708 104932 249760 104984
rect 281080 104932 281132 104984
rect 287980 104932 288032 104984
rect 167736 104864 167788 104916
rect 248788 104864 248840 104916
rect 283840 104864 283892 104916
rect 288348 104864 288400 104916
rect 303804 104796 303856 104848
rect 314752 104796 314804 104848
rect 272892 104184 272944 104236
rect 282920 104184 282972 104236
rect 169116 104116 169168 104168
rect 211896 104116 211948 104168
rect 264428 104116 264480 104168
rect 283748 104116 283800 104168
rect 266360 104048 266412 104100
rect 269948 104048 270000 104100
rect 171968 103504 172020 103556
rect 249708 103504 249760 103556
rect 266452 103436 266504 103488
rect 284944 103436 284996 103488
rect 266360 103368 266412 103420
rect 271236 103368 271288 103420
rect 281540 102280 281592 102332
rect 285220 102280 285272 102332
rect 278136 102212 278188 102264
rect 282460 102212 282512 102264
rect 285036 102212 285088 102264
rect 288348 102212 288400 102264
rect 174728 102144 174780 102196
rect 249708 102144 249760 102196
rect 271512 102144 271564 102196
rect 278412 102144 278464 102196
rect 284300 102144 284352 102196
rect 288256 102144 288308 102196
rect 303712 102076 303764 102128
rect 323032 102076 323084 102128
rect 266360 102008 266412 102060
rect 270040 102008 270092 102060
rect 166448 101396 166500 101448
rect 200856 101396 200908 101448
rect 218796 101396 218848 101448
rect 251824 101396 251876 101448
rect 284944 100784 284996 100836
rect 287612 100784 287664 100836
rect 177488 100716 177540 100768
rect 249156 100716 249208 100768
rect 265624 100716 265676 100768
rect 272064 100716 272116 100768
rect 279700 100716 279752 100768
rect 288348 100716 288400 100768
rect 266360 100648 266412 100700
rect 282368 100648 282420 100700
rect 266452 100580 266504 100632
rect 272800 100580 272852 100632
rect 164976 99968 165028 100020
rect 249064 99968 249116 100020
rect 284116 99424 284168 99476
rect 288256 99424 288308 99476
rect 214656 99356 214708 99408
rect 249708 99356 249760 99408
rect 272616 99356 272668 99408
rect 288348 99356 288400 99408
rect 266452 99288 266504 99340
rect 274272 99288 274324 99340
rect 276940 98676 276992 98728
rect 282920 98676 282972 98728
rect 273904 98608 273956 98660
rect 281540 98608 281592 98660
rect 283656 98132 283708 98184
rect 287888 98132 287940 98184
rect 203524 98064 203576 98116
rect 249708 98064 249760 98116
rect 282368 98064 282420 98116
rect 286784 98064 286836 98116
rect 171876 97996 171928 98048
rect 249616 97996 249668 98048
rect 264060 97996 264112 98048
rect 268292 97996 268344 98048
rect 3424 97928 3476 97980
rect 21364 97928 21416 97980
rect 210424 97928 210476 97980
rect 252192 97928 252244 97980
rect 265808 97724 265860 97776
rect 267280 97724 267332 97776
rect 178868 97248 178920 97300
rect 209228 97248 209280 97300
rect 165528 96636 165580 96688
rect 249708 96636 249760 96688
rect 252192 96636 252244 96688
rect 264060 96772 264112 96824
rect 288348 97248 288400 97300
rect 257804 96024 257856 96076
rect 257896 96024 257948 96076
rect 303896 96568 303948 96620
rect 334072 96568 334124 96620
rect 261024 96024 261076 96076
rect 165620 95956 165672 96008
rect 214564 95956 214616 96008
rect 224868 95956 224920 96008
rect 290924 95956 290976 96008
rect 168656 95888 168708 95940
rect 247868 95888 247920 95940
rect 258724 95888 258776 95940
rect 266268 95888 266320 95940
rect 271144 95208 271196 95260
rect 278320 95208 278372 95260
rect 246396 95140 246448 95192
rect 301504 95140 301556 95192
rect 289728 95072 289780 95124
rect 291292 95072 291344 95124
rect 67732 94460 67784 94512
rect 100024 94460 100076 94512
rect 181536 94460 181588 94512
rect 248788 94460 248840 94512
rect 257344 94460 257396 94512
rect 264152 94460 264204 94512
rect 162860 94392 162912 94444
rect 165620 94392 165672 94444
rect 124036 93848 124088 93900
rect 238116 93848 238168 93900
rect 267740 93780 267792 93832
rect 295984 93780 296036 93832
rect 290924 93712 290976 93764
rect 303804 93712 303856 93764
rect 67364 93168 67416 93220
rect 88984 93168 89036 93220
rect 119712 93168 119764 93220
rect 166264 93168 166316 93220
rect 170588 93168 170640 93220
rect 177580 93168 177632 93220
rect 184388 93168 184440 93220
rect 206376 93168 206428 93220
rect 246304 93168 246356 93220
rect 265900 93168 265952 93220
rect 66076 93100 66128 93152
rect 106188 93100 106240 93152
rect 121736 93100 121788 93152
rect 185676 93100 185728 93152
rect 260104 93100 260156 93152
rect 283840 93100 283892 93152
rect 136088 92420 136140 92472
rect 173348 92420 173400 92472
rect 250720 92420 250772 92472
rect 303620 92420 303672 92472
rect 151360 92352 151412 92404
rect 162860 92352 162912 92404
rect 117228 91740 117280 91792
rect 126888 91740 126940 91792
rect 164148 91740 164200 91792
rect 235264 91740 235316 91792
rect 235908 91740 235960 91792
rect 266452 91740 266504 91792
rect 267096 91740 267148 91792
rect 274640 91740 274692 91792
rect 86868 91128 86920 91180
rect 106924 91128 106976 91180
rect 114468 91128 114520 91180
rect 134708 91128 134760 91180
rect 89076 91060 89128 91112
rect 116584 91060 116636 91112
rect 127992 91060 128044 91112
rect 129004 91060 129056 91112
rect 109960 90992 110012 91044
rect 224316 90992 224368 91044
rect 236736 90992 236788 91044
rect 303712 90992 303764 91044
rect 111616 90924 111668 90976
rect 170680 90924 170732 90976
rect 65984 90312 66036 90364
rect 111064 90312 111116 90364
rect 175924 90312 175976 90364
rect 196716 90312 196768 90364
rect 198096 90312 198148 90364
rect 286508 90312 286560 90364
rect 122840 89632 122892 89684
rect 232596 89632 232648 89684
rect 251824 89632 251876 89684
rect 301136 89632 301188 89684
rect 107476 89564 107528 89616
rect 158720 89564 158772 89616
rect 98736 88952 98788 89004
rect 122196 88952 122248 89004
rect 160100 88952 160152 89004
rect 176016 88952 176068 89004
rect 196716 88952 196768 89004
rect 264428 88952 264480 89004
rect 102600 88272 102652 88324
rect 235356 88272 235408 88324
rect 134708 88204 134760 88256
rect 164148 88204 164200 88256
rect 164976 87592 165028 87644
rect 243636 87592 243688 87644
rect 260196 87592 260248 87644
rect 272892 87592 272944 87644
rect 75920 86912 75972 86964
rect 249340 86912 249392 86964
rect 113456 86844 113508 86896
rect 182916 86844 182968 86896
rect 253204 86300 253256 86352
rect 270132 86300 270184 86352
rect 66168 86232 66220 86284
rect 107016 86232 107068 86284
rect 191104 86232 191156 86284
rect 278136 86232 278188 86284
rect 3148 85484 3200 85536
rect 29644 85484 29696 85536
rect 125416 85484 125468 85536
rect 166448 85484 166500 85536
rect 151636 85416 151688 85468
rect 160100 85416 160152 85468
rect 206284 84872 206336 84924
rect 275560 84872 275612 84924
rect 160744 84804 160796 84856
rect 263048 84804 263100 84856
rect 95056 84124 95108 84176
rect 231308 84124 231360 84176
rect 97908 84056 97960 84108
rect 180248 84056 180300 84108
rect 255964 83512 256016 83564
rect 276940 83512 276992 83564
rect 221464 83444 221516 83496
rect 295984 83444 296036 83496
rect 96528 82764 96580 82816
rect 211804 82764 211856 82816
rect 114284 82696 114336 82748
rect 167644 82696 167696 82748
rect 95148 81336 95200 81388
rect 234160 81336 234212 81388
rect 151084 81268 151136 81320
rect 162216 81268 162268 81320
rect 162124 80656 162176 80708
rect 264336 80656 264388 80708
rect 122196 79976 122248 80028
rect 163504 79976 163556 80028
rect 151728 79908 151780 79960
rect 178776 79908 178828 79960
rect 88984 78616 89036 78668
rect 200764 78616 200816 78668
rect 324964 78616 325016 78668
rect 325700 78616 325752 78668
rect 125508 78548 125560 78600
rect 170404 78548 170456 78600
rect 229744 77936 229796 77988
rect 275284 77936 275336 77988
rect 91008 77188 91060 77240
rect 167736 77188 167788 77240
rect 118516 77120 118568 77172
rect 181444 77120 181496 77172
rect 121368 75828 121420 75880
rect 173440 75828 173492 75880
rect 97908 75148 97960 75200
rect 278228 75148 278280 75200
rect 116584 74468 116636 74520
rect 214656 74468 214708 74520
rect 153108 74400 153160 74452
rect 233976 74400 234028 74452
rect 86776 73788 86828 73840
rect 105544 73788 105596 73840
rect 100024 73108 100076 73160
rect 209136 73108 209188 73160
rect 124128 73040 124180 73092
rect 174636 73040 174688 73092
rect 3424 71680 3476 71732
rect 18604 71680 18656 71732
rect 119988 71680 120040 71732
rect 177396 71680 177448 71732
rect 113088 71000 113140 71052
rect 274088 71000 274140 71052
rect 129648 70320 129700 70372
rect 175924 70320 175976 70372
rect 119988 69640 120040 69692
rect 272708 69640 272760 69692
rect 108856 68960 108908 69012
rect 184388 68960 184440 69012
rect 133788 68892 133840 68944
rect 198004 68892 198056 68944
rect 110328 67532 110380 67584
rect 170588 67532 170640 67584
rect 71044 66852 71096 66904
rect 245016 66852 245068 66904
rect 112996 66172 113048 66224
rect 186964 66172 187016 66224
rect 106924 66104 106976 66156
rect 171876 66104 171928 66156
rect 251824 65492 251876 65544
rect 268660 65492 268712 65544
rect 88156 64812 88208 64864
rect 199476 64812 199528 64864
rect 103428 64744 103480 64796
rect 213276 64744 213328 64796
rect 126704 63452 126756 63504
rect 220176 63452 220228 63504
rect 104808 63384 104860 63436
rect 178868 63384 178920 63436
rect 115848 62024 115900 62076
rect 238024 62024 238076 62076
rect 59176 61344 59228 61396
rect 274180 61344 274232 61396
rect 105544 60664 105596 60716
rect 203524 60664 203576 60716
rect 129004 60596 129056 60648
rect 191196 60596 191248 60648
rect 3056 59304 3108 59356
rect 17224 59304 17276 59356
rect 108948 59304 109000 59356
rect 202328 59304 202380 59356
rect 126796 59236 126848 59288
rect 188436 59236 188488 59288
rect 214656 58624 214708 58676
rect 236000 58624 236052 58676
rect 101956 57876 102008 57928
rect 195336 57876 195388 57928
rect 77208 57196 77260 57248
rect 280988 57196 281040 57248
rect 126888 56516 126940 56568
rect 242256 56516 242308 56568
rect 91008 55836 91060 55888
rect 267188 55836 267240 55888
rect 102048 55156 102100 55208
rect 244924 55156 244976 55208
rect 95056 54476 95108 54528
rect 286324 54476 286376 54528
rect 118608 53728 118660 53780
rect 239404 53728 239456 53780
rect 102048 53048 102100 53100
rect 273996 53048 274048 53100
rect 117228 52368 117280 52420
rect 225604 52368 225656 52420
rect 104808 51688 104860 51740
rect 283564 51688 283616 51740
rect 174544 50396 174596 50448
rect 273260 50396 273312 50448
rect 86868 50328 86920 50380
rect 289084 50328 289136 50380
rect 107568 49036 107620 49088
rect 250536 49036 250588 49088
rect 37188 48968 37240 49020
rect 276756 48968 276808 49020
rect 71688 47608 71740 47660
rect 265808 47608 265860 47660
rect 39948 47540 40000 47592
rect 236644 47540 236696 47592
rect 238024 47540 238076 47592
rect 249064 47540 249116 47592
rect 119896 46248 119948 46300
rect 268568 46248 268620 46300
rect 126244 46180 126296 46232
rect 282368 46180 282420 46232
rect 2780 45500 2832 45552
rect 4804 45500 4856 45552
rect 115848 44820 115900 44872
rect 260196 44820 260248 44872
rect 84108 43460 84160 43512
rect 271328 43460 271380 43512
rect 75828 43392 75880 43444
rect 283656 43392 283708 43444
rect 12256 42100 12308 42152
rect 272616 42100 272668 42152
rect 5448 42032 5500 42084
rect 291200 42032 291252 42084
rect 205088 40740 205140 40792
rect 214656 40740 214708 40792
rect 217324 40740 217376 40792
rect 291200 40740 291252 40792
rect 57244 40672 57296 40724
rect 253204 40672 253256 40724
rect 74448 39380 74500 39432
rect 160744 39380 160796 39432
rect 213184 39380 213236 39432
rect 276020 39380 276072 39432
rect 146944 39312 146996 39364
rect 260104 39312 260156 39364
rect 55036 37884 55088 37936
rect 282276 37884 282328 37936
rect 79324 36592 79376 36644
rect 251824 36592 251876 36644
rect 3976 36524 4028 36576
rect 262864 36524 262916 36576
rect 204904 35232 204956 35284
rect 287060 35232 287112 35284
rect 1400 35164 1452 35216
rect 229836 35164 229888 35216
rect 142804 33804 142856 33856
rect 206284 33804 206336 33856
rect 41328 33736 41380 33788
rect 147036 33736 147088 33788
rect 199384 33736 199436 33788
rect 269120 33736 269172 33788
rect 3516 33056 3568 33108
rect 39304 33056 39356 33108
rect 189724 32444 189776 32496
rect 271328 32444 271380 32496
rect 124128 32376 124180 32428
rect 280804 32376 280856 32428
rect 196624 31084 196676 31136
rect 259460 31084 259512 31136
rect 118608 31016 118660 31068
rect 232596 31016 232648 31068
rect 122748 29656 122800 29708
rect 198096 29656 198148 29708
rect 185584 29588 185636 29640
rect 267740 29588 267792 29640
rect 130384 28296 130436 28348
rect 168380 28296 168432 28348
rect 182824 28296 182876 28348
rect 271420 28296 271472 28348
rect 53656 28228 53708 28280
rect 279516 28228 279568 28280
rect 114560 26936 114612 26988
rect 205088 26936 205140 26988
rect 44088 26868 44140 26920
rect 151084 26868 151136 26920
rect 204996 26868 205048 26920
rect 263600 26868 263652 26920
rect 209044 25576 209096 25628
rect 295340 25576 295392 25628
rect 96528 25508 96580 25560
rect 271236 25508 271288 25560
rect 117228 24148 117280 24200
rect 268476 24148 268528 24200
rect 81348 24080 81400 24132
rect 264244 24080 264296 24132
rect 111616 22788 111668 22840
rect 278044 22788 278096 22840
rect 56508 22720 56560 22772
rect 276664 22720 276716 22772
rect 125508 21428 125560 21480
rect 267096 21428 267148 21480
rect 50988 21360 51040 21412
rect 251272 21360 251324 21412
rect 3424 20612 3476 20664
rect 36544 20612 36596 20664
rect 112444 20136 112496 20188
rect 114560 20136 114612 20188
rect 188344 20000 188396 20052
rect 242900 20000 242952 20052
rect 49608 19932 49660 19984
rect 267004 19932 267056 19984
rect 178684 18640 178736 18692
rect 281540 18640 281592 18692
rect 60648 18572 60700 18624
rect 238024 18572 238076 18624
rect 20 17280 72 17332
rect 116584 17280 116636 17332
rect 236644 17280 236696 17332
rect 347044 17280 347096 17332
rect 106924 17212 106976 17264
rect 238024 17212 238076 17264
rect 68928 15920 68980 15972
rect 104164 15920 104216 15972
rect 240784 15920 240836 15972
rect 264980 15920 265032 15972
rect 35164 15852 35216 15904
rect 79324 15852 79376 15904
rect 88984 15852 89036 15904
rect 246304 15852 246356 15904
rect 9588 14492 9640 14544
rect 224224 14492 224276 14544
rect 63408 14424 63460 14476
rect 314660 14424 314712 14476
rect 92388 13132 92440 13184
rect 272524 13132 272576 13184
rect 23020 13064 23072 13116
rect 214564 13064 214616 13116
rect 110328 11772 110380 11824
rect 269764 11772 269816 11824
rect 37004 11704 37056 11756
rect 269856 11704 269908 11756
rect 108948 10344 109000 10396
rect 142804 10344 142856 10396
rect 202144 10344 202196 10396
rect 284944 10344 284996 10396
rect 31300 10276 31352 10328
rect 255964 10276 256016 10328
rect 9956 8984 10008 9036
rect 162124 8984 162176 9036
rect 66720 8916 66772 8968
rect 254584 8916 254636 8968
rect 44272 7624 44324 7676
rect 71044 7624 71096 7676
rect 92756 7624 92808 7676
rect 271144 7624 271196 7676
rect 61936 7556 61988 7608
rect 268292 7556 268344 7608
rect 3424 6604 3476 6656
rect 7564 6604 7616 6656
rect 89168 6196 89220 6248
rect 112444 6196 112496 6248
rect 114008 6196 114060 6248
rect 279424 6196 279476 6248
rect 30104 6128 30156 6180
rect 196808 6128 196860 6180
rect 233884 6128 233936 6180
rect 260656 6128 260708 6180
rect 304264 6128 304316 6180
rect 342168 6128 342220 6180
rect 69112 4836 69164 4888
rect 146944 4836 146996 4888
rect 184204 4836 184256 4888
rect 303160 4836 303212 4888
rect 11152 4768 11204 4820
rect 35164 4768 35216 4820
rect 45468 4768 45520 4820
rect 291292 4768 291344 4820
rect 338672 4768 338724 4820
rect 360200 4768 360252 4820
rect 27712 3612 27764 3664
rect 28908 3612 28960 3664
rect 35992 3544 36044 3596
rect 37096 3544 37148 3596
rect 51356 3544 51408 3596
rect 57152 3544 57204 3596
rect 60832 3544 60884 3596
rect 62028 3544 62080 3596
rect 102232 3544 102284 3596
rect 122104 3544 122156 3596
rect 228364 3544 228416 3596
rect 239312 3544 239364 3596
rect 251180 3544 251232 3596
rect 252376 3544 252428 3596
rect 299572 3544 299624 3596
rect 300768 3544 300820 3596
rect 2872 3476 2924 3528
rect 3976 3476 4028 3528
rect 8760 3476 8812 3528
rect 9588 3476 9640 3528
rect 15936 3476 15988 3528
rect 16488 3476 16540 3528
rect 18236 3476 18288 3528
rect 19248 3476 19300 3528
rect 20628 3476 20680 3528
rect 22744 3476 22796 3528
rect 24216 3476 24268 3528
rect 24768 3476 24820 3528
rect 25320 3476 25372 3528
rect 26148 3476 26200 3528
rect 28908 3476 28960 3528
rect 29644 3476 29696 3528
rect 32404 3476 32456 3528
rect 33048 3476 33100 3528
rect 33600 3476 33652 3528
rect 34428 3476 34480 3528
rect 34796 3476 34848 3528
rect 35808 3476 35860 3528
rect 40684 3476 40736 3528
rect 41328 3476 41380 3528
rect 41880 3476 41932 3528
rect 42708 3476 42760 3528
rect 43076 3476 43128 3528
rect 44088 3476 44140 3528
rect 48964 3476 49016 3528
rect 49608 3476 49660 3528
rect 50160 3476 50212 3528
rect 50896 3476 50948 3528
rect 52552 3476 52604 3528
rect 53656 3476 53708 3528
rect 56048 3476 56100 3528
rect 56508 3476 56560 3528
rect 57244 3476 57296 3528
rect 57796 3476 57848 3528
rect 58440 3476 58492 3528
rect 59176 3476 59228 3528
rect 59636 3476 59688 3528
rect 60648 3476 60700 3528
rect 63224 3476 63276 3528
rect 7656 3408 7708 3460
rect 33784 3408 33836 3460
rect 64328 3408 64380 3460
rect 64788 3408 64840 3460
rect 65524 3408 65576 3460
rect 66168 3408 66220 3460
rect 67916 3408 67968 3460
rect 68928 3408 68980 3460
rect 72608 3408 72660 3460
rect 73068 3408 73120 3460
rect 73804 3408 73856 3460
rect 74448 3408 74500 3460
rect 75000 3408 75052 3460
rect 75828 3408 75880 3460
rect 76196 3408 76248 3460
rect 77208 3408 77260 3460
rect 80888 3408 80940 3460
rect 81348 3408 81400 3460
rect 83280 3408 83332 3460
rect 84108 3408 84160 3460
rect 85672 3408 85724 3460
rect 86776 3408 86828 3460
rect 91560 3408 91612 3460
rect 92388 3408 92440 3460
rect 97448 3476 97500 3528
rect 97908 3476 97960 3528
rect 98644 3476 98696 3528
rect 99288 3476 99340 3528
rect 99840 3476 99892 3528
rect 100668 3476 100720 3528
rect 101036 3476 101088 3528
rect 102048 3476 102100 3528
rect 106924 3476 106976 3528
rect 107568 3476 107620 3528
rect 108120 3476 108172 3528
rect 108948 3476 109000 3528
rect 109316 3476 109368 3528
rect 110328 3476 110380 3528
rect 110512 3476 110564 3528
rect 111708 3476 111760 3528
rect 115204 3476 115256 3528
rect 115848 3476 115900 3528
rect 116400 3476 116452 3528
rect 117228 3476 117280 3528
rect 117596 3476 117648 3528
rect 118608 3476 118660 3528
rect 118792 3476 118844 3528
rect 119804 3476 119856 3528
rect 122288 3476 122340 3528
rect 122748 3476 122800 3528
rect 123484 3476 123536 3528
rect 124128 3476 124180 3528
rect 124680 3476 124732 3528
rect 125508 3476 125560 3528
rect 129372 3476 129424 3528
rect 130384 3476 130436 3528
rect 231124 3476 231176 3528
rect 247592 3476 247644 3528
rect 250444 3476 250496 3528
rect 271236 3476 271288 3528
rect 271420 3476 271472 3528
rect 272432 3476 272484 3528
rect 307760 3476 307812 3528
rect 309048 3476 309100 3528
rect 322204 3476 322256 3528
rect 323308 3476 323360 3528
rect 324320 3476 324372 3528
rect 325608 3476 325660 3528
rect 332600 3476 332652 3528
rect 333888 3476 333940 3528
rect 337476 3476 337528 3528
rect 338120 3476 338172 3528
rect 350448 3476 350500 3528
rect 353300 3476 353352 3528
rect 582196 3476 582248 3528
rect 583484 3476 583536 3528
rect 105544 3408 105596 3460
rect 105728 3408 105780 3460
rect 229744 3408 229796 3460
rect 242164 3408 242216 3460
rect 293684 3408 293736 3460
rect 295984 3408 296036 3460
rect 304356 3408 304408 3460
rect 306748 3408 306800 3460
rect 317420 3408 317472 3460
rect 77392 3340 77444 3392
rect 88984 3340 89036 3392
rect 298744 3272 298796 3324
rect 301964 3272 302016 3324
rect 316224 3272 316276 3324
rect 320180 3272 320232 3324
rect 346952 3272 347004 3324
rect 351920 3272 351972 3324
rect 17040 3204 17092 3256
rect 17868 3204 17920 3256
rect 280804 3068 280856 3120
rect 283104 3068 283156 3120
rect 347044 3068 347096 3120
rect 349252 3068 349304 3120
rect 90364 3000 90416 3052
rect 91008 3000 91060 3052
rect 93952 3000 94004 3052
rect 95056 3000 95108 3052
rect 581000 3000 581052 3052
rect 583576 3000 583628 3052
rect 332692 2932 332744 2984
rect 335360 2932 335412 2984
rect 84476 2116 84528 2168
rect 196716 2116 196768 2168
rect 238024 2116 238076 2168
rect 305552 2116 305604 2168
rect 26516 2048 26568 2100
rect 265624 2048 265676 2100
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 702642 8156 703520
rect 8116 702636 8168 702642
rect 8116 702578 8168 702584
rect 24320 698970 24348 703520
rect 24308 698964 24360 698970
rect 24308 698906 24360 698912
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 2778 658200 2834 658209
rect 2778 658135 2834 658144
rect 2792 657014 2820 658135
rect 2780 657008 2832 657014
rect 2780 656950 2832 656956
rect 2780 580508 2832 580514
rect 2780 580450 2832 580456
rect 2792 580009 2820 580450
rect 2778 580000 2834 580009
rect 2778 579935 2834 579944
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 3436 547194 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 22744 670744 22796 670750
rect 22744 670686 22796 670692
rect 4804 657008 4856 657014
rect 4804 656950 4856 656956
rect 3516 632120 3568 632126
rect 3514 632088 3516 632097
rect 3568 632088 3570 632097
rect 3514 632023 3570 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 4816 592686 4844 656950
rect 4804 592680 4856 592686
rect 4804 592622 4856 592628
rect 4804 589348 4856 589354
rect 4804 589290 4856 589296
rect 4816 580514 4844 589290
rect 4804 580508 4856 580514
rect 4804 580450 4856 580456
rect 3514 553888 3570 553897
rect 3514 553823 3516 553832
rect 3568 553823 3570 553832
rect 7564 553852 7616 553858
rect 3516 553794 3568 553800
rect 7564 553794 7616 553800
rect 3424 547188 3476 547194
rect 3424 547130 3476 547136
rect 3424 538348 3476 538354
rect 3424 538290 3476 538296
rect 3436 527921 3464 538290
rect 7576 538218 7604 553794
rect 22756 541686 22784 670686
rect 25504 632120 25556 632126
rect 25504 632062 25556 632068
rect 25516 576162 25544 632062
rect 36544 618316 36596 618322
rect 36544 618258 36596 618264
rect 25504 576156 25556 576162
rect 25504 576098 25556 576104
rect 35808 561740 35860 561746
rect 35808 561682 35860 561688
rect 22744 541680 22796 541686
rect 22744 541622 22796 541628
rect 7564 538212 7616 538218
rect 7564 538154 7616 538160
rect 8208 534744 8260 534750
rect 8208 534686 8260 534692
rect 4804 533384 4856 533390
rect 4804 533326 4856 533332
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 4816 501906 4844 533326
rect 2780 501900 2832 501906
rect 2780 501842 2832 501848
rect 4804 501900 4856 501906
rect 4804 501842 4856 501848
rect 2792 501809 2820 501842
rect 2778 501800 2834 501809
rect 2778 501735 2834 501744
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3344 475386 3372 475623
rect 8220 475386 8248 534686
rect 23388 530596 23440 530602
rect 23388 530538 23440 530544
rect 11704 514820 11756 514826
rect 11704 514762 11756 514768
rect 3332 475380 3384 475386
rect 3332 475322 3384 475328
rect 8208 475380 8260 475386
rect 8208 475322 8260 475328
rect 2778 462632 2834 462641
rect 2778 462567 2780 462576
rect 2832 462567 2834 462576
rect 4804 462596 4856 462602
rect 2780 462538 2832 462544
rect 4804 462538 4856 462544
rect 4816 451246 4844 462538
rect 4804 451240 4856 451246
rect 4804 451182 4856 451188
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 11716 448526 11744 514762
rect 17224 475380 17276 475386
rect 17224 475322 17276 475328
rect 11704 448520 11756 448526
rect 11704 448462 11756 448468
rect 4804 444440 4856 444446
rect 4804 444382 4856 444388
rect 3424 423632 3476 423638
rect 3422 423600 3424 423609
rect 3476 423600 3478 423609
rect 3422 423535 3478 423544
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 2780 398744 2832 398750
rect 2780 398686 2832 398692
rect 2792 397497 2820 398686
rect 2778 397488 2834 397497
rect 2778 397423 2834 397432
rect 3436 389842 3464 410479
rect 4816 398750 4844 444382
rect 15844 428460 15896 428466
rect 15844 428402 15896 428408
rect 4804 398744 4856 398750
rect 4804 398686 4856 398692
rect 3424 389836 3476 389842
rect 3424 389778 3476 389784
rect 7562 382936 7618 382945
rect 7562 382871 7618 382880
rect 4804 381540 4856 381546
rect 4804 381482 4856 381488
rect 3424 373312 3476 373318
rect 3424 373254 3476 373260
rect 3146 371376 3202 371385
rect 3146 371311 3202 371320
rect 3160 370530 3188 371311
rect 3148 370524 3200 370530
rect 3148 370466 3200 370472
rect 3436 358465 3464 373254
rect 3422 358456 3478 358465
rect 3422 358391 3478 358400
rect 3148 346384 3200 346390
rect 3148 346326 3200 346332
rect 3160 345409 3188 346326
rect 3146 345400 3202 345409
rect 3146 345335 3202 345344
rect 4816 320142 4844 381482
rect 7576 370530 7604 382871
rect 7564 370524 7616 370530
rect 7564 370466 7616 370472
rect 11704 370524 11756 370530
rect 11704 370466 11756 370472
rect 7562 327312 7618 327321
rect 7562 327247 7618 327256
rect 4068 320136 4120 320142
rect 4068 320078 4120 320084
rect 4804 320136 4856 320142
rect 4804 320078 4856 320084
rect 4080 319297 4108 320078
rect 4066 319288 4122 319297
rect 4066 319223 4122 319232
rect 3424 306332 3476 306338
rect 3424 306274 3476 306280
rect 3436 306241 3464 306274
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 2778 293176 2834 293185
rect 2778 293111 2834 293120
rect 2792 292874 2820 293111
rect 2780 292868 2832 292874
rect 2780 292810 2832 292816
rect 4080 269822 4108 319223
rect 4804 292868 4856 292874
rect 4804 292810 4856 292816
rect 4068 269816 4120 269822
rect 4068 269758 4120 269764
rect 3422 267200 3478 267209
rect 3422 267135 3478 267144
rect 3436 267034 3464 267135
rect 3424 267028 3476 267034
rect 3424 266970 3476 266976
rect 3424 255264 3476 255270
rect 3424 255206 3476 255212
rect 3436 254153 3464 255206
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3424 241460 3476 241466
rect 3424 241402 3476 241408
rect 3436 241097 3464 241402
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 4816 237386 4844 292810
rect 4804 237380 4856 237386
rect 4804 237322 4856 237328
rect 4802 222320 4858 222329
rect 4802 222255 4858 222264
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3514 206272 3570 206281
rect 3514 206207 3570 206216
rect 3424 202836 3476 202842
rect 3424 202778 3476 202784
rect 3436 201929 3464 202778
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3528 200114 3556 206207
rect 3436 200086 3556 200114
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3436 110673 3464 200086
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 150408 3568 150414
rect 3516 150350 3568 150356
rect 3528 149841 3556 150350
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 4066 76528 4122 76537
rect 4066 76463 4122 76472
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 2780 45552 2832 45558
rect 2778 45520 2780 45529
rect 2832 45520 2834 45529
rect 2778 45455 2834 45464
rect 3976 36576 4028 36582
rect 3976 36518 4028 36524
rect 1400 35216 1452 35222
rect 1400 35158 1452 35164
rect 20 17332 72 17338
rect 20 17274 72 17280
rect 32 16574 60 17274
rect 1412 16574 1440 35158
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 32 16546 152 16574
rect 1412 16546 1716 16574
rect 124 490 152 16546
rect 400 598 612 626
rect 400 490 428 598
rect 124 462 428 490
rect 584 480 612 598
rect 1688 480 1716 16546
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 6497 3464 6598
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 3988 3534 4016 36518
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 2884 480 2912 3470
rect 4080 480 4108 76463
rect 4816 45558 4844 222255
rect 4804 45552 4856 45558
rect 4804 45494 4856 45500
rect 5448 42084 5500 42090
rect 5448 42026 5500 42032
rect 5460 6914 5488 42026
rect 6826 18592 6882 18601
rect 6826 18527 6882 18536
rect 6840 6914 6868 18527
rect 5276 6886 5488 6914
rect 6472 6886 6868 6914
rect 5276 480 5304 6886
rect 6472 480 6500 6886
rect 7576 6662 7604 327247
rect 11716 318102 11744 370466
rect 11704 318096 11756 318102
rect 11704 318038 11756 318044
rect 14464 308440 14516 308446
rect 14464 308382 14516 308388
rect 14476 255270 14504 308382
rect 15856 267034 15884 428402
rect 17236 391241 17264 475322
rect 23400 454034 23428 530538
rect 22744 454028 22796 454034
rect 22744 453970 22796 453976
rect 23388 454028 23440 454034
rect 23388 453970 23440 453976
rect 22756 452674 22784 453970
rect 22744 452668 22796 452674
rect 22744 452610 22796 452616
rect 22756 423638 22784 452610
rect 35820 429146 35848 561682
rect 36556 536110 36584 618258
rect 40052 598262 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 67640 703520 67692 703526
rect 72946 703520 73058 704960
rect 75828 703656 75880 703662
rect 75828 703598 75880 703604
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 67640 703462 67692 703468
rect 59268 703384 59320 703390
rect 59268 703326 59320 703332
rect 57888 702976 57940 702982
rect 57888 702918 57940 702924
rect 55128 702568 55180 702574
rect 55128 702510 55180 702516
rect 40040 598256 40092 598262
rect 40040 598198 40092 598204
rect 53654 590744 53710 590753
rect 53654 590679 53710 590688
rect 52368 587920 52420 587926
rect 52368 587862 52420 587868
rect 48228 585200 48280 585206
rect 48228 585142 48280 585148
rect 47860 576156 47912 576162
rect 47860 576098 47912 576104
rect 47872 575550 47900 576098
rect 47860 575544 47912 575550
rect 47860 575486 47912 575492
rect 48136 575544 48188 575550
rect 48136 575486 48188 575492
rect 43444 565888 43496 565894
rect 43444 565830 43496 565836
rect 39948 560312 40000 560318
rect 39948 560254 40000 560260
rect 36544 536104 36596 536110
rect 36544 536046 36596 536052
rect 39960 511290 39988 560254
rect 41236 547188 41288 547194
rect 41236 547130 41288 547136
rect 41328 547188 41380 547194
rect 41328 547130 41380 547136
rect 41248 542434 41276 547130
rect 41236 542428 41288 542434
rect 41236 542370 41288 542376
rect 39948 511284 40000 511290
rect 39948 511226 40000 511232
rect 39856 435396 39908 435402
rect 39856 435338 39908 435344
rect 34520 429140 34572 429146
rect 34520 429082 34572 429088
rect 35808 429140 35860 429146
rect 35808 429082 35860 429088
rect 34532 428466 34560 429082
rect 34520 428460 34572 428466
rect 34520 428402 34572 428408
rect 22744 423632 22796 423638
rect 22744 423574 22796 423580
rect 17222 391232 17278 391241
rect 17222 391167 17278 391176
rect 33782 387016 33838 387025
rect 33782 386951 33838 386960
rect 33796 346390 33824 386951
rect 39868 375426 39896 435338
rect 39960 425746 39988 511226
rect 40684 448588 40736 448594
rect 40684 448530 40736 448536
rect 39948 425740 40000 425746
rect 39948 425682 40000 425688
rect 39856 375420 39908 375426
rect 39856 375362 39908 375368
rect 39868 373994 39896 375362
rect 39868 373966 39988 373994
rect 33784 346384 33836 346390
rect 33784 346326 33836 346332
rect 25504 330540 25556 330546
rect 25504 330482 25556 330488
rect 17222 328536 17278 328545
rect 17222 328471 17278 328480
rect 15844 267028 15896 267034
rect 15844 266970 15896 266976
rect 14464 255264 14516 255270
rect 14464 255206 14516 255212
rect 15856 231810 15884 266970
rect 15844 231804 15896 231810
rect 15844 231746 15896 231752
rect 14464 220108 14516 220114
rect 14464 220050 14516 220056
rect 14476 150414 14504 220050
rect 14464 150408 14516 150414
rect 14464 150350 14516 150356
rect 16486 77888 16542 77897
rect 16486 77823 16542 77832
rect 13726 69592 13782 69601
rect 13726 69527 13782 69536
rect 12256 42152 12308 42158
rect 12256 42094 12308 42100
rect 12268 16574 12296 42094
rect 12268 16546 12388 16574
rect 9588 14544 9640 14550
rect 9588 14486 9640 14492
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 9600 3534 9628 14486
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 7656 3460 7708 3466
rect 7656 3402 7708 3408
rect 7668 480 7696 3402
rect 8772 480 8800 3470
rect 9968 480 9996 8978
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11164 480 11192 4762
rect 12360 480 12388 16546
rect 13740 6914 13768 69527
rect 15106 53136 15162 53145
rect 15106 53071 15162 53080
rect 15120 6914 15148 53071
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 16500 3534 16528 77823
rect 17236 59362 17264 328471
rect 22744 327140 22796 327146
rect 22744 327082 22796 327088
rect 21362 326224 21418 326233
rect 21362 326159 21418 326168
rect 18604 307080 18656 307086
rect 18604 307022 18656 307028
rect 18616 71738 18644 307022
rect 21376 97986 21404 326159
rect 22756 215286 22784 327082
rect 22744 215280 22796 215286
rect 22744 215222 22796 215228
rect 25516 137970 25544 330482
rect 36544 329112 36596 329118
rect 36544 329054 36596 329060
rect 32404 328500 32456 328506
rect 32404 328442 32456 328448
rect 29644 278792 29696 278798
rect 29644 278734 29696 278740
rect 25504 137964 25556 137970
rect 25504 137906 25556 137912
rect 21364 97980 21416 97986
rect 21364 97922 21416 97928
rect 29656 85542 29684 278734
rect 32416 241466 32444 328442
rect 35164 315308 35216 315314
rect 35164 315250 35216 315256
rect 33784 294024 33836 294030
rect 33784 293966 33836 293972
rect 32404 241460 32456 241466
rect 32404 241402 32456 241408
rect 33796 164218 33824 293966
rect 35176 189038 35204 315250
rect 36556 306338 36584 329054
rect 36544 306332 36596 306338
rect 36544 306274 36596 306280
rect 39960 296682 39988 373966
rect 39948 296676 40000 296682
rect 39948 296618 40000 296624
rect 40696 292534 40724 448530
rect 41340 405006 41368 547130
rect 43456 536790 43484 565830
rect 44088 542428 44140 542434
rect 44088 542370 44140 542376
rect 43444 536784 43496 536790
rect 43444 536726 43496 536732
rect 41328 405000 41380 405006
rect 41328 404942 41380 404948
rect 43996 398132 44048 398138
rect 43996 398074 44048 398080
rect 40684 292528 40736 292534
rect 40684 292470 40736 292476
rect 35900 269816 35952 269822
rect 35900 269758 35952 269764
rect 35912 261526 35940 269758
rect 41328 264988 41380 264994
rect 41328 264930 41380 264936
rect 35900 261520 35952 261526
rect 35900 261462 35952 261468
rect 39304 211812 39356 211818
rect 39304 211754 39356 211760
rect 36542 197976 36598 197985
rect 36542 197911 36598 197920
rect 35164 189032 35216 189038
rect 35164 188974 35216 188980
rect 33784 164212 33836 164218
rect 33784 164154 33836 164160
rect 29644 85536 29696 85542
rect 29644 85478 29696 85484
rect 22006 83464 22062 83473
rect 22006 83399 22062 83408
rect 18604 71732 18656 71738
rect 18604 71674 18656 71680
rect 19246 68232 19302 68241
rect 19246 68167 19302 68176
rect 17224 59356 17276 59362
rect 17224 59298 17276 59304
rect 17866 48920 17922 48929
rect 17866 48855 17922 48864
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 15948 480 15976 3470
rect 17880 3262 17908 48855
rect 19260 3534 19288 68167
rect 22020 6914 22048 83399
rect 34426 82104 34482 82113
rect 34426 82039 34482 82048
rect 22742 78024 22798 78033
rect 22742 77959 22798 77968
rect 21836 6886 22048 6914
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 17040 3256 17092 3262
rect 17040 3198 17092 3204
rect 17868 3256 17920 3262
rect 17868 3198 17920 3204
rect 17052 480 17080 3198
rect 18248 480 18276 3470
rect 19430 3360 19486 3369
rect 19430 3295 19486 3304
rect 19444 480 19472 3295
rect 20640 480 20668 3470
rect 21836 480 21864 6886
rect 22756 3534 22784 77959
rect 26146 59936 26202 59945
rect 26146 59871 26202 59880
rect 24766 21312 24822 21321
rect 24766 21247 24822 21256
rect 23020 13116 23072 13122
rect 23020 13058 23072 13064
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 23032 480 23060 13058
rect 24780 3534 24808 21247
rect 26160 3534 26188 59871
rect 33046 55992 33102 56001
rect 33046 55927 33102 55936
rect 29642 37904 29698 37913
rect 29642 37839 29698 37848
rect 28906 30968 28962 30977
rect 28906 30903 28962 30912
rect 28920 3670 28948 30903
rect 27712 3664 27764 3670
rect 27712 3606 27764 3612
rect 28908 3664 28960 3670
rect 28908 3606 28960 3612
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 24228 480 24256 3470
rect 25332 480 25360 3470
rect 26516 2100 26568 2106
rect 26516 2042 26568 2048
rect 26528 480 26556 2042
rect 27724 480 27752 3606
rect 29656 3534 29684 37839
rect 31300 10328 31352 10334
rect 31300 10270 31352 10276
rect 30104 6180 30156 6186
rect 30104 6122 30156 6128
rect 28908 3528 28960 3534
rect 28908 3470 28960 3476
rect 29644 3528 29696 3534
rect 29644 3470 29696 3476
rect 28920 480 28948 3470
rect 30116 480 30144 6122
rect 31312 480 31340 10270
rect 33060 3534 33088 55927
rect 33782 39264 33838 39273
rect 33782 39199 33838 39208
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 32416 480 32444 3470
rect 33612 480 33640 3470
rect 33796 3466 33824 39199
rect 34440 3534 34468 82039
rect 35806 79520 35862 79529
rect 35806 79455 35862 79464
rect 35164 15904 35216 15910
rect 35164 15846 35216 15852
rect 35176 4826 35204 15846
rect 35164 4820 35216 4826
rect 35164 4762 35216 4768
rect 35820 3534 35848 79455
rect 36556 20670 36584 197911
rect 37188 49020 37240 49026
rect 37188 48962 37240 48968
rect 36544 20664 36596 20670
rect 36544 20606 36596 20612
rect 37004 11756 37056 11762
rect 37004 11698 37056 11704
rect 35992 3596 36044 3602
rect 35992 3538 36044 3544
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 34796 3528 34848 3534
rect 34796 3470 34848 3476
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 33784 3460 33836 3466
rect 33784 3402 33836 3408
rect 34808 480 34836 3470
rect 36004 480 36032 3538
rect 37016 3482 37044 11698
rect 37200 6914 37228 48962
rect 38566 46200 38622 46209
rect 38566 46135 38622 46144
rect 38580 6914 38608 46135
rect 39316 33114 39344 211754
rect 41340 66881 41368 264930
rect 43904 258120 43956 258126
rect 43904 258062 43956 258068
rect 41326 66872 41382 66881
rect 41326 66807 41382 66816
rect 39948 47592 40000 47598
rect 39948 47534 40000 47540
rect 39304 33108 39356 33114
rect 39304 33050 39356 33056
rect 39960 6914 39988 47534
rect 42706 44840 42762 44849
rect 42706 44775 42762 44784
rect 41328 33788 41380 33794
rect 41328 33730 41380 33736
rect 37108 6886 37228 6914
rect 38396 6886 38608 6914
rect 39592 6886 39988 6914
rect 37108 3602 37136 6886
rect 37096 3596 37148 3602
rect 37096 3538 37148 3544
rect 37016 3454 37228 3482
rect 37200 480 37228 3454
rect 38396 480 38424 6886
rect 39592 480 39620 6886
rect 41340 3534 41368 33730
rect 42720 3534 42748 44775
rect 43916 25537 43944 258062
rect 44008 239465 44036 398074
rect 44100 396778 44128 542370
rect 48148 454714 48176 575486
rect 48240 460222 48268 585142
rect 50896 582412 50948 582418
rect 50896 582354 50948 582360
rect 49608 536104 49660 536110
rect 49608 536046 49660 536052
rect 48228 460216 48280 460222
rect 48228 460158 48280 460164
rect 48136 454708 48188 454714
rect 48136 454650 48188 454656
rect 48136 431996 48188 432002
rect 48136 431938 48188 431944
rect 44088 396772 44140 396778
rect 44088 396714 44140 396720
rect 46848 294092 46900 294098
rect 46848 294034 46900 294040
rect 43994 239456 44050 239465
rect 43994 239391 44050 239400
rect 46860 213246 46888 294034
rect 48148 227662 48176 431938
rect 49620 389162 49648 536046
rect 50804 451308 50856 451314
rect 50804 451250 50856 451256
rect 49608 389156 49660 389162
rect 49608 389098 49660 389104
rect 49608 344344 49660 344350
rect 49608 344286 49660 344292
rect 48228 285728 48280 285734
rect 48228 285670 48280 285676
rect 48136 227656 48188 227662
rect 48136 227598 48188 227604
rect 46848 213240 46900 213246
rect 46848 213182 46900 213188
rect 48134 62792 48190 62801
rect 48134 62727 48190 62736
rect 44088 26920 44140 26926
rect 44088 26862 44140 26868
rect 43902 25528 43958 25537
rect 43902 25463 43958 25472
rect 44100 3534 44128 26862
rect 46846 22672 46902 22681
rect 46846 22607 46902 22616
rect 44272 7676 44324 7682
rect 44272 7618 44324 7624
rect 40684 3528 40736 3534
rect 40684 3470 40736 3476
rect 41328 3528 41380 3534
rect 41328 3470 41380 3476
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 44088 3528 44140 3534
rect 44088 3470 44140 3476
rect 40696 480 40724 3470
rect 41892 480 41920 3470
rect 43088 480 43116 3470
rect 44284 480 44312 7618
rect 46860 6914 46888 22607
rect 48148 6914 48176 62727
rect 46676 6886 46888 6914
rect 47872 6886 48176 6914
rect 45468 4820 45520 4826
rect 45468 4762 45520 4768
rect 45480 480 45508 4762
rect 46676 480 46704 6886
rect 47872 480 47900 6886
rect 48240 2009 48268 285670
rect 49620 220726 49648 344286
rect 50816 329798 50844 451250
rect 50908 449886 50936 582354
rect 51724 564392 51776 564398
rect 51724 564334 51776 564340
rect 50988 557592 51040 557598
rect 50988 557534 51040 557540
rect 50896 449880 50948 449886
rect 50896 449822 50948 449828
rect 51000 421598 51028 557534
rect 51736 431934 51764 564334
rect 52276 461644 52328 461650
rect 52276 461586 52328 461592
rect 52184 433356 52236 433362
rect 52184 433298 52236 433304
rect 51724 431928 51776 431934
rect 51724 431870 51776 431876
rect 50988 421592 51040 421598
rect 50988 421534 51040 421540
rect 50896 401600 50948 401606
rect 50896 401542 50948 401548
rect 50528 329792 50580 329798
rect 50528 329734 50580 329740
rect 50804 329792 50856 329798
rect 50804 329734 50856 329740
rect 50540 329118 50568 329734
rect 50528 329112 50580 329118
rect 50528 329054 50580 329060
rect 50804 298784 50856 298790
rect 50804 298726 50856 298732
rect 50816 227633 50844 298726
rect 50908 239601 50936 401542
rect 52196 376038 52224 433298
rect 52288 386374 52316 461586
rect 52380 458250 52408 587862
rect 53668 465730 53696 590679
rect 55036 574796 55088 574802
rect 55036 574738 55088 574744
rect 53748 566500 53800 566506
rect 53748 566442 53800 566448
rect 53656 465724 53708 465730
rect 53656 465666 53708 465672
rect 52368 458244 52420 458250
rect 52368 458186 52420 458192
rect 53564 458244 53616 458250
rect 53564 458186 53616 458192
rect 52460 436076 52512 436082
rect 52460 436018 52512 436024
rect 52472 435402 52500 436018
rect 52460 435396 52512 435402
rect 52460 435338 52512 435344
rect 52276 386368 52328 386374
rect 52276 386310 52328 386316
rect 52276 384328 52328 384334
rect 52276 384270 52328 384276
rect 52184 376032 52236 376038
rect 52184 375974 52236 375980
rect 50988 282940 51040 282946
rect 50988 282882 51040 282888
rect 50894 239592 50950 239601
rect 50894 239527 50950 239536
rect 50802 227624 50858 227633
rect 50802 227559 50858 227568
rect 49608 220720 49660 220726
rect 49608 220662 49660 220668
rect 49620 220114 49648 220662
rect 49608 220108 49660 220114
rect 49608 220050 49660 220056
rect 50894 79384 50950 79393
rect 50894 79319 50950 79328
rect 49608 19984 49660 19990
rect 49608 19926 49660 19932
rect 49620 3534 49648 19926
rect 50908 3534 50936 79319
rect 51000 21418 51028 282882
rect 52184 271924 52236 271930
rect 52184 271866 52236 271872
rect 52092 267028 52144 267034
rect 52092 266970 52144 266976
rect 52104 236609 52132 266970
rect 52090 236600 52146 236609
rect 52090 236535 52146 236544
rect 52196 218006 52224 271866
rect 52288 262886 52316 384270
rect 53576 378826 53604 458186
rect 53654 446040 53710 446049
rect 53654 445975 53710 445984
rect 53564 378820 53616 378826
rect 53564 378762 53616 378768
rect 53668 345014 53696 445975
rect 53760 436082 53788 566442
rect 55048 450566 55076 574738
rect 55140 564398 55168 702510
rect 57796 567248 57848 567254
rect 57796 567190 57848 567196
rect 55128 564392 55180 564398
rect 55128 564334 55180 564340
rect 56508 558952 56560 558958
rect 56508 558894 56560 558900
rect 55128 539640 55180 539646
rect 55128 539582 55180 539588
rect 55036 450560 55088 450566
rect 55036 450502 55088 450508
rect 55034 445904 55090 445913
rect 55034 445839 55090 445848
rect 53748 436076 53800 436082
rect 53748 436018 53800 436024
rect 53668 344986 53788 345014
rect 53760 331362 53788 344986
rect 54852 337408 54904 337414
rect 54852 337350 54904 337356
rect 53748 331356 53800 331362
rect 53748 331298 53800 331304
rect 52368 324352 52420 324358
rect 52368 324294 52420 324300
rect 52276 262880 52328 262886
rect 52276 262822 52328 262828
rect 52276 253972 52328 253978
rect 52276 253914 52328 253920
rect 52184 218000 52236 218006
rect 52184 217942 52236 217948
rect 52288 195974 52316 253914
rect 52276 195968 52328 195974
rect 52276 195910 52328 195916
rect 52380 33833 52408 324294
rect 53564 313336 53616 313342
rect 53564 313278 53616 313284
rect 53576 224913 53604 313278
rect 53656 309188 53708 309194
rect 53656 309130 53708 309136
rect 53562 224904 53618 224913
rect 53562 224839 53618 224848
rect 53668 208350 53696 309130
rect 53760 290057 53788 331298
rect 53840 318096 53892 318102
rect 53840 318038 53892 318044
rect 53852 317490 53880 318038
rect 53840 317484 53892 317490
rect 53840 317426 53892 317432
rect 53746 290048 53802 290057
rect 53746 289983 53802 289992
rect 53748 270564 53800 270570
rect 53748 270506 53800 270512
rect 53656 208344 53708 208350
rect 53656 208286 53708 208292
rect 53760 72457 53788 270506
rect 54864 237386 54892 337350
rect 54944 317484 54996 317490
rect 54944 317426 54996 317432
rect 54852 237380 54904 237386
rect 54852 237322 54904 237328
rect 54956 198665 54984 317426
rect 55048 264246 55076 445839
rect 55140 393310 55168 539582
rect 56520 534070 56548 558894
rect 57520 545760 57572 545766
rect 57520 545702 57572 545708
rect 56508 534064 56560 534070
rect 56508 534006 56560 534012
rect 56520 424386 56548 534006
rect 56508 424380 56560 424386
rect 56508 424322 56560 424328
rect 56508 419552 56560 419558
rect 56508 419494 56560 419500
rect 55128 393304 55180 393310
rect 55128 393246 55180 393252
rect 56520 331226 56548 419494
rect 57532 401606 57560 545702
rect 57612 471300 57664 471306
rect 57612 471242 57664 471248
rect 57520 401600 57572 401606
rect 57520 401542 57572 401548
rect 57624 389230 57652 471242
rect 57808 438190 57836 567190
rect 57900 543794 57928 702918
rect 59176 586560 59228 586566
rect 59176 586502 59228 586508
rect 58900 554804 58952 554810
rect 58900 554746 58952 554752
rect 57888 543788 57940 543794
rect 57888 543730 57940 543736
rect 57796 438184 57848 438190
rect 57796 438126 57848 438132
rect 58912 418130 58940 554746
rect 59084 468512 59136 468518
rect 59084 468454 59136 468460
rect 58992 425740 59044 425746
rect 58992 425682 59044 425688
rect 59004 425134 59032 425682
rect 58992 425128 59044 425134
rect 58992 425070 59044 425076
rect 58900 418124 58952 418130
rect 58900 418066 58952 418072
rect 57796 414724 57848 414730
rect 57796 414666 57848 414672
rect 57704 405000 57756 405006
rect 57704 404942 57756 404948
rect 57716 403646 57744 404942
rect 57704 403640 57756 403646
rect 57704 403582 57756 403588
rect 57612 389224 57664 389230
rect 57612 389166 57664 389172
rect 56508 331220 56560 331226
rect 56508 331162 56560 331168
rect 56520 330546 56548 331162
rect 56508 330540 56560 330546
rect 56508 330482 56560 330488
rect 56508 317552 56560 317558
rect 56508 317494 56560 317500
rect 55128 285796 55180 285802
rect 55128 285738 55180 285744
rect 55036 264240 55088 264246
rect 55036 264182 55088 264188
rect 55036 263696 55088 263702
rect 55036 263638 55088 263644
rect 55048 219201 55076 263638
rect 55034 219192 55090 219201
rect 55034 219127 55090 219136
rect 54942 198656 54998 198665
rect 54942 198591 54998 198600
rect 53746 72448 53802 72457
rect 53746 72383 53802 72392
rect 53746 64152 53802 64161
rect 53746 64087 53802 64096
rect 52366 33824 52422 33833
rect 52366 33759 52422 33768
rect 53656 28280 53708 28286
rect 53656 28222 53708 28228
rect 50988 21412 51040 21418
rect 50988 21354 51040 21360
rect 51356 3596 51408 3602
rect 51356 3538 51408 3544
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 49608 3528 49660 3534
rect 49608 3470 49660 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50896 3528 50948 3534
rect 50896 3470 50948 3476
rect 48226 2000 48282 2009
rect 48226 1935 48282 1944
rect 48976 480 49004 3470
rect 50172 480 50200 3470
rect 51368 480 51396 3538
rect 53668 3534 53696 28222
rect 52552 3528 52604 3534
rect 52552 3470 52604 3476
rect 53656 3528 53708 3534
rect 53656 3470 53708 3476
rect 52564 480 52592 3470
rect 53760 480 53788 64087
rect 55036 37936 55088 37942
rect 55036 37878 55088 37884
rect 55048 6914 55076 37878
rect 55140 29617 55168 285738
rect 56416 281580 56468 281586
rect 56416 281522 56468 281528
rect 56324 258188 56376 258194
rect 56324 258130 56376 258136
rect 56336 231169 56364 258130
rect 56322 231160 56378 231169
rect 56322 231095 56378 231104
rect 56428 217977 56456 281522
rect 56414 217968 56470 217977
rect 56414 217903 56470 217912
rect 56520 71233 56548 317494
rect 57612 273964 57664 273970
rect 57612 273906 57664 273912
rect 57624 229090 57652 273906
rect 57716 244934 57744 403582
rect 57704 244928 57756 244934
rect 57704 244870 57756 244876
rect 57808 241505 57836 414666
rect 59004 358057 59032 425070
rect 59096 391270 59124 468454
rect 59188 463010 59216 586502
rect 59280 553518 59308 703326
rect 62028 703180 62080 703186
rect 62028 703122 62080 703128
rect 61934 590880 61990 590889
rect 61934 590815 61990 590824
rect 60556 568608 60608 568614
rect 60556 568550 60608 568556
rect 59268 553512 59320 553518
rect 59268 553454 59320 553460
rect 59176 463004 59228 463010
rect 59176 462946 59228 462952
rect 60464 446412 60516 446418
rect 60464 446354 60516 446360
rect 59176 444508 59228 444514
rect 59176 444450 59228 444456
rect 59084 391264 59136 391270
rect 59084 391206 59136 391212
rect 58990 358048 59046 358057
rect 58990 357983 59046 357992
rect 59084 325712 59136 325718
rect 59084 325654 59136 325660
rect 57888 303680 57940 303686
rect 57888 303622 57940 303628
rect 57794 241496 57850 241505
rect 57794 241431 57850 241440
rect 57612 229084 57664 229090
rect 57612 229026 57664 229032
rect 56506 71224 56562 71233
rect 56506 71159 56562 71168
rect 57244 40724 57296 40730
rect 57244 40666 57296 40672
rect 55126 29608 55182 29617
rect 55126 29543 55182 29552
rect 56508 22772 56560 22778
rect 56508 22714 56560 22720
rect 54956 6886 55076 6914
rect 54956 480 54984 6886
rect 56520 3534 56548 22714
rect 57256 6914 57284 40666
rect 57794 35184 57850 35193
rect 57794 35119 57850 35128
rect 57164 6886 57284 6914
rect 57164 3602 57192 6886
rect 57152 3596 57204 3602
rect 57152 3538 57204 3544
rect 57808 3534 57836 35119
rect 57900 32473 57928 303622
rect 58992 261520 59044 261526
rect 58992 261462 59044 261468
rect 59004 260914 59032 261462
rect 58992 260908 59044 260914
rect 58992 260850 59044 260856
rect 59004 232558 59032 260850
rect 58992 232552 59044 232558
rect 58992 232494 59044 232500
rect 59096 230489 59124 325654
rect 59188 252686 59216 444450
rect 60372 442264 60424 442270
rect 60372 442206 60424 442212
rect 60384 370530 60412 442206
rect 60476 383654 60504 446354
rect 60568 439074 60596 568550
rect 60648 549296 60700 549302
rect 60648 549238 60700 549244
rect 60556 439068 60608 439074
rect 60556 439010 60608 439016
rect 60660 408474 60688 549238
rect 61844 456068 61896 456074
rect 61844 456010 61896 456016
rect 61752 453348 61804 453354
rect 61752 453290 61804 453296
rect 60648 408468 60700 408474
rect 60648 408410 60700 408416
rect 61764 386306 61792 453290
rect 61856 389094 61884 456010
rect 61948 451926 61976 590815
rect 62040 547806 62068 703122
rect 66168 702500 66220 702506
rect 66168 702442 66220 702448
rect 66074 581632 66130 581641
rect 66074 581567 66130 581576
rect 64788 579692 64840 579698
rect 64788 579634 64840 579640
rect 63316 571396 63368 571402
rect 63316 571338 63368 571344
rect 62028 547800 62080 547806
rect 62028 547742 62080 547748
rect 62040 547194 62068 547742
rect 62028 547188 62080 547194
rect 62028 547130 62080 547136
rect 62028 543788 62080 543794
rect 62028 543730 62080 543736
rect 61936 451920 61988 451926
rect 61936 451862 61988 451868
rect 62040 398138 62068 543730
rect 63328 475522 63356 571338
rect 64144 553512 64196 553518
rect 64144 553454 64196 553460
rect 63408 547936 63460 547942
rect 63408 547878 63460 547884
rect 63316 475516 63368 475522
rect 63316 475458 63368 475464
rect 63316 457496 63368 457502
rect 63316 457438 63368 457444
rect 63224 424380 63276 424386
rect 63224 424322 63276 424328
rect 62028 398132 62080 398138
rect 62028 398074 62080 398080
rect 61936 393304 61988 393310
rect 61934 393272 61936 393281
rect 61988 393272 61990 393281
rect 61934 393207 61990 393216
rect 61844 389088 61896 389094
rect 61844 389030 61896 389036
rect 61752 386300 61804 386306
rect 61752 386242 61804 386248
rect 60464 383648 60516 383654
rect 60464 383590 60516 383596
rect 60372 370524 60424 370530
rect 60372 370466 60424 370472
rect 62028 369164 62080 369170
rect 62028 369106 62080 369112
rect 61752 341012 61804 341018
rect 61752 340954 61804 340960
rect 60556 340944 60608 340950
rect 60556 340886 60608 340892
rect 60464 334620 60516 334626
rect 60464 334562 60516 334568
rect 59268 334008 59320 334014
rect 59268 333950 59320 333956
rect 59176 252680 59228 252686
rect 59176 252622 59228 252628
rect 59176 247104 59228 247110
rect 59176 247046 59228 247052
rect 59082 230480 59138 230489
rect 59082 230415 59138 230424
rect 59188 75313 59216 247046
rect 59174 75304 59230 75313
rect 59174 75239 59230 75248
rect 59176 61396 59228 61402
rect 59176 61338 59228 61344
rect 57886 32464 57942 32473
rect 57886 32399 57942 32408
rect 59188 3534 59216 61338
rect 59280 54505 59308 333950
rect 60476 303618 60504 334562
rect 60464 303612 60516 303618
rect 60464 303554 60516 303560
rect 60568 300830 60596 340886
rect 60648 322992 60700 322998
rect 60648 322934 60700 322940
rect 60556 300824 60608 300830
rect 60556 300766 60608 300772
rect 60556 287088 60608 287094
rect 60556 287030 60608 287036
rect 60464 278792 60516 278798
rect 60464 278734 60516 278740
rect 60476 237969 60504 278734
rect 60462 237960 60518 237969
rect 60462 237895 60518 237904
rect 60568 216617 60596 287030
rect 60554 216608 60610 216617
rect 60554 216543 60610 216552
rect 60660 65521 60688 322934
rect 61658 313440 61714 313449
rect 61658 313375 61714 313384
rect 61672 313342 61700 313375
rect 61660 313336 61712 313342
rect 61660 313278 61712 313284
rect 61764 306406 61792 340954
rect 61844 335436 61896 335442
rect 61844 335378 61896 335384
rect 61752 306400 61804 306406
rect 61752 306342 61804 306348
rect 61856 289270 61884 335378
rect 61936 321632 61988 321638
rect 61936 321574 61988 321580
rect 61844 289264 61896 289270
rect 61844 289206 61896 289212
rect 61752 271992 61804 271998
rect 61752 271934 61804 271940
rect 61764 235278 61792 271934
rect 61844 256760 61896 256766
rect 61844 256702 61896 256708
rect 61752 235272 61804 235278
rect 61752 235214 61804 235220
rect 61856 193225 61884 256702
rect 61948 235346 61976 321574
rect 62040 267714 62068 369106
rect 63236 362273 63264 424322
rect 63328 385014 63356 457438
rect 63420 406638 63448 547878
rect 64156 414730 64184 553454
rect 64800 532030 64828 579634
rect 65982 572928 66038 572937
rect 65982 572863 66038 572872
rect 65522 564496 65578 564505
rect 65522 564431 65578 564440
rect 64788 532024 64840 532030
rect 64788 531966 64840 531972
rect 64696 449200 64748 449206
rect 64696 449142 64748 449148
rect 64144 414724 64196 414730
rect 64144 414666 64196 414672
rect 63408 406632 63460 406638
rect 63408 406574 63460 406580
rect 64604 406632 64656 406638
rect 64604 406574 64656 406580
rect 64616 406162 64644 406574
rect 64604 406156 64656 406162
rect 64604 406098 64656 406104
rect 64616 385665 64644 406098
rect 64708 387802 64736 449142
rect 65536 433362 65564 564431
rect 65996 539714 66024 572863
rect 65984 539708 66036 539714
rect 65984 539650 66036 539656
rect 66088 464370 66116 581567
rect 66180 546417 66208 702442
rect 67456 599616 67508 599622
rect 67456 599558 67508 599564
rect 66810 588296 66866 588305
rect 66810 588231 66866 588240
rect 66824 587926 66852 588231
rect 66812 587920 66864 587926
rect 66812 587862 66864 587868
rect 66260 586560 66312 586566
rect 66258 586528 66260 586537
rect 66312 586528 66314 586537
rect 66258 586463 66314 586472
rect 66810 582448 66866 582457
rect 66810 582383 66812 582392
rect 66864 582383 66866 582392
rect 66812 582354 66864 582360
rect 66810 579728 66866 579737
rect 66810 579663 66812 579672
rect 66864 579663 66866 579672
rect 66812 579634 66864 579640
rect 66902 575648 66958 575657
rect 66902 575583 66958 575592
rect 66916 575550 66944 575583
rect 66904 575544 66956 575550
rect 66904 575486 66956 575492
rect 67468 575385 67496 599558
rect 67548 596828 67600 596834
rect 67548 596770 67600 596776
rect 67454 575376 67510 575385
rect 67454 575311 67510 575320
rect 67468 574802 67496 575311
rect 67456 574796 67508 574802
rect 67456 574738 67508 574744
rect 66442 571840 66498 571849
rect 66442 571775 66498 571784
rect 66456 571402 66484 571775
rect 66444 571396 66496 571402
rect 66444 571338 66496 571344
rect 67362 570208 67418 570217
rect 67362 570143 67418 570152
rect 66902 568848 66958 568857
rect 66902 568783 66958 568792
rect 66916 568614 66944 568783
rect 66904 568608 66956 568614
rect 66904 568550 66956 568556
rect 66902 567488 66958 567497
rect 66902 567423 66958 567432
rect 66916 567254 66944 567423
rect 66904 567248 66956 567254
rect 66904 567190 66956 567196
rect 66812 564392 66864 564398
rect 66810 564360 66812 564369
rect 66864 564360 66866 564369
rect 66810 564295 66866 564304
rect 66810 561776 66866 561785
rect 66810 561711 66812 561720
rect 66864 561711 66866 561720
rect 66812 561682 66864 561688
rect 66534 560552 66590 560561
rect 66534 560487 66590 560496
rect 66548 560318 66576 560487
rect 66536 560312 66588 560318
rect 66536 560254 66588 560260
rect 66534 559192 66590 559201
rect 66534 559127 66590 559136
rect 66548 558958 66576 559127
rect 66536 558952 66588 558958
rect 66536 558894 66588 558900
rect 66902 556336 66958 556345
rect 66902 556271 66958 556280
rect 66626 554976 66682 554985
rect 66626 554911 66682 554920
rect 66640 554810 66668 554911
rect 66628 554804 66680 554810
rect 66628 554746 66680 554752
rect 66534 553752 66590 553761
rect 66534 553687 66590 553696
rect 66548 553518 66576 553687
rect 66536 553512 66588 553518
rect 66536 553454 66588 553460
rect 66442 549672 66498 549681
rect 66442 549607 66498 549616
rect 66456 549302 66484 549607
rect 66444 549296 66496 549302
rect 66444 549238 66496 549244
rect 66534 548312 66590 548321
rect 66534 548247 66590 548256
rect 66548 547942 66576 548247
rect 66536 547936 66588 547942
rect 66536 547878 66588 547884
rect 66628 547800 66680 547806
rect 66628 547742 66680 547748
rect 66640 547641 66668 547742
rect 66626 547632 66682 547641
rect 66626 547567 66682 547576
rect 66166 546408 66222 546417
rect 66166 546343 66222 546352
rect 66180 545766 66208 546343
rect 66168 545760 66220 545766
rect 66168 545702 66220 545708
rect 66810 544096 66866 544105
rect 66810 544031 66866 544040
rect 66824 543794 66852 544031
rect 66812 543788 66864 543794
rect 66812 543730 66864 543736
rect 66810 542736 66866 542745
rect 66810 542671 66866 542680
rect 66824 542434 66852 542671
rect 66812 542428 66864 542434
rect 66812 542370 66864 542376
rect 66168 529236 66220 529242
rect 66168 529178 66220 529184
rect 66076 464364 66128 464370
rect 66076 464306 66128 464312
rect 65982 448624 66038 448633
rect 65982 448559 66038 448568
rect 65524 433356 65576 433362
rect 65524 433298 65576 433304
rect 64788 421592 64840 421598
rect 64788 421534 64840 421540
rect 64696 387796 64748 387802
rect 64696 387738 64748 387744
rect 64602 385656 64658 385665
rect 64602 385591 64658 385600
rect 63316 385008 63368 385014
rect 63316 384950 63368 384956
rect 63222 362264 63278 362273
rect 63222 362199 63278 362208
rect 64800 350849 64828 421534
rect 65524 418124 65576 418130
rect 65524 418066 65576 418072
rect 64786 350840 64842 350849
rect 64786 350775 64842 350784
rect 63316 349852 63368 349858
rect 63316 349794 63368 349800
rect 63224 339584 63276 339590
rect 63224 339526 63276 339532
rect 63236 306338 63264 339526
rect 63328 315994 63356 349794
rect 64602 337376 64658 337385
rect 64602 337311 64658 337320
rect 63408 329860 63460 329866
rect 63408 329802 63460 329808
rect 63316 315988 63368 315994
rect 63316 315930 63368 315936
rect 63328 315314 63356 315930
rect 63316 315308 63368 315314
rect 63316 315250 63368 315256
rect 63224 306332 63276 306338
rect 63224 306274 63276 306280
rect 63316 299600 63368 299606
rect 63316 299542 63368 299548
rect 63132 280220 63184 280226
rect 63132 280162 63184 280168
rect 62028 267708 62080 267714
rect 62028 267650 62080 267656
rect 62120 262880 62172 262886
rect 62120 262822 62172 262828
rect 62132 262274 62160 262822
rect 62120 262268 62172 262274
rect 62120 262210 62172 262216
rect 62028 248464 62080 248470
rect 62028 248406 62080 248412
rect 61936 235340 61988 235346
rect 61936 235282 61988 235288
rect 61842 193216 61898 193225
rect 61842 193151 61898 193160
rect 62040 69737 62068 248406
rect 63144 233918 63172 280162
rect 63224 262268 63276 262274
rect 63224 262210 63276 262216
rect 63132 233912 63184 233918
rect 63132 233854 63184 233860
rect 63236 200025 63264 262210
rect 63328 223553 63356 299542
rect 63314 223544 63370 223553
rect 63314 223479 63370 223488
rect 63222 200016 63278 200025
rect 63222 199951 63278 199960
rect 62026 69728 62082 69737
rect 62026 69663 62082 69672
rect 60646 65512 60702 65521
rect 60646 65447 60702 65456
rect 59266 54496 59322 54505
rect 59266 54431 59322 54440
rect 62026 50280 62082 50289
rect 62026 50215 62082 50224
rect 60648 18624 60700 18630
rect 60648 18566 60700 18572
rect 60660 3534 60688 18566
rect 61936 7608 61988 7614
rect 61936 7550 61988 7556
rect 60832 3596 60884 3602
rect 60832 3538 60884 3544
rect 56048 3528 56100 3534
rect 56048 3470 56100 3476
rect 56508 3528 56560 3534
rect 56508 3470 56560 3476
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 57796 3528 57848 3534
rect 57796 3470 57848 3476
rect 58440 3528 58492 3534
rect 58440 3470 58492 3476
rect 59176 3528 59228 3534
rect 59176 3470 59228 3476
rect 59636 3528 59688 3534
rect 59636 3470 59688 3476
rect 60648 3528 60700 3534
rect 60648 3470 60700 3476
rect 56060 480 56088 3470
rect 57256 480 57284 3470
rect 58452 480 58480 3470
rect 59648 480 59676 3470
rect 60844 480 60872 3538
rect 61948 3482 61976 7550
rect 62040 3602 62068 50215
rect 63420 14482 63448 329802
rect 64420 318844 64472 318850
rect 64420 318786 64472 318792
rect 64432 68377 64460 318786
rect 64616 311846 64644 337311
rect 64694 335608 64750 335617
rect 64694 335543 64750 335552
rect 64604 311840 64656 311846
rect 64604 311782 64656 311788
rect 64708 302190 64736 335543
rect 64800 313274 64828 350775
rect 64788 313268 64840 313274
rect 64788 313210 64840 313216
rect 64696 302184 64748 302190
rect 64696 302126 64748 302132
rect 65536 291174 65564 418066
rect 65996 388929 66024 448559
rect 66076 438184 66128 438190
rect 66076 438126 66128 438132
rect 65982 388920 66038 388929
rect 65982 388855 66038 388864
rect 66088 360913 66116 438126
rect 66180 388385 66208 529178
rect 66536 438184 66588 438190
rect 66536 438126 66588 438132
rect 66548 437753 66576 438126
rect 66534 437744 66590 437753
rect 66534 437679 66590 437688
rect 66812 436076 66864 436082
rect 66812 436018 66864 436024
rect 66824 435305 66852 436018
rect 66810 435296 66866 435305
rect 66810 435231 66866 435240
rect 66444 433288 66496 433294
rect 66444 433230 66496 433236
rect 66456 433129 66484 433230
rect 66442 433120 66498 433129
rect 66442 433055 66498 433064
rect 66812 431928 66864 431934
rect 66812 431870 66864 431876
rect 66824 430953 66852 431870
rect 66810 430944 66866 430953
rect 66810 430879 66866 430888
rect 66812 429140 66864 429146
rect 66812 429082 66864 429088
rect 66824 428505 66852 429082
rect 66810 428496 66866 428505
rect 66810 428431 66866 428440
rect 66810 426320 66866 426329
rect 66810 426255 66866 426264
rect 66824 425134 66852 426255
rect 66812 425128 66864 425134
rect 66812 425070 66864 425076
rect 66812 424380 66864 424386
rect 66812 424322 66864 424328
rect 66824 424153 66852 424322
rect 66810 424144 66866 424153
rect 66810 424079 66866 424088
rect 66810 421968 66866 421977
rect 66810 421903 66866 421912
rect 66824 421598 66852 421903
rect 66812 421592 66864 421598
rect 66812 421534 66864 421540
rect 66916 419558 66944 556271
rect 67086 541784 67142 541793
rect 67086 541719 67142 541728
rect 67100 541686 67128 541719
rect 67088 541680 67140 541686
rect 67088 541622 67140 541628
rect 67100 539510 67128 541622
rect 67088 539504 67140 539510
rect 67088 539446 67140 539452
rect 67376 442950 67404 570143
rect 67560 566817 67588 596770
rect 67546 566808 67602 566817
rect 67546 566743 67602 566752
rect 67560 566506 67588 566743
rect 67548 566500 67600 566506
rect 67548 566442 67600 566448
rect 67652 558929 67680 703462
rect 71044 702840 71096 702846
rect 71044 702782 71096 702788
rect 69020 592680 69072 592686
rect 69020 592622 69072 592628
rect 67730 589928 67786 589937
rect 67730 589863 67786 589872
rect 67744 585857 67772 589863
rect 69032 588962 69060 592622
rect 71056 590889 71084 702782
rect 72988 699825 73016 703520
rect 73068 703316 73120 703322
rect 73068 703258 73120 703264
rect 72974 699816 73030 699825
rect 72974 699751 73030 699760
rect 73080 596174 73108 703258
rect 75840 596174 75868 703598
rect 86868 703588 86920 703594
rect 86868 703530 86920 703536
rect 83464 700324 83516 700330
rect 83464 700266 83516 700272
rect 79324 698964 79376 698970
rect 79324 698906 79376 698912
rect 79336 600302 79364 698906
rect 79324 600296 79376 600302
rect 79324 600238 79376 600244
rect 79968 600296 80020 600302
rect 79968 600238 80020 600244
rect 79980 599010 80008 600238
rect 79968 599004 80020 599010
rect 79968 598946 80020 598952
rect 72988 596146 73108 596174
rect 75748 596146 75868 596174
rect 72988 592034 73016 596146
rect 75644 592136 75696 592142
rect 75644 592078 75696 592084
rect 72896 592006 73016 592034
rect 72422 591016 72478 591025
rect 72422 590951 72478 590960
rect 71042 590880 71098 590889
rect 71042 590815 71098 590824
rect 70308 590776 70360 590782
rect 70308 590718 70360 590724
rect 70320 589098 70348 590718
rect 70104 589070 70348 589098
rect 71056 589098 71084 590815
rect 72436 589098 72464 590951
rect 72896 589422 72924 592006
rect 75184 590776 75236 590782
rect 73618 590744 73674 590753
rect 75184 590718 75236 590724
rect 73618 590679 73674 590688
rect 72884 589416 72936 589422
rect 72884 589358 72936 589364
rect 71056 589070 71208 589098
rect 72128 589070 72464 589098
rect 69032 588934 69520 588962
rect 69492 588674 69520 588934
rect 72896 588826 72924 589358
rect 73632 589098 73660 590679
rect 75196 589966 75224 590718
rect 75184 589960 75236 589966
rect 75184 589902 75236 589908
rect 75656 589354 75684 592078
rect 74862 589348 74914 589354
rect 74862 589290 74914 589296
rect 75644 589348 75696 589354
rect 75644 589290 75696 589296
rect 73632 589070 73968 589098
rect 74874 589084 74902 589290
rect 75748 589234 75776 596146
rect 79784 594856 79836 594862
rect 79784 594798 79836 594804
rect 77944 592068 77996 592074
rect 77944 592010 77996 592016
rect 77022 590744 77078 590753
rect 77022 590679 77078 590688
rect 75656 589206 75776 589234
rect 75656 588849 75684 589206
rect 77036 589098 77064 590679
rect 77956 589098 77984 592010
rect 78404 590708 78456 590714
rect 78404 590650 78456 590656
rect 76728 589070 77064 589098
rect 77648 589070 77984 589098
rect 75642 588840 75698 588849
rect 72896 588798 73048 588826
rect 78416 588826 78444 590650
rect 79796 589098 79824 594798
rect 79980 590730 80008 598946
rect 83476 596174 83504 700266
rect 83476 596146 83780 596174
rect 83462 592104 83518 592113
rect 83462 592039 83518 592048
rect 82542 590880 82598 590889
rect 82542 590815 82598 590824
rect 79980 590702 80100 590730
rect 79488 589070 79824 589098
rect 80072 589098 80100 590702
rect 81346 590608 81402 590617
rect 81346 590543 81402 590552
rect 81360 589274 81388 590543
rect 81314 589246 81388 589274
rect 80072 589070 80408 589098
rect 81314 589084 81342 589246
rect 82556 589098 82584 590815
rect 82634 590744 82690 590753
rect 82634 590679 82690 590688
rect 82648 589286 82676 590679
rect 82636 589280 82688 589286
rect 82636 589222 82688 589228
rect 83476 589098 83504 592039
rect 83752 591025 83780 596146
rect 86224 593428 86276 593434
rect 86224 593370 86276 593376
rect 83738 591016 83794 591025
rect 83738 590951 83794 590960
rect 82248 589070 82584 589098
rect 83168 589070 83504 589098
rect 78416 588798 78568 588826
rect 75642 588775 75698 588784
rect 75656 588690 75684 588775
rect 69480 588668 69532 588674
rect 75656 588662 75808 588690
rect 69480 588610 69532 588616
rect 83752 588470 83780 590951
rect 84108 590776 84160 590782
rect 84108 590718 84160 590724
rect 84120 589274 84148 590718
rect 84074 589246 84148 589274
rect 84074 589084 84102 589246
rect 86236 589098 86264 593370
rect 86880 592034 86908 703530
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 89180 700330 89208 703520
rect 93768 703452 93820 703458
rect 93768 703394 93820 703400
rect 89812 702636 89864 702642
rect 89812 702578 89864 702584
rect 89168 700324 89220 700330
rect 89168 700266 89220 700272
rect 88984 700256 89036 700262
rect 88984 700198 89036 700204
rect 87604 605872 87656 605878
rect 87604 605814 87656 605820
rect 87616 594454 87644 605814
rect 88996 599622 89024 700198
rect 88984 599616 89036 599622
rect 88984 599558 89036 599564
rect 88892 598256 88944 598262
rect 88892 598198 88944 598204
rect 88904 596174 88932 598198
rect 88904 596146 89116 596174
rect 88984 595468 89036 595474
rect 88984 595410 89036 595416
rect 87604 594448 87656 594454
rect 87604 594390 87656 594396
rect 86880 592006 87092 592034
rect 86866 591016 86922 591025
rect 86866 590951 86922 590960
rect 86880 589274 86908 590951
rect 85928 589070 86264 589098
rect 86834 589246 86908 589274
rect 86960 589280 87012 589286
rect 86834 589084 86862 589246
rect 86960 589222 87012 589228
rect 86972 588849 87000 589222
rect 86958 588840 87014 588849
rect 86958 588775 87014 588784
rect 87064 588606 87092 592006
rect 88996 590617 89024 595410
rect 88982 590608 89038 590617
rect 88982 590543 89038 590552
rect 85304 588600 85356 588606
rect 85008 588548 85304 588554
rect 85008 588542 85356 588548
rect 87052 588600 87104 588606
rect 88062 588568 88118 588577
rect 87052 588542 87104 588548
rect 85008 588526 85344 588542
rect 87768 588526 88062 588554
rect 88062 588503 88118 588512
rect 83740 588464 83792 588470
rect 83740 588406 83792 588412
rect 88688 588390 89024 588418
rect 88892 588328 88944 588334
rect 88892 588270 88944 588276
rect 67730 585848 67786 585857
rect 67730 585783 67786 585792
rect 67744 585206 67772 585783
rect 67732 585200 67784 585206
rect 67732 585142 67784 585148
rect 88904 582374 88932 588270
rect 88996 583001 89024 588390
rect 88982 582992 89038 583001
rect 88982 582927 89038 582936
rect 88904 582346 89024 582374
rect 88996 581754 89024 582346
rect 88812 581726 89024 581754
rect 67730 578368 67786 578377
rect 67730 578303 67786 578312
rect 67638 558920 67694 558929
rect 67638 558855 67694 558864
rect 67652 557598 67680 558855
rect 67640 557592 67692 557598
rect 67640 557534 67692 557540
rect 67454 552256 67510 552265
rect 67454 552191 67510 552200
rect 67364 442944 67416 442950
rect 67364 442886 67416 442892
rect 66994 439920 67050 439929
rect 66994 439855 67050 439864
rect 67008 439074 67036 439855
rect 66996 439068 67048 439074
rect 66996 439010 67048 439016
rect 67364 439068 67416 439074
rect 67364 439010 67416 439016
rect 66904 419552 66956 419558
rect 66902 419520 66904 419529
rect 66956 419520 66958 419529
rect 66902 419455 66958 419464
rect 66444 418124 66496 418130
rect 66444 418066 66496 418072
rect 66456 417353 66484 418066
rect 66442 417344 66498 417353
rect 66442 417279 66498 417288
rect 66810 415168 66866 415177
rect 66810 415103 66866 415112
rect 66824 414730 66852 415103
rect 66812 414724 66864 414730
rect 66812 414666 66864 414672
rect 66258 406192 66314 406201
rect 66258 406127 66260 406136
rect 66312 406127 66314 406136
rect 66260 406098 66312 406104
rect 66258 403744 66314 403753
rect 66258 403679 66314 403688
rect 66272 403646 66300 403679
rect 66260 403640 66312 403646
rect 66260 403582 66312 403588
rect 66260 401600 66312 401606
rect 66258 401568 66260 401577
rect 66312 401568 66314 401577
rect 66258 401503 66314 401512
rect 66442 399392 66498 399401
rect 66442 399327 66498 399336
rect 66456 398138 66484 399327
rect 66444 398132 66496 398138
rect 66444 398074 66496 398080
rect 66994 396944 67050 396953
rect 66994 396879 67050 396888
rect 67008 396778 67036 396879
rect 66996 396772 67048 396778
rect 66996 396714 67048 396720
rect 67272 396772 67324 396778
rect 67272 396714 67324 396720
rect 66812 393304 66864 393310
rect 66812 393246 66864 393252
rect 66824 392601 66852 393246
rect 66810 392592 66866 392601
rect 66810 392527 66866 392536
rect 66166 388376 66222 388385
rect 66166 388311 66222 388320
rect 66074 360904 66130 360913
rect 66074 360839 66130 360848
rect 65616 353320 65668 353326
rect 65616 353262 65668 353268
rect 65628 321570 65656 353262
rect 66076 346452 66128 346458
rect 66076 346394 66128 346400
rect 65616 321564 65668 321570
rect 65616 321506 65668 321512
rect 66088 312089 66116 346394
rect 67284 345098 67312 396714
rect 67272 345092 67324 345098
rect 67272 345034 67324 345040
rect 66168 337476 66220 337482
rect 66168 337418 66220 337424
rect 66074 312080 66130 312089
rect 66074 312015 66130 312024
rect 64696 291168 64748 291174
rect 64696 291110 64748 291116
rect 65524 291168 65576 291174
rect 65524 291110 65576 291116
rect 64708 289950 64736 291110
rect 64696 289944 64748 289950
rect 64696 289886 64748 289892
rect 64512 269136 64564 269142
rect 64512 269078 64564 269084
rect 64524 240786 64552 269078
rect 64604 252680 64656 252686
rect 64604 252622 64656 252628
rect 64512 240780 64564 240786
rect 64512 240722 64564 240728
rect 64616 219337 64644 252622
rect 64708 234569 64736 289886
rect 66180 276185 66208 337418
rect 67178 326768 67234 326777
rect 67178 326703 67234 326712
rect 67192 325718 67220 326703
rect 67180 325712 67232 325718
rect 67180 325654 67232 325660
rect 66902 324864 66958 324873
rect 66902 324799 66958 324808
rect 66916 324358 66944 324799
rect 66904 324352 66956 324358
rect 66904 324294 66956 324300
rect 66810 323776 66866 323785
rect 66810 323711 66866 323720
rect 66824 322998 66852 323711
rect 66812 322992 66864 322998
rect 66812 322934 66864 322940
rect 66444 321564 66496 321570
rect 66444 321506 66496 321512
rect 66456 320521 66484 321506
rect 66442 320512 66498 320521
rect 66442 320447 66498 320456
rect 66810 319424 66866 319433
rect 66810 319359 66866 319368
rect 66824 318850 66852 319359
rect 66812 318844 66864 318850
rect 66812 318786 66864 318792
rect 66902 318336 66958 318345
rect 66902 318271 66958 318280
rect 66812 317552 66864 317558
rect 66810 317520 66812 317529
rect 66864 317520 66866 317529
rect 66916 317490 66944 318271
rect 66810 317455 66866 317464
rect 66904 317484 66956 317490
rect 66904 317426 66956 317432
rect 67284 316441 67312 345034
rect 67376 338473 67404 439010
rect 67468 412729 67496 552191
rect 67548 540932 67600 540938
rect 67548 540874 67600 540880
rect 67560 539646 67588 540874
rect 67548 539640 67600 539646
rect 67548 539582 67600 539588
rect 67548 539504 67600 539510
rect 67548 539446 67600 539452
rect 67454 412720 67510 412729
rect 67454 412655 67510 412664
rect 67362 338464 67418 338473
rect 67362 338399 67418 338408
rect 67376 327049 67404 338399
rect 67362 327040 67418 327049
rect 67362 326975 67418 326984
rect 67364 325644 67416 325650
rect 67364 325586 67416 325592
rect 67376 321609 67404 325586
rect 67362 321600 67418 321609
rect 67362 321535 67418 321544
rect 67364 320884 67416 320890
rect 67364 320826 67416 320832
rect 67270 316432 67326 316441
rect 67270 316367 67326 316376
rect 66812 315988 66864 315994
rect 66812 315930 66864 315936
rect 66824 315353 66852 315930
rect 66810 315344 66866 315353
rect 66810 315279 66866 315288
rect 66902 314256 66958 314265
rect 66902 314191 66958 314200
rect 66916 313342 66944 314191
rect 66904 313336 66956 313342
rect 66904 313278 66956 313284
rect 66812 313268 66864 313274
rect 66812 313210 66864 313216
rect 66824 313177 66852 313210
rect 66810 313168 66866 313177
rect 66810 313103 66866 313112
rect 66444 311840 66496 311846
rect 66444 311782 66496 311788
rect 66456 311001 66484 311782
rect 66442 310992 66498 311001
rect 66442 310927 66498 310936
rect 66810 309904 66866 309913
rect 66810 309839 66866 309848
rect 66824 309194 66852 309839
rect 66812 309188 66864 309194
rect 66812 309130 66864 309136
rect 66718 308000 66774 308009
rect 66718 307935 66774 307944
rect 66732 307086 66760 307935
rect 66720 307080 66772 307086
rect 66720 307022 66772 307028
rect 66996 306400 67048 306406
rect 66996 306342 67048 306348
rect 66904 306332 66956 306338
rect 66904 306274 66956 306280
rect 66916 305833 66944 306274
rect 66902 305824 66958 305833
rect 66902 305759 66958 305768
rect 66902 304736 66958 304745
rect 66902 304671 66958 304680
rect 66260 303680 66312 303686
rect 66258 303648 66260 303657
rect 66312 303648 66314 303657
rect 66258 303583 66314 303592
rect 66812 303612 66864 303618
rect 66812 303554 66864 303560
rect 66824 302569 66852 303554
rect 66810 302560 66866 302569
rect 66810 302495 66866 302504
rect 66812 302184 66864 302190
rect 66812 302126 66864 302132
rect 66824 301481 66852 302126
rect 66810 301472 66866 301481
rect 66810 301407 66866 301416
rect 66812 300824 66864 300830
rect 66812 300766 66864 300772
rect 66258 300656 66314 300665
rect 66258 300591 66314 300600
rect 66272 299606 66300 300591
rect 66260 299600 66312 299606
rect 66824 299577 66852 300766
rect 66260 299542 66312 299548
rect 66810 299568 66866 299577
rect 66810 299503 66866 299512
rect 66916 298790 66944 304671
rect 66904 298784 66956 298790
rect 66904 298726 66956 298732
rect 66444 296676 66496 296682
rect 66444 296618 66496 296624
rect 66456 296313 66484 296618
rect 66442 296304 66498 296313
rect 66442 296239 66498 296248
rect 66258 294128 66314 294137
rect 66258 294063 66260 294072
rect 66312 294063 66314 294072
rect 66260 294034 66312 294040
rect 66902 293040 66958 293049
rect 66902 292975 66958 292984
rect 66812 292528 66864 292534
rect 66812 292470 66864 292476
rect 66824 292233 66852 292470
rect 66810 292224 66866 292233
rect 66810 292159 66866 292168
rect 66810 290048 66866 290057
rect 66810 289983 66866 289992
rect 66824 289950 66852 289983
rect 66812 289944 66864 289950
rect 66812 289886 66864 289892
rect 66260 289264 66312 289270
rect 66260 289206 66312 289212
rect 66272 288969 66300 289206
rect 66258 288960 66314 288969
rect 66258 288895 66314 288904
rect 66810 287872 66866 287881
rect 66810 287807 66866 287816
rect 66824 287094 66852 287807
rect 66812 287088 66864 287094
rect 66812 287030 66864 287036
rect 66812 285728 66864 285734
rect 66810 285696 66812 285705
rect 66864 285696 66866 285705
rect 66810 285631 66866 285640
rect 66626 283792 66682 283801
rect 66626 283727 66682 283736
rect 66640 282946 66668 283727
rect 66628 282940 66680 282946
rect 66628 282882 66680 282888
rect 66350 282704 66406 282713
rect 66350 282639 66406 282648
rect 66364 281586 66392 282639
rect 66352 281580 66404 281586
rect 66352 281522 66404 281528
rect 66810 280528 66866 280537
rect 66810 280463 66866 280472
rect 66824 280226 66852 280463
rect 66812 280220 66864 280226
rect 66812 280162 66864 280168
rect 66626 279440 66682 279449
rect 66626 279375 66682 279384
rect 66640 278798 66668 279375
rect 66628 278792 66680 278798
rect 66628 278734 66680 278740
rect 66258 277264 66314 277273
rect 66258 277199 66314 277208
rect 66166 276176 66222 276185
rect 66166 276111 66222 276120
rect 65984 264240 66036 264246
rect 65984 264182 66036 264188
rect 65996 242078 66024 264182
rect 66074 256320 66130 256329
rect 66074 256255 66130 256264
rect 65984 242072 66036 242078
rect 65984 242014 66036 242020
rect 64694 234560 64750 234569
rect 64694 234495 64750 234504
rect 66088 229770 66116 256255
rect 66076 229764 66128 229770
rect 66076 229706 66128 229712
rect 64602 219328 64658 219337
rect 64602 219263 64658 219272
rect 66180 202881 66208 276111
rect 66272 273970 66300 277199
rect 66260 273964 66312 273970
rect 66260 273906 66312 273912
rect 66810 272096 66866 272105
rect 66810 272031 66866 272040
rect 66824 271930 66852 272031
rect 66812 271924 66864 271930
rect 66812 271866 66864 271872
rect 66810 271008 66866 271017
rect 66810 270943 66866 270952
rect 66824 270570 66852 270943
rect 66812 270564 66864 270570
rect 66812 270506 66864 270512
rect 66442 269920 66498 269929
rect 66442 269855 66498 269864
rect 66456 269142 66484 269855
rect 66444 269136 66496 269142
rect 66444 269078 66496 269084
rect 66442 267744 66498 267753
rect 66442 267679 66444 267688
rect 66496 267679 66498 267688
rect 66444 267650 66496 267656
rect 66916 267034 66944 292975
rect 67008 287054 67036 306342
rect 67008 287026 67128 287054
rect 66994 286784 67050 286793
rect 66994 286719 67050 286728
rect 67008 285802 67036 286719
rect 66996 285796 67048 285802
rect 66996 285738 67048 285744
rect 67100 284617 67128 287026
rect 67086 284608 67142 284617
rect 67086 284543 67142 284552
rect 67376 278361 67404 320826
rect 67468 309097 67496 412655
rect 67560 394777 67588 539446
rect 67640 533452 67692 533458
rect 67640 533394 67692 533400
rect 67546 394768 67602 394777
rect 67546 394703 67602 394712
rect 67560 372706 67588 394703
rect 67652 389094 67680 533394
rect 67744 476066 67772 578303
rect 67822 577008 67878 577017
rect 67822 576943 67878 576952
rect 67836 538966 67864 576943
rect 68652 540932 68704 540938
rect 68652 540874 68704 540880
rect 68664 540841 68692 540874
rect 68650 540832 68706 540841
rect 68650 540767 68706 540776
rect 69848 539640 69900 539646
rect 69848 539582 69900 539588
rect 68480 539158 68816 539186
rect 69676 539158 69736 539186
rect 67824 538960 67876 538966
rect 67824 538902 67876 538908
rect 68480 533458 68508 539158
rect 69676 536790 69704 539158
rect 69664 536784 69716 536790
rect 69664 536726 69716 536732
rect 69676 535537 69704 536726
rect 69662 535528 69718 535537
rect 69662 535463 69718 535472
rect 68468 533452 68520 533458
rect 68468 533394 68520 533400
rect 67732 476060 67784 476066
rect 67732 476002 67784 476008
rect 67824 475516 67876 475522
rect 67824 475458 67876 475464
rect 67836 445777 67864 475458
rect 69860 462330 69888 539582
rect 70656 539158 70716 539186
rect 70688 538218 70716 539158
rect 71240 539158 71576 539186
rect 72436 539158 72496 539186
rect 73172 539158 73416 539186
rect 74000 539158 74336 539186
rect 74644 539158 75256 539186
rect 76176 539158 76512 539186
rect 70676 538212 70728 538218
rect 70676 538154 70728 538160
rect 70688 535537 70716 538154
rect 70674 535528 70730 535537
rect 70674 535463 70730 535472
rect 71240 528554 71268 539158
rect 72436 537538 72464 539158
rect 72424 537532 72476 537538
rect 72424 537474 72476 537480
rect 70504 528526 71268 528554
rect 69020 462324 69072 462330
rect 69020 462266 69072 462272
rect 69848 462324 69900 462330
rect 69848 462266 69900 462272
rect 69032 460970 69060 462266
rect 69020 460964 69072 460970
rect 69072 460912 69888 460934
rect 69020 460906 69888 460912
rect 68376 447160 68428 447166
rect 68376 447102 68428 447108
rect 67822 445768 67878 445777
rect 67822 445703 67878 445712
rect 67732 442944 67784 442950
rect 67732 442886 67784 442892
rect 67744 442105 67772 442886
rect 68388 442270 68416 447102
rect 68466 445768 68522 445777
rect 68466 445703 68522 445712
rect 68480 444258 68508 445703
rect 69860 444394 69888 460906
rect 70504 456074 70532 528526
rect 70492 456068 70544 456074
rect 70492 456010 70544 456016
rect 71780 450560 71832 450566
rect 71780 450502 71832 450508
rect 71792 447273 71820 450502
rect 72436 448633 72464 537474
rect 73172 536110 73200 539158
rect 73160 536104 73212 536110
rect 73160 536046 73212 536052
rect 74000 535498 74028 539158
rect 73160 535492 73212 535498
rect 73160 535434 73212 535440
rect 73988 535492 74040 535498
rect 73988 535434 74040 535440
rect 73172 461650 73200 535434
rect 73160 461644 73212 461650
rect 73160 461586 73212 461592
rect 73160 454708 73212 454714
rect 73160 454650 73212 454656
rect 73172 454102 73200 454650
rect 73160 454096 73212 454102
rect 73160 454038 73212 454044
rect 72422 448624 72478 448633
rect 72422 448559 72478 448568
rect 71778 447264 71834 447273
rect 71778 447199 71834 447208
rect 71792 444530 71820 447199
rect 73172 444666 73200 454038
rect 74644 449206 74672 539158
rect 74724 538960 74776 538966
rect 74724 538902 74776 538908
rect 74736 451314 74764 538902
rect 76484 536761 76512 539158
rect 76760 539158 77096 539186
rect 77312 539158 78016 539186
rect 78784 539158 78936 539186
rect 79520 539158 79856 539186
rect 80776 539158 80836 539186
rect 76760 538121 76788 539158
rect 76746 538112 76802 538121
rect 76746 538047 76802 538056
rect 76470 536752 76526 536761
rect 76470 536687 76526 536696
rect 75918 535528 75974 535537
rect 75918 535463 75974 535472
rect 75932 468518 75960 535463
rect 76484 529242 76512 536687
rect 76760 535537 76788 538047
rect 76746 535528 76802 535537
rect 76746 535463 76802 535472
rect 76472 529236 76524 529242
rect 76472 529178 76524 529184
rect 76564 476060 76616 476066
rect 76564 476002 76616 476008
rect 75920 468512 75972 468518
rect 75920 468454 75972 468460
rect 74724 451308 74776 451314
rect 74724 451250 74776 451256
rect 74632 449200 74684 449206
rect 74632 449142 74684 449148
rect 73172 444638 73246 444666
rect 71746 444502 71820 444530
rect 69860 444366 70288 444394
rect 71746 444380 71774 444502
rect 73218 444380 73246 444638
rect 74736 444394 74764 451250
rect 76576 445806 76604 476002
rect 77312 446418 77340 539158
rect 78680 533452 78732 533458
rect 78680 533394 78732 533400
rect 77944 532024 77996 532030
rect 77944 531966 77996 531972
rect 77956 455394 77984 531966
rect 78692 471306 78720 533394
rect 78680 471300 78732 471306
rect 78680 471242 78732 471248
rect 78680 464364 78732 464370
rect 78680 464306 78732 464312
rect 77392 455388 77444 455394
rect 77392 455330 77444 455336
rect 77944 455388 77996 455394
rect 77944 455330 77996 455336
rect 77404 454170 77432 455330
rect 77392 454164 77444 454170
rect 77392 454106 77444 454112
rect 77300 446412 77352 446418
rect 77300 446354 77352 446360
rect 76564 445800 76616 445806
rect 76564 445742 76616 445748
rect 76576 444394 76604 445742
rect 74736 444366 74888 444394
rect 76360 444366 76604 444394
rect 77404 444394 77432 454106
rect 78692 445913 78720 464306
rect 78784 453354 78812 539158
rect 79520 533458 79548 539158
rect 80808 538286 80836 539158
rect 81452 539158 81696 539186
rect 82616 539158 82768 539186
rect 83536 539158 84148 539186
rect 84456 539158 84792 539186
rect 85376 539158 85528 539186
rect 86296 539158 86632 539186
rect 80336 538280 80388 538286
rect 80336 538222 80388 538228
rect 80796 538280 80848 538286
rect 80796 538222 80848 538228
rect 79508 533452 79560 533458
rect 79508 533394 79560 533400
rect 80348 528554 80376 538222
rect 80072 528526 80376 528554
rect 80072 457502 80100 528526
rect 81452 461553 81480 539158
rect 82740 536790 82768 539158
rect 82728 536784 82780 536790
rect 82728 536726 82780 536732
rect 81438 461544 81494 461553
rect 81438 461479 81494 461488
rect 80060 457496 80112 457502
rect 80060 457438 80112 457444
rect 82082 457464 82138 457473
rect 82082 457399 82138 457408
rect 78772 453348 78824 453354
rect 78772 453290 78824 453296
rect 80888 449880 80940 449886
rect 80888 449822 80940 449828
rect 78678 445904 78734 445913
rect 78678 445839 78734 445848
rect 78692 444394 78720 445839
rect 80900 444530 80928 449822
rect 82096 445913 82124 457399
rect 82740 456249 82768 536726
rect 82820 460216 82872 460222
rect 84120 460193 84148 539158
rect 84764 536081 84792 539158
rect 85500 536246 85528 539158
rect 86604 538214 86632 539158
rect 87064 539158 87400 539186
rect 88320 539158 88656 539186
rect 86868 538214 86920 538218
rect 86604 538212 86920 538214
rect 86604 538186 86868 538212
rect 86868 538154 86920 538160
rect 85488 536240 85540 536246
rect 85488 536182 85540 536188
rect 86224 536240 86276 536246
rect 86224 536182 86276 536188
rect 84750 536072 84806 536081
rect 84750 536007 84806 536016
rect 85580 463004 85632 463010
rect 85580 462946 85632 462952
rect 82820 460158 82872 460164
rect 84106 460184 84162 460193
rect 82726 456240 82782 456249
rect 82726 456175 82782 456184
rect 82832 452742 82860 460158
rect 84106 460119 84162 460128
rect 82820 452736 82872 452742
rect 82820 452678 82872 452684
rect 83464 452736 83516 452742
rect 83464 452678 83516 452684
rect 82082 445904 82138 445913
rect 82082 445839 82138 445848
rect 80900 444502 80974 444530
rect 77404 444366 77832 444394
rect 78692 444366 79488 444394
rect 80946 444380 80974 444502
rect 82096 444394 82124 445839
rect 83476 444394 83504 452678
rect 85592 446049 85620 462946
rect 86236 449177 86264 536182
rect 86880 462913 86908 538154
rect 86866 462904 86922 462913
rect 86866 462839 86922 462848
rect 86960 458244 87012 458250
rect 86960 458186 87012 458192
rect 86222 449168 86278 449177
rect 86222 449103 86278 449112
rect 85578 446040 85634 446049
rect 85578 445975 85634 445984
rect 85592 444666 85620 445975
rect 85546 444638 85620 444666
rect 86972 444666 87000 458186
rect 87064 457473 87092 539158
rect 88628 535498 88656 539158
rect 88616 535492 88668 535498
rect 88616 535434 88668 535440
rect 87050 457464 87106 457473
rect 87050 457399 87106 457408
rect 88812 447166 88840 581726
rect 89088 576858 89116 596146
rect 89720 589960 89772 589966
rect 89720 589902 89772 589908
rect 88904 576830 89116 576858
rect 88904 567293 88932 576830
rect 88890 567284 88946 567293
rect 88890 567219 88892 567228
rect 88944 567219 88946 567228
rect 88892 567190 88944 567196
rect 89536 539572 89588 539578
rect 89536 539514 89588 539520
rect 89548 538354 89576 539514
rect 89536 538348 89588 538354
rect 89536 538290 89588 538296
rect 89548 465798 89576 538290
rect 89628 535492 89680 535498
rect 89628 535434 89680 535440
rect 89536 465792 89588 465798
rect 89536 465734 89588 465740
rect 89640 456113 89668 535434
rect 89626 456104 89682 456113
rect 89626 456039 89682 456048
rect 88800 447160 88852 447166
rect 88800 447102 88852 447108
rect 86972 444638 87046 444666
rect 82096 444366 82432 444394
rect 83476 444366 83904 444394
rect 85546 444380 85574 444638
rect 87018 444380 87046 444638
rect 88812 444394 88840 447102
rect 88504 444366 88840 444394
rect 89732 444394 89760 589902
rect 89824 560153 89852 702578
rect 91192 594448 91244 594454
rect 91192 594390 91244 594396
rect 89902 585848 89958 585857
rect 89902 585783 89958 585792
rect 89810 560144 89866 560153
rect 89810 560079 89866 560088
rect 89916 539578 89944 585783
rect 91098 581632 91154 581641
rect 91098 581567 91154 581576
rect 91112 581058 91140 581567
rect 91100 581052 91152 581058
rect 91100 580994 91152 581000
rect 91098 578912 91154 578921
rect 91098 578847 91154 578856
rect 91112 578270 91140 578847
rect 91100 578264 91152 578270
rect 91100 578206 91152 578212
rect 91098 577552 91154 577561
rect 91098 577487 91154 577496
rect 91112 576910 91140 577487
rect 91100 576904 91152 576910
rect 91100 576846 91152 576852
rect 91204 576745 91232 594390
rect 92480 587852 92532 587858
rect 92480 587794 92532 587800
rect 91926 584624 91982 584633
rect 91926 584559 91982 584568
rect 91940 584458 91968 584559
rect 91928 584452 91980 584458
rect 91928 584394 91980 584400
rect 91836 583704 91888 583710
rect 91834 583672 91836 583681
rect 91888 583672 91890 583681
rect 91834 583607 91890 583616
rect 91190 576736 91246 576745
rect 91190 576671 91246 576680
rect 91204 576162 91232 576671
rect 91192 576156 91244 576162
rect 91192 576098 91244 576104
rect 91098 575104 91154 575113
rect 91098 575039 91154 575048
rect 91112 574802 91140 575039
rect 91100 574796 91152 574802
rect 91100 574738 91152 574744
rect 91098 573472 91154 573481
rect 91098 573407 91154 573416
rect 91112 572762 91140 573407
rect 91100 572756 91152 572762
rect 91100 572698 91152 572704
rect 91190 572112 91246 572121
rect 91190 572047 91246 572056
rect 91204 571470 91232 572047
rect 91192 571464 91244 571470
rect 91098 571432 91154 571441
rect 91192 571406 91244 571412
rect 91098 571367 91100 571376
rect 91152 571367 91154 571376
rect 91100 571338 91152 571344
rect 91098 570072 91154 570081
rect 91098 570007 91154 570016
rect 91112 569974 91140 570007
rect 91100 569968 91152 569974
rect 91100 569910 91152 569916
rect 92202 568712 92258 568721
rect 92202 568647 92258 568656
rect 91100 565888 91152 565894
rect 91098 565856 91100 565865
rect 91152 565856 91154 565865
rect 91098 565791 91154 565800
rect 91742 564496 91798 564505
rect 91742 564431 91798 564440
rect 91098 563136 91154 563145
rect 91098 563071 91100 563080
rect 91152 563071 91154 563080
rect 91100 563042 91152 563048
rect 91098 560960 91154 560969
rect 91098 560895 91154 560904
rect 89996 546440 90048 546446
rect 89996 546382 90048 546388
rect 91008 546440 91060 546446
rect 91008 546382 91060 546388
rect 90008 545329 90036 546382
rect 89994 545320 90050 545329
rect 89994 545255 90050 545264
rect 89904 539572 89956 539578
rect 89904 539514 89956 539520
rect 91020 458833 91048 546382
rect 91112 530602 91140 560895
rect 91190 558240 91246 558249
rect 91190 558175 91246 558184
rect 91204 557598 91232 558175
rect 91192 557592 91244 557598
rect 91192 557534 91244 557540
rect 91190 556880 91246 556889
rect 91190 556815 91246 556824
rect 91204 556238 91232 556815
rect 91192 556232 91244 556238
rect 91192 556174 91244 556180
rect 91190 555520 91246 555529
rect 91190 555455 91246 555464
rect 91204 554810 91232 555455
rect 91192 554804 91244 554810
rect 91192 554746 91244 554752
rect 91190 552936 91246 552945
rect 91190 552871 91246 552880
rect 91204 552362 91232 552871
rect 91192 552356 91244 552362
rect 91192 552298 91244 552304
rect 91190 552120 91246 552129
rect 91190 552055 91192 552064
rect 91244 552055 91246 552064
rect 91192 552026 91244 552032
rect 91190 549400 91246 549409
rect 91190 549335 91246 549344
rect 91204 549302 91232 549335
rect 91192 549296 91244 549302
rect 91192 549238 91244 549244
rect 91282 547904 91338 547913
rect 91282 547839 91338 547848
rect 91192 544400 91244 544406
rect 91192 544342 91244 544348
rect 91204 544105 91232 544342
rect 91190 544096 91246 544105
rect 91190 544031 91246 544040
rect 91190 542464 91246 542473
rect 91190 542399 91192 542408
rect 91244 542399 91246 542408
rect 91192 542370 91244 542376
rect 91192 541680 91244 541686
rect 91192 541622 91244 541628
rect 91204 541385 91232 541622
rect 91190 541376 91246 541385
rect 91190 541311 91246 541320
rect 91190 539744 91246 539753
rect 91190 539679 91192 539688
rect 91244 539679 91246 539688
rect 91192 539650 91244 539656
rect 91296 534750 91324 547839
rect 91374 546544 91430 546553
rect 91374 546479 91430 546488
rect 91284 534744 91336 534750
rect 91284 534686 91336 534692
rect 91388 533390 91416 546479
rect 91376 533384 91428 533390
rect 91376 533326 91428 533332
rect 91100 530596 91152 530602
rect 91100 530538 91152 530544
rect 91006 458824 91062 458833
rect 91006 458759 91062 458768
rect 91560 451920 91612 451926
rect 91756 451897 91784 564431
rect 92216 562358 92244 568647
rect 92204 562352 92256 562358
rect 92204 562294 92256 562300
rect 91834 560144 91890 560153
rect 91834 560079 91890 560088
rect 91848 548554 91876 560079
rect 91836 548548 91888 548554
rect 91836 548490 91888 548496
rect 91560 451862 91612 451868
rect 91742 451888 91798 451897
rect 91572 448633 91600 451862
rect 91742 451823 91798 451832
rect 91558 448624 91614 448633
rect 91558 448559 91614 448568
rect 91572 444666 91600 448559
rect 91572 444638 91646 444666
rect 90132 444544 90188 444553
rect 90132 444479 90188 444488
rect 90146 444394 90174 444479
rect 89732 444380 90174 444394
rect 91618 444380 91646 444638
rect 92492 444514 92520 587794
rect 93780 584458 93808 703394
rect 98736 703112 98788 703118
rect 98736 703054 98788 703060
rect 97908 702772 97960 702778
rect 97908 702714 97960 702720
rect 94504 702636 94556 702642
rect 94504 702578 94556 702584
rect 93860 589416 93912 589422
rect 93860 589358 93912 589364
rect 93768 584452 93820 584458
rect 93768 584394 93820 584400
rect 93768 583704 93820 583710
rect 93768 583646 93820 583652
rect 93124 539708 93176 539714
rect 93124 539650 93176 539656
rect 93136 460193 93164 539650
rect 93780 469849 93808 583646
rect 93766 469840 93822 469849
rect 93766 469775 93822 469784
rect 93122 460184 93178 460193
rect 93122 460119 93178 460128
rect 93872 445777 93900 589358
rect 94516 583710 94544 702578
rect 96620 592136 96672 592142
rect 96620 592078 96672 592084
rect 95884 590776 95936 590782
rect 95884 590718 95936 590724
rect 94504 583704 94556 583710
rect 94504 583646 94556 583652
rect 95148 574796 95200 574802
rect 95148 574738 95200 574744
rect 95160 558210 95188 574738
rect 95896 565146 95924 590718
rect 95884 565140 95936 565146
rect 95884 565082 95936 565088
rect 95148 558204 95200 558210
rect 95148 558146 95200 558152
rect 95240 552356 95292 552362
rect 95240 552298 95292 552304
rect 95148 544400 95200 544406
rect 95148 544342 95200 544348
rect 95160 467129 95188 544342
rect 95146 467120 95202 467129
rect 95146 467055 95202 467064
rect 95252 446457 95280 552298
rect 95884 465724 95936 465730
rect 95884 465666 95936 465672
rect 95896 455569 95924 465666
rect 95882 455560 95938 455569
rect 95882 455495 95938 455504
rect 95896 451274 95924 455495
rect 95804 451246 95924 451274
rect 95238 446448 95294 446457
rect 95238 446383 95294 446392
rect 93858 445768 93914 445777
rect 93858 445703 93914 445712
rect 94502 445768 94558 445777
rect 94502 445703 94558 445712
rect 92480 444508 92532 444514
rect 92480 444450 92532 444456
rect 93078 444508 93130 444514
rect 93078 444450 93130 444456
rect 93090 444380 93118 444450
rect 94516 444394 94544 445703
rect 95804 444394 95832 451246
rect 96632 445777 96660 592078
rect 97920 580961 97948 702714
rect 98642 588704 98698 588713
rect 98642 588639 98698 588648
rect 97906 580952 97962 580961
rect 97906 580887 97962 580896
rect 97920 580281 97948 580887
rect 97906 580272 97962 580281
rect 97906 580207 97962 580216
rect 98656 451314 98684 588639
rect 98748 574802 98776 703054
rect 105464 700330 105492 703520
rect 130384 703248 130436 703254
rect 130384 703190 130436 703196
rect 124864 703044 124916 703050
rect 124864 702986 124916 702992
rect 105452 700324 105504 700330
rect 105452 700266 105504 700272
rect 114560 599004 114612 599010
rect 114560 598946 114612 598952
rect 108304 595468 108356 595474
rect 108304 595410 108356 595416
rect 105544 594856 105596 594862
rect 105544 594798 105596 594804
rect 102140 592068 102192 592074
rect 102140 592010 102192 592016
rect 100760 590708 100812 590714
rect 100760 590650 100812 590656
rect 100772 588198 100800 590650
rect 101402 588840 101458 588849
rect 101402 588775 101458 588784
rect 100760 588192 100812 588198
rect 100760 588134 100812 588140
rect 98736 574796 98788 574802
rect 98736 574738 98788 574744
rect 100668 554804 100720 554810
rect 100668 554746 100720 554752
rect 98736 549296 98788 549302
rect 98736 549238 98788 549244
rect 98748 461553 98776 549238
rect 100680 462913 100708 554746
rect 100666 462904 100722 462913
rect 100666 462839 100722 462848
rect 98734 461544 98790 461553
rect 98734 461479 98790 461488
rect 98644 451308 98696 451314
rect 98644 451250 98696 451256
rect 96618 445768 96674 445777
rect 96618 445703 96674 445712
rect 97354 445768 97410 445777
rect 97354 445703 97410 445712
rect 97368 444394 97396 445703
rect 98656 444394 98684 451250
rect 101416 444514 101444 588775
rect 102152 445777 102180 592010
rect 103520 588192 103572 588198
rect 103520 588134 103572 588140
rect 103532 451246 103560 588134
rect 104164 581052 104216 581058
rect 104164 580994 104216 581000
rect 103520 451240 103572 451246
rect 103520 451182 103572 451188
rect 104176 450537 104204 580994
rect 104256 542428 104308 542434
rect 104256 542370 104308 542376
rect 104268 459649 104296 542370
rect 104254 459640 104310 459649
rect 104254 459575 104310 459584
rect 104624 451240 104676 451246
rect 104624 451182 104676 451188
rect 104162 450528 104218 450537
rect 104162 450463 104218 450472
rect 104636 450022 104664 451182
rect 104072 450016 104124 450022
rect 104072 449958 104124 449964
rect 104624 450016 104676 450022
rect 104624 449958 104676 449964
rect 102138 445768 102194 445777
rect 102138 445703 102194 445712
rect 101404 444508 101456 444514
rect 101404 444450 101456 444456
rect 101416 444394 101444 444450
rect 89732 444366 90160 444380
rect 94516 444366 94760 444394
rect 95804 444366 96232 444394
rect 97368 444366 97704 444394
rect 98656 444366 99176 444394
rect 100832 444366 101444 444394
rect 102152 444394 102180 445703
rect 104084 444394 104112 449958
rect 105556 446049 105584 594798
rect 107014 590880 107070 590889
rect 107014 590815 107070 590824
rect 105636 576156 105688 576162
rect 105636 576098 105688 576104
rect 105648 447846 105676 576098
rect 107028 553110 107056 590815
rect 107016 553104 107068 553110
rect 107016 553046 107068 553052
rect 106924 552084 106976 552090
rect 106924 552026 106976 552032
rect 106280 458856 106332 458862
rect 106280 458798 106332 458804
rect 105636 447840 105688 447846
rect 105636 447782 105688 447788
rect 105542 446040 105598 446049
rect 105542 445975 105598 445984
rect 105556 444394 105584 445975
rect 102152 444366 102304 444394
rect 103776 444366 104112 444394
rect 105432 444366 105584 444394
rect 106292 444394 106320 458798
rect 106936 456113 106964 552026
rect 106922 456104 106978 456113
rect 106922 456039 106978 456048
rect 108316 448594 108344 595410
rect 110418 592104 110474 592113
rect 110418 592039 110474 592048
rect 108396 571464 108448 571470
rect 108396 571406 108448 571412
rect 108304 448588 108356 448594
rect 108304 448530 108356 448536
rect 108316 444666 108344 448530
rect 108408 447817 108436 571406
rect 109040 553104 109092 553110
rect 109040 553046 109092 553052
rect 108394 447808 108450 447817
rect 108394 447743 108450 447752
rect 109052 444689 109080 553046
rect 110432 445777 110460 592039
rect 112442 591016 112498 591025
rect 112442 590951 112498 590960
rect 111800 565140 111852 565146
rect 111800 565082 111852 565088
rect 111812 448526 111840 565082
rect 112456 458930 112484 590951
rect 113180 588600 113232 588606
rect 113180 588542 113232 588548
rect 112444 458924 112496 458930
rect 112444 458866 112496 458872
rect 111800 448520 111852 448526
rect 111800 448462 111852 448468
rect 111812 445874 111840 448462
rect 111800 445868 111852 445874
rect 111800 445810 111852 445816
rect 112996 445868 113048 445874
rect 112996 445810 113048 445816
rect 110418 445768 110474 445777
rect 110418 445703 110474 445712
rect 111154 445768 111210 445777
rect 111154 445703 111210 445712
rect 109038 444680 109094 444689
rect 108316 444638 108390 444666
rect 106292 444366 106904 444394
rect 108362 444380 108390 444638
rect 109038 444615 109094 444624
rect 109052 444394 109080 444615
rect 111168 444394 111196 445703
rect 113008 444530 113036 445810
rect 113192 445777 113220 588542
rect 114572 458862 114600 598946
rect 118698 585712 118754 585721
rect 118698 585647 118754 585656
rect 116584 569968 116636 569974
rect 116584 569910 116636 569916
rect 114560 458856 114612 458862
rect 114560 458798 114612 458804
rect 116596 449206 116624 569910
rect 117320 458924 117372 458930
rect 117320 458866 117372 458872
rect 116584 449200 116636 449206
rect 116584 449142 116636 449148
rect 116398 445904 116454 445913
rect 116398 445839 116454 445848
rect 113178 445768 113234 445777
rect 113178 445703 113234 445712
rect 114098 445768 114154 445777
rect 114098 445703 114154 445712
rect 112962 444502 113036 444530
rect 109052 444366 109848 444394
rect 111168 444366 111504 444394
rect 112962 444380 112990 444502
rect 114112 444394 114140 445703
rect 116412 444394 116440 445839
rect 117332 445777 117360 458866
rect 117318 445768 117374 445777
rect 117318 445703 117374 445712
rect 114112 444366 114448 444394
rect 116104 444366 116440 444394
rect 117332 444394 117360 445703
rect 118712 444446 118740 585647
rect 124220 584452 124272 584458
rect 124220 584394 124272 584400
rect 123482 582992 123538 583001
rect 123482 582927 123538 582936
rect 121644 578264 121696 578270
rect 121644 578206 121696 578212
rect 120632 572756 120684 572762
rect 120632 572698 120684 572704
rect 119020 444680 119076 444689
rect 119020 444615 119076 444624
rect 118700 444440 118752 444446
rect 117332 444366 117576 444394
rect 119034 444394 119062 444615
rect 118752 444388 119062 444394
rect 118700 444382 119062 444388
rect 118712 444380 119062 444382
rect 118712 444366 119048 444380
rect 68650 444272 68706 444281
rect 68480 444230 68650 444258
rect 68706 444230 68816 444258
rect 68650 444207 68706 444216
rect 68664 444147 68692 444207
rect 68376 442264 68428 442270
rect 68376 442206 68428 442212
rect 67730 442096 67786 442105
rect 67730 442031 67786 442040
rect 67640 389088 67692 389094
rect 67640 389030 67692 389036
rect 67548 372700 67600 372706
rect 67548 372642 67600 372648
rect 67454 309088 67510 309097
rect 67454 309023 67510 309032
rect 67560 298489 67588 372642
rect 67652 353326 67680 389030
rect 67744 380186 67772 442031
rect 120644 419393 120672 572698
rect 120724 562352 120776 562358
rect 120724 562294 120776 562300
rect 120630 419384 120686 419393
rect 120630 419319 120686 419328
rect 120630 416800 120686 416809
rect 120630 416735 120686 416744
rect 67822 410544 67878 410553
rect 67822 410479 67878 410488
rect 67836 389881 67864 410479
rect 68376 408468 68428 408474
rect 68376 408410 68428 408416
rect 68388 408377 68416 408410
rect 68374 408368 68430 408377
rect 68374 408303 68430 408312
rect 81440 390992 81492 390998
rect 81440 390934 81492 390940
rect 82084 390992 82136 390998
rect 92754 390960 92810 390969
rect 82136 390940 82432 390946
rect 82084 390934 82432 390940
rect 73232 390646 73384 390674
rect 69938 390416 69994 390425
rect 68480 390374 68816 390402
rect 67822 389872 67878 389881
rect 67822 389807 67878 389816
rect 68480 389094 68508 390374
rect 71870 390416 71926 390425
rect 69994 390388 70288 390402
rect 69994 390374 70302 390388
rect 71760 390374 71870 390402
rect 69938 390351 69994 390360
rect 70274 390130 70302 390374
rect 71926 390374 72096 390402
rect 71870 390351 71926 390360
rect 71884 390291 71912 390351
rect 70274 390102 70348 390130
rect 68468 389088 68520 389094
rect 68468 389030 68520 389036
rect 67732 380180 67784 380186
rect 67732 380122 67784 380128
rect 70320 374678 70348 390102
rect 72068 389065 72096 390374
rect 72054 389056 72110 389065
rect 72054 388991 72110 389000
rect 73066 389056 73122 389065
rect 73356 389026 73384 390646
rect 74552 390374 74888 390402
rect 76360 390374 76696 390402
rect 77832 390374 77984 390402
rect 73066 388991 73122 389000
rect 73160 389020 73212 389026
rect 70308 374672 70360 374678
rect 70308 374614 70360 374620
rect 71688 374264 71740 374270
rect 71688 374206 71740 374212
rect 71596 359508 71648 359514
rect 71596 359450 71648 359456
rect 70400 356788 70452 356794
rect 70400 356730 70452 356736
rect 67640 353320 67692 353326
rect 67640 353262 67692 353268
rect 69848 353320 69900 353326
rect 69848 353262 69900 353268
rect 67640 342304 67692 342310
rect 67640 342246 67692 342252
rect 67652 322697 67680 342246
rect 69860 335354 69888 353262
rect 70306 347984 70362 347993
rect 70306 347919 70362 347928
rect 70320 335354 70348 347919
rect 70412 345014 70440 356730
rect 71608 349858 71636 359450
rect 71700 356794 71728 374206
rect 71688 356788 71740 356794
rect 71688 356730 71740 356736
rect 71700 356114 71728 356730
rect 71688 356108 71740 356114
rect 71688 356050 71740 356056
rect 71596 349852 71648 349858
rect 71596 349794 71648 349800
rect 70412 344986 70808 345014
rect 69584 335326 69888 335354
rect 70136 335326 70348 335354
rect 69386 331256 69442 331265
rect 69386 331191 69442 331200
rect 68282 329080 68338 329089
rect 68282 329015 68338 329024
rect 67824 328432 67876 328438
rect 67824 328374 67876 328380
rect 67732 326936 67784 326942
rect 67732 326878 67784 326884
rect 67744 325650 67772 326878
rect 67732 325644 67784 325650
rect 67732 325586 67784 325592
rect 67638 322688 67694 322697
rect 67638 322623 67694 322632
rect 67836 316034 67864 328374
rect 68296 320890 68324 329015
rect 68650 327176 68706 327185
rect 68706 327134 69000 327162
rect 68650 327111 68706 327120
rect 68652 327072 68704 327078
rect 68652 327014 68704 327020
rect 68560 327004 68612 327010
rect 68560 326946 68612 326952
rect 68572 326505 68600 326946
rect 68558 326496 68614 326505
rect 68558 326431 68614 326440
rect 68664 326233 68692 327014
rect 69400 327010 69428 331191
rect 69388 327004 69440 327010
rect 69388 326946 69440 326952
rect 69584 326942 69612 335326
rect 70136 327570 70164 335326
rect 70674 332616 70730 332625
rect 70674 332551 70730 332560
rect 70688 327570 70716 332551
rect 69736 327542 70164 327570
rect 70472 327542 70716 327570
rect 70780 327570 70808 344986
rect 71780 338156 71832 338162
rect 71780 338098 71832 338104
rect 71792 327570 71820 338098
rect 72974 334248 73030 334257
rect 72974 334183 73030 334192
rect 71872 332648 71924 332654
rect 71872 332590 71924 332596
rect 71884 328438 71912 332590
rect 71872 328432 71924 328438
rect 71872 328374 71924 328380
rect 72988 327570 73016 334183
rect 73080 332654 73108 388991
rect 73160 388962 73212 388968
rect 73344 389020 73396 389026
rect 73344 388962 73396 388968
rect 73172 374270 73200 388962
rect 74552 388929 74580 390374
rect 76668 389162 76696 390374
rect 76656 389156 76708 389162
rect 76656 389098 76708 389104
rect 74538 388920 74594 388929
rect 74538 388855 74594 388864
rect 73160 374264 73212 374270
rect 73160 374206 73212 374212
rect 73160 369912 73212 369918
rect 73160 369854 73212 369860
rect 73068 332648 73120 332654
rect 73068 332590 73120 332596
rect 70780 327542 71208 327570
rect 71792 327542 71944 327570
rect 72680 327542 73016 327570
rect 73172 327570 73200 369854
rect 74356 340196 74408 340202
rect 74356 340138 74408 340144
rect 74368 327570 74396 340138
rect 74552 337482 74580 388855
rect 76562 387152 76618 387161
rect 76562 387087 76618 387096
rect 75920 378820 75972 378826
rect 75920 378762 75972 378768
rect 74998 341456 75054 341465
rect 74998 341391 75054 341400
rect 74540 337476 74592 337482
rect 74540 337418 74592 337424
rect 74540 329860 74592 329866
rect 74540 329802 74592 329808
rect 73172 327542 73416 327570
rect 73968 327542 74396 327570
rect 74552 327434 74580 329802
rect 75012 327570 75040 341391
rect 75932 327570 75960 378762
rect 75012 327556 75440 327570
rect 75012 327542 75454 327556
rect 75932 327542 76512 327570
rect 74552 327406 74704 327434
rect 75426 327162 75454 327542
rect 76484 327214 76512 327542
rect 76472 327208 76524 327214
rect 75734 327176 75790 327185
rect 75426 327148 75734 327162
rect 75440 327134 75734 327148
rect 76472 327150 76524 327156
rect 75734 327111 75790 327120
rect 70030 327040 70086 327049
rect 76576 327010 76604 387087
rect 76668 366353 76696 389098
rect 77956 386374 77984 390374
rect 79336 390374 79488 390402
rect 80624 390374 80960 390402
rect 79336 387802 79364 390374
rect 79966 388376 80022 388385
rect 79966 388311 80022 388320
rect 79980 387870 80008 388311
rect 80624 387870 80652 390374
rect 79968 387864 80020 387870
rect 79968 387806 80020 387812
rect 80612 387864 80664 387870
rect 80612 387806 80664 387812
rect 79324 387796 79376 387802
rect 79324 387738 79376 387744
rect 77944 386368 77996 386374
rect 77944 386310 77996 386316
rect 76654 366344 76710 366353
rect 76654 366279 76710 366288
rect 77956 355473 77984 386310
rect 78680 370524 78732 370530
rect 78680 370466 78732 370472
rect 78692 365770 78720 370466
rect 78680 365764 78732 365770
rect 78680 365706 78732 365712
rect 77942 355464 77998 355473
rect 77942 355399 77998 355408
rect 78588 347064 78640 347070
rect 78588 347006 78640 347012
rect 77206 342408 77262 342417
rect 77206 342343 77262 342352
rect 77220 327570 77248 342343
rect 78600 327570 78628 347006
rect 78692 331158 78720 365706
rect 79336 365022 79364 387738
rect 79980 370530 80008 387806
rect 81452 371278 81480 390934
rect 82096 390918 82432 390934
rect 102598 390960 102654 390969
rect 92810 390918 93440 390946
rect 102304 390918 102598 390946
rect 92754 390895 92810 390904
rect 89810 390416 89866 390425
rect 82832 390374 83904 390402
rect 82832 383654 82860 390374
rect 85546 390130 85574 390388
rect 87018 390130 87046 390388
rect 88504 390374 89024 390402
rect 85546 390102 85620 390130
rect 85488 389836 85540 389842
rect 85488 389778 85540 389784
rect 85500 389065 85528 389778
rect 85486 389056 85542 389065
rect 85486 388991 85542 389000
rect 85592 386306 85620 390102
rect 86972 390102 87046 390130
rect 86972 389230 87000 390102
rect 86960 389224 87012 389230
rect 86960 389166 87012 389172
rect 85580 386300 85632 386306
rect 85580 386242 85632 386248
rect 82820 383648 82872 383654
rect 82820 383590 82872 383596
rect 81440 371272 81492 371278
rect 81440 371214 81492 371220
rect 79968 370524 80020 370530
rect 79968 370466 80020 370472
rect 81346 369064 81402 369073
rect 81346 368999 81402 369008
rect 79966 367704 80022 367713
rect 79966 367639 80022 367648
rect 79324 365016 79376 365022
rect 79324 364958 79376 364964
rect 79980 361622 80008 367639
rect 81360 362982 81388 368999
rect 80060 362976 80112 362982
rect 80060 362918 80112 362924
rect 81348 362976 81400 362982
rect 81348 362918 81400 362924
rect 78772 361616 78824 361622
rect 78772 361558 78824 361564
rect 79968 361616 80020 361622
rect 79968 361558 80020 361564
rect 78680 331152 78732 331158
rect 78680 331094 78732 331100
rect 76912 327542 77248 327570
rect 78384 327542 78628 327570
rect 78784 327570 78812 361558
rect 79324 331152 79376 331158
rect 79324 331094 79376 331100
rect 79336 327570 79364 331094
rect 80072 327570 80100 362918
rect 80702 339552 80758 339561
rect 80702 339487 80758 339496
rect 80716 327570 80744 339487
rect 81452 327570 81480 371214
rect 82832 344350 82860 383590
rect 84014 383072 84070 383081
rect 84014 383007 84070 383016
rect 84028 353569 84056 383007
rect 84106 374640 84162 374649
rect 84106 374575 84162 374584
rect 83462 353560 83518 353569
rect 83462 353495 83518 353504
rect 84014 353560 84070 353569
rect 84014 353495 84070 353504
rect 82820 344344 82872 344350
rect 82820 344286 82872 344292
rect 83476 331158 83504 353495
rect 82728 331152 82780 331158
rect 82728 331094 82780 331100
rect 83464 331152 83516 331158
rect 83464 331094 83516 331100
rect 82740 327570 82768 331094
rect 84120 330585 84148 374575
rect 85592 351121 85620 386242
rect 85762 352608 85818 352617
rect 85762 352543 85818 352552
rect 85578 351112 85634 351121
rect 85578 351047 85634 351056
rect 85488 350600 85540 350606
rect 85488 350542 85540 350548
rect 85500 335354 85528 350542
rect 85776 345137 85804 352543
rect 85762 345128 85818 345137
rect 85762 345063 85818 345072
rect 85776 345014 85804 345063
rect 85776 344986 86448 345014
rect 85224 335326 85528 335354
rect 84106 330576 84162 330585
rect 84106 330511 84162 330520
rect 83646 327720 83702 327729
rect 83646 327655 83702 327664
rect 83660 327570 83688 327655
rect 85224 327570 85252 335326
rect 86314 333296 86370 333305
rect 86314 333231 86370 333240
rect 85856 330540 85908 330546
rect 85856 330482 85908 330488
rect 85868 327570 85896 330482
rect 86328 327570 86356 333231
rect 78784 327542 79120 327570
rect 79336 327542 79672 327570
rect 80072 327542 80408 327570
rect 80716 327542 81144 327570
rect 81452 327542 81880 327570
rect 82616 327542 82768 327570
rect 83352 327542 83688 327570
rect 84824 327542 85252 327570
rect 85560 327542 85896 327570
rect 86112 327542 86356 327570
rect 86420 327570 86448 344986
rect 86972 337414 87000 389166
rect 88996 385014 89024 390374
rect 91282 390416 91338 390425
rect 89866 390374 90404 390402
rect 89810 390351 89866 390360
rect 90376 389065 90404 390374
rect 91338 390374 92060 390402
rect 91282 390351 91338 390360
rect 90362 389056 90418 389065
rect 90362 388991 90418 389000
rect 88984 385008 89036 385014
rect 88984 384950 89036 384956
rect 88996 352617 89024 384950
rect 89626 358864 89682 358873
rect 89626 358799 89682 358808
rect 88982 352608 89038 352617
rect 88982 352543 89038 352552
rect 89442 338328 89498 338337
rect 89442 338263 89498 338272
rect 86960 337408 87012 337414
rect 86960 337350 87012 337356
rect 87142 336832 87198 336841
rect 87142 336767 87198 336776
rect 87156 327570 87184 336767
rect 88616 329996 88668 330002
rect 88616 329938 88668 329944
rect 88628 327570 88656 329938
rect 89456 327570 89484 338263
rect 89640 330002 89668 358799
rect 90376 354822 90404 388991
rect 92032 383654 92060 390374
rect 93412 388482 93440 390918
rect 102598 390895 102654 390904
rect 110418 390960 110474 390969
rect 110418 390895 110474 390904
rect 111154 390960 111210 390969
rect 111210 390918 111504 390946
rect 111154 390895 111210 390904
rect 100666 390552 100722 390561
rect 100722 390524 100832 390538
rect 100722 390510 100846 390524
rect 100666 390487 100722 390496
rect 97354 390416 97410 390425
rect 94240 390374 94576 390402
rect 95896 390374 96232 390402
rect 93400 388476 93452 388482
rect 93400 388418 93452 388424
rect 93766 388376 93822 388385
rect 93766 388311 93822 388320
rect 93676 388068 93728 388074
rect 93676 388010 93728 388016
rect 92032 383626 92336 383654
rect 91006 371376 91062 371385
rect 91006 371311 91062 371320
rect 90364 354816 90416 354822
rect 90364 354758 90416 354764
rect 90376 350606 90404 354758
rect 90364 350600 90416 350606
rect 90364 350542 90416 350548
rect 89904 334008 89956 334014
rect 89904 333950 89956 333956
rect 89628 329996 89680 330002
rect 89628 329938 89680 329944
rect 86420 327542 86848 327570
rect 87156 327542 87584 327570
rect 88320 327542 88656 327570
rect 89056 327542 89484 327570
rect 89916 327298 89944 333950
rect 91020 332586 91048 371311
rect 92308 349110 92336 383626
rect 93688 365702 93716 388010
rect 93124 365696 93176 365702
rect 93124 365638 93176 365644
rect 93676 365696 93728 365702
rect 93676 365638 93728 365644
rect 92296 349104 92348 349110
rect 92296 349046 92348 349052
rect 93136 347070 93164 365638
rect 93780 350713 93808 388311
rect 94240 388074 94268 390374
rect 95896 389065 95924 390374
rect 98826 390416 98882 390425
rect 97410 390374 97856 390402
rect 97354 390351 97410 390360
rect 95882 389056 95938 389065
rect 95882 388991 95938 389000
rect 94228 388068 94280 388074
rect 94228 388010 94280 388016
rect 94502 369880 94558 369889
rect 94502 369815 94558 369824
rect 93214 350704 93270 350713
rect 93214 350639 93270 350648
rect 93766 350704 93822 350713
rect 93766 350639 93822 350648
rect 93124 347064 93176 347070
rect 93124 347006 93176 347012
rect 92388 345704 92440 345710
rect 92388 345646 92440 345652
rect 92400 335354 92428 345646
rect 93228 340202 93256 350639
rect 93216 340196 93268 340202
rect 93216 340138 93268 340144
rect 92848 336864 92900 336870
rect 92848 336806 92900 336812
rect 92216 335326 92428 335354
rect 91560 333124 91612 333130
rect 91560 333066 91612 333072
rect 91008 332580 91060 332586
rect 91008 332522 91060 332528
rect 90822 331392 90878 331401
rect 90822 331327 90878 331336
rect 90836 327570 90864 331327
rect 91572 327570 91600 333066
rect 92216 327570 92244 335326
rect 92754 334384 92810 334393
rect 92754 334319 92810 334328
rect 92768 327570 92796 334319
rect 90528 327542 90864 327570
rect 91264 327542 91600 327570
rect 91816 327542 92244 327570
rect 92552 327542 92796 327570
rect 92860 327570 92888 336806
rect 94516 333130 94544 369815
rect 97828 352578 97856 390374
rect 98882 390374 99328 390402
rect 98826 390351 98882 390360
rect 98642 368384 98698 368393
rect 98642 368319 98698 368328
rect 98656 367169 98684 368319
rect 99300 367810 99328 390374
rect 100818 390130 100846 390510
rect 100772 390102 100846 390130
rect 100114 389872 100170 389881
rect 100114 389807 100170 389816
rect 99288 367804 99340 367810
rect 99288 367746 99340 367752
rect 98642 367160 98698 367169
rect 98642 367095 98698 367104
rect 97816 352572 97868 352578
rect 97816 352514 97868 352520
rect 96528 348424 96580 348430
rect 96528 348366 96580 348372
rect 96436 347064 96488 347070
rect 96436 347006 96488 347012
rect 95146 341048 95202 341057
rect 95146 340983 95202 340992
rect 94504 333124 94556 333130
rect 94504 333066 94556 333072
rect 93860 332580 93912 332586
rect 93860 332522 93912 332528
rect 93872 327570 93900 332522
rect 95160 327570 95188 340983
rect 96448 331158 96476 347006
rect 95792 331152 95844 331158
rect 95792 331094 95844 331100
rect 96436 331152 96488 331158
rect 96436 331094 96488 331100
rect 95804 327570 95832 331094
rect 96540 327570 96568 348366
rect 97264 343664 97316 343670
rect 97264 343606 97316 343612
rect 97276 330546 97304 343606
rect 97906 339824 97962 339833
rect 97906 339759 97962 339768
rect 97264 330540 97316 330546
rect 97264 330482 97316 330488
rect 97264 330132 97316 330138
rect 97264 330074 97316 330080
rect 97276 327570 97304 330074
rect 97920 327570 97948 339759
rect 98656 333305 98684 367095
rect 98736 363044 98788 363050
rect 98736 362986 98788 362992
rect 98642 333296 98698 333305
rect 98642 333231 98698 333240
rect 98550 332752 98606 332761
rect 98550 332687 98606 332696
rect 98564 327570 98592 332687
rect 98748 330138 98776 362986
rect 100128 343738 100156 389807
rect 99380 343732 99432 343738
rect 99380 343674 99432 343680
rect 100116 343732 100168 343738
rect 100116 343674 100168 343680
rect 99286 330440 99342 330449
rect 99286 330375 99342 330384
rect 98736 330132 98788 330138
rect 98736 330074 98788 330080
rect 99300 327570 99328 330375
rect 92860 327542 93288 327570
rect 93872 327542 94024 327570
rect 94760 327542 95188 327570
rect 95496 327542 95832 327570
rect 96232 327542 96568 327570
rect 96968 327542 97304 327570
rect 97520 327542 97948 327570
rect 98256 327542 98592 327570
rect 98992 327542 99328 327570
rect 93872 327321 93900 327542
rect 89792 327270 89944 327298
rect 93858 327312 93914 327321
rect 93858 327247 93914 327256
rect 77298 327176 77354 327185
rect 83922 327176 83978 327185
rect 77354 327134 77648 327162
rect 77298 327111 77354 327120
rect 83978 327134 84088 327162
rect 83922 327111 83978 327120
rect 99392 327078 99420 343674
rect 100772 341465 100800 390102
rect 102612 389065 102640 390895
rect 105082 390416 105138 390425
rect 103776 390374 104112 390402
rect 104084 389162 104112 390374
rect 106554 390416 106610 390425
rect 105138 390374 105676 390402
rect 105082 390351 105138 390360
rect 104072 389156 104124 389162
rect 104072 389098 104124 389104
rect 102598 389056 102654 389065
rect 102598 388991 102654 389000
rect 105542 389056 105598 389065
rect 105542 388991 105598 389000
rect 104900 376780 104952 376786
rect 104900 376722 104952 376728
rect 102046 360224 102102 360233
rect 102046 360159 102102 360168
rect 101402 346488 101458 346497
rect 101402 346423 101458 346432
rect 100758 341456 100814 341465
rect 100758 341391 100814 341400
rect 101416 330138 101444 346423
rect 101496 330540 101548 330546
rect 101496 330482 101548 330488
rect 100024 330132 100076 330138
rect 100024 330074 100076 330080
rect 101404 330132 101456 330138
rect 101404 330074 101456 330080
rect 100036 327570 100064 330074
rect 101508 327570 101536 330482
rect 102060 327570 102088 360159
rect 102140 356176 102192 356182
rect 102140 356118 102192 356124
rect 99728 327542 100064 327570
rect 101200 327542 101536 327570
rect 101936 327542 102088 327570
rect 102152 327570 102180 356118
rect 104808 351280 104860 351286
rect 104808 351222 104860 351228
rect 102782 342272 102838 342281
rect 102782 342207 102838 342216
rect 102796 327570 102824 342207
rect 104256 334008 104308 334014
rect 104256 333950 104308 333956
rect 104268 327570 104296 333950
rect 104820 327570 104848 351222
rect 104912 345014 104940 376722
rect 105556 347041 105584 388991
rect 105648 387025 105676 390374
rect 108026 390416 108082 390425
rect 106610 390374 107332 390402
rect 106554 390351 106610 390360
rect 105634 387016 105690 387025
rect 105634 386951 105690 386960
rect 105648 358086 105676 386951
rect 107304 383654 107332 390374
rect 109498 390416 109554 390425
rect 108082 390374 108804 390402
rect 108026 390351 108082 390360
rect 108302 389328 108358 389337
rect 108302 389263 108358 389272
rect 108316 388385 108344 389263
rect 108302 388376 108358 388385
rect 108302 388311 108358 388320
rect 108302 385656 108358 385665
rect 108302 385591 108358 385600
rect 107304 383626 107516 383654
rect 107488 369238 107516 383626
rect 107476 369232 107528 369238
rect 107476 369174 107528 369180
rect 108316 364334 108344 385591
rect 108776 382974 108804 390374
rect 109554 390374 110276 390402
rect 109498 390351 109554 390360
rect 110248 383654 110276 390374
rect 110248 383626 110368 383654
rect 108764 382968 108816 382974
rect 108764 382910 108816 382916
rect 107856 364306 108344 364334
rect 107856 363089 107884 364306
rect 107842 363080 107898 363089
rect 107842 363015 107898 363024
rect 105636 358080 105688 358086
rect 105636 358022 105688 358028
rect 106922 352064 106978 352073
rect 106922 351999 106978 352008
rect 105542 347032 105598 347041
rect 105542 346967 105598 346976
rect 104912 344986 105032 345014
rect 102152 327542 102672 327570
rect 102796 327542 103224 327570
rect 103960 327542 104296 327570
rect 104696 327542 104848 327570
rect 105004 327570 105032 344986
rect 106186 342544 106242 342553
rect 106186 342479 106242 342488
rect 106200 327842 106228 342479
rect 106936 330449 106964 351999
rect 107750 335472 107806 335481
rect 107750 335407 107806 335416
rect 107200 331288 107252 331294
rect 107200 331230 107252 331236
rect 106922 330440 106978 330449
rect 106922 330375 106978 330384
rect 106154 327814 106228 327842
rect 105004 327542 105432 327570
rect 106154 327556 106182 327814
rect 107212 327570 107240 331230
rect 107764 330410 107792 335407
rect 107752 330404 107804 330410
rect 107752 330346 107804 330352
rect 107856 327570 107884 363015
rect 110340 351218 110368 383626
rect 110432 380254 110460 390895
rect 115848 390584 115900 390590
rect 115848 390526 115900 390532
rect 112640 390374 112976 390402
rect 114112 390374 114448 390402
rect 112640 389065 112668 390374
rect 114112 389337 114140 390374
rect 114098 389328 114154 389337
rect 114098 389263 114154 389272
rect 111798 389056 111854 389065
rect 111798 388991 111854 389000
rect 112626 389056 112682 389065
rect 112626 388991 112682 389000
rect 111708 387116 111760 387122
rect 111708 387058 111760 387064
rect 110420 380248 110472 380254
rect 110420 380190 110472 380196
rect 110328 351212 110380 351218
rect 110328 351154 110380 351160
rect 111720 347857 111748 387058
rect 111812 369170 111840 388991
rect 112444 388476 112496 388482
rect 112444 388418 112496 388424
rect 111800 369164 111852 369170
rect 111800 369106 111852 369112
rect 112456 356697 112484 388418
rect 115860 360262 115888 390526
rect 115938 390416 115994 390425
rect 120262 390416 120318 390425
rect 115994 390374 116104 390402
rect 117576 390374 117820 390402
rect 115938 390351 115994 390360
rect 115204 360256 115256 360262
rect 115204 360198 115256 360204
rect 115848 360256 115900 360262
rect 115848 360198 115900 360204
rect 112442 356688 112498 356697
rect 112442 356623 112498 356632
rect 112442 353696 112498 353705
rect 112442 353631 112498 353640
rect 110418 347848 110474 347857
rect 110418 347783 110474 347792
rect 111706 347848 111762 347857
rect 111706 347783 111762 347792
rect 110432 345014 110460 347783
rect 110432 344986 110736 345014
rect 108762 334112 108818 334121
rect 108762 334047 108818 334056
rect 108028 330404 108080 330410
rect 108028 330346 108080 330352
rect 106904 327542 107240 327570
rect 107640 327542 107884 327570
rect 108040 327570 108068 330346
rect 108040 327542 108376 327570
rect 108776 327298 108804 334047
rect 109958 331120 110014 331129
rect 109958 331055 110014 331064
rect 109972 327570 110000 331055
rect 110604 330132 110656 330138
rect 110604 330074 110656 330080
rect 110616 327570 110644 330074
rect 109664 327542 110000 327570
rect 110400 327542 110644 327570
rect 110708 327570 110736 344986
rect 111706 343768 111762 343777
rect 111706 343703 111762 343712
rect 111720 330138 111748 343703
rect 111798 339688 111854 339697
rect 111798 339623 111854 339632
rect 111708 330132 111760 330138
rect 111708 330074 111760 330080
rect 111812 327842 111840 339623
rect 112456 336025 112484 353631
rect 113086 349208 113142 349217
rect 113086 349143 113142 349152
rect 112442 336016 112498 336025
rect 112442 335951 112498 335960
rect 113100 335354 113128 349143
rect 114466 343904 114522 343913
rect 114466 343839 114522 343848
rect 113180 336048 113232 336054
rect 113180 335990 113232 335996
rect 113008 335326 113128 335354
rect 111812 327814 111886 327842
rect 110708 327542 111136 327570
rect 111858 327556 111886 327814
rect 113008 327570 113036 335326
rect 113192 334626 113220 335990
rect 113180 334620 113232 334626
rect 113180 334562 113232 334568
rect 113640 332716 113692 332722
rect 113640 332658 113692 332664
rect 113652 327570 113680 332658
rect 114480 327570 114508 343839
rect 115216 335354 115244 360198
rect 115952 349761 115980 390351
rect 117792 389230 117820 390374
rect 118712 390374 119048 390402
rect 120184 390374 120262 390402
rect 118712 389473 118740 390374
rect 118698 389464 118754 389473
rect 118698 389399 118754 389408
rect 117780 389224 117832 389230
rect 117778 389192 117780 389201
rect 117832 389192 117834 389201
rect 117778 389127 117834 389136
rect 118712 374746 118740 389399
rect 120184 389094 120212 390374
rect 120318 390374 120520 390402
rect 120262 390351 120318 390360
rect 120276 390291 120304 390351
rect 119436 389088 119488 389094
rect 119436 389030 119488 389036
rect 120172 389088 120224 389094
rect 120172 389030 120224 389036
rect 119342 386336 119398 386345
rect 119342 386271 119398 386280
rect 118700 374740 118752 374746
rect 118700 374682 118752 374688
rect 118712 373994 118740 374682
rect 118620 373966 118740 373994
rect 118620 373318 118648 373966
rect 118608 373312 118660 373318
rect 118608 373254 118660 373260
rect 117318 365664 117374 365673
rect 117318 365599 117374 365608
rect 117332 364449 117360 365599
rect 117318 364440 117374 364449
rect 117318 364375 117374 364384
rect 117228 361616 117280 361622
rect 117228 361558 117280 361564
rect 116582 355328 116638 355337
rect 116582 355263 116638 355272
rect 115938 349752 115994 349761
rect 115938 349687 115994 349696
rect 116596 347070 116624 355263
rect 116584 347064 116636 347070
rect 116584 347006 116636 347012
rect 115294 346624 115350 346633
rect 115294 346559 115350 346568
rect 115032 335326 115244 335354
rect 115032 328545 115060 335326
rect 115308 331129 115336 346559
rect 115940 339516 115992 339522
rect 115940 339458 115992 339464
rect 115664 334076 115716 334082
rect 115664 334018 115716 334024
rect 115294 331120 115350 331129
rect 115294 331055 115350 331064
rect 115018 328536 115074 328545
rect 115018 328471 115074 328480
rect 115032 327570 115060 328471
rect 115676 327570 115704 334018
rect 112608 327542 113036 327570
rect 113344 327542 113680 327570
rect 114080 327542 114508 327570
rect 114632 327542 115060 327570
rect 115368 327542 115704 327570
rect 115952 327570 115980 339458
rect 117240 327570 117268 361558
rect 117332 345014 117360 364375
rect 119356 349178 119384 386271
rect 119448 374649 119476 389030
rect 120644 387122 120672 416735
rect 120736 411097 120764 562294
rect 121460 556232 121512 556238
rect 121460 556174 121512 556180
rect 120814 419520 120870 419529
rect 120814 419455 120870 419464
rect 120722 411088 120778 411097
rect 120722 411023 120778 411032
rect 120828 390590 120856 419455
rect 121182 410544 121238 410553
rect 121182 410479 121238 410488
rect 121196 409902 121224 410479
rect 121184 409896 121236 409902
rect 121184 409838 121236 409844
rect 121472 392601 121500 556174
rect 121552 548548 121604 548554
rect 121552 548490 121604 548496
rect 121564 396953 121592 548490
rect 121656 428505 121684 578206
rect 123208 558204 123260 558210
rect 123208 558146 123260 558152
rect 123114 450528 123170 450537
rect 123114 450463 123170 450472
rect 122932 447840 122984 447846
rect 122932 447782 122984 447788
rect 123022 447808 123078 447817
rect 122746 430944 122802 430953
rect 122746 430879 122802 430888
rect 121642 428496 121698 428505
rect 121642 428431 121698 428440
rect 121550 396944 121606 396953
rect 121550 396879 121606 396888
rect 121564 396098 121592 396879
rect 121552 396092 121604 396098
rect 121552 396034 121604 396040
rect 121458 392592 121514 392601
rect 121458 392527 121514 392536
rect 120816 390584 120868 390590
rect 120816 390526 120868 390532
rect 120632 387116 120684 387122
rect 120632 387058 120684 387064
rect 119434 374640 119490 374649
rect 119434 374575 119490 374584
rect 121366 364576 121422 364585
rect 121366 364511 121422 364520
rect 120722 360360 120778 360369
rect 120722 360295 120778 360304
rect 119434 357504 119490 357513
rect 119434 357439 119490 357448
rect 118700 349172 118752 349178
rect 118700 349114 118752 349120
rect 119344 349172 119396 349178
rect 119344 349114 119396 349120
rect 117332 344986 117912 345014
rect 117780 331152 117832 331158
rect 117780 331094 117832 331100
rect 117792 327570 117820 331094
rect 115952 327542 116104 327570
rect 116840 327542 117268 327570
rect 117576 327542 117820 327570
rect 117884 327570 117912 344986
rect 118606 340912 118662 340921
rect 118606 340847 118662 340856
rect 118620 331158 118648 340847
rect 118712 331158 118740 349114
rect 119448 349110 119476 357439
rect 120736 351286 120764 360295
rect 120724 351280 120776 351286
rect 120724 351222 120776 351228
rect 118792 349104 118844 349110
rect 118792 349046 118844 349052
rect 119436 349104 119488 349110
rect 119436 349046 119488 349052
rect 118608 331152 118660 331158
rect 118608 331094 118660 331100
rect 118700 331152 118752 331158
rect 118700 331094 118752 331100
rect 118804 327570 118832 349046
rect 120080 337408 120132 337414
rect 120080 337350 120132 337356
rect 119436 331152 119488 331158
rect 119436 331094 119488 331100
rect 119448 327570 119476 331094
rect 120092 327570 120120 337350
rect 121380 327570 121408 364511
rect 122760 353433 122788 430879
rect 122944 424153 122972 447782
rect 123022 447743 123078 447752
rect 122930 424144 122986 424153
rect 122930 424079 122986 424088
rect 122944 412634 122972 424079
rect 123036 417353 123064 447743
rect 123128 433129 123156 450463
rect 123114 433120 123170 433129
rect 123114 433055 123170 433064
rect 123114 428496 123170 428505
rect 123114 428431 123170 428440
rect 123022 417344 123078 417353
rect 123022 417279 123078 417288
rect 123022 412720 123078 412729
rect 123022 412655 123078 412664
rect 122852 412606 122972 412634
rect 123036 412622 123064 412655
rect 123024 412616 123076 412622
rect 122852 378729 122880 412606
rect 123024 412558 123076 412564
rect 123036 411330 123064 412558
rect 123024 411324 123076 411330
rect 123024 411266 123076 411272
rect 122930 394768 122986 394777
rect 122930 394703 122986 394712
rect 122944 384334 122972 394703
rect 122932 384328 122984 384334
rect 122932 384270 122984 384276
rect 122838 378720 122894 378729
rect 122838 378655 122894 378664
rect 122932 365016 122984 365022
rect 122932 364958 122984 364964
rect 122944 358902 122972 364958
rect 123128 359514 123156 428431
rect 123220 421977 123248 558146
rect 123496 447681 123524 582927
rect 123482 447672 123538 447681
rect 123482 447607 123538 447616
rect 124126 439920 124182 439929
rect 124126 439855 124182 439864
rect 124140 439550 124168 439855
rect 124128 439544 124180 439550
rect 124128 439486 124180 439492
rect 124232 438190 124260 584394
rect 124876 536761 124904 702986
rect 126244 702908 126296 702914
rect 126244 702850 126296 702856
rect 125600 557592 125652 557598
rect 125600 557534 125652 557540
rect 124862 536752 124918 536761
rect 124862 536687 124918 536696
rect 124956 452668 125008 452674
rect 124956 452610 125008 452616
rect 124864 445800 124916 445806
rect 124864 445742 124916 445748
rect 123668 438184 123720 438190
rect 123668 438126 123720 438132
rect 124220 438184 124272 438190
rect 124220 438126 124272 438132
rect 123680 437753 123708 438126
rect 123666 437744 123722 437753
rect 123666 437679 123722 437688
rect 123850 433120 123906 433129
rect 123850 433055 123906 433064
rect 123864 432614 123892 433055
rect 123852 432608 123904 432614
rect 123852 432550 123904 432556
rect 123206 421968 123262 421977
rect 123206 421903 123262 421912
rect 123220 421598 123248 421903
rect 123208 421592 123260 421598
rect 123208 421534 123260 421540
rect 124128 415200 124180 415206
rect 124126 415168 124128 415177
rect 124180 415168 124182 415177
rect 124126 415103 124182 415112
rect 123484 411324 123536 411330
rect 123484 411266 123536 411272
rect 123496 381546 123524 411266
rect 124126 408368 124182 408377
rect 124126 408303 124182 408312
rect 124140 407794 124168 408303
rect 124128 407788 124180 407794
rect 124128 407730 124180 407736
rect 124126 406192 124182 406201
rect 124126 406127 124128 406136
rect 124180 406127 124182 406136
rect 124128 406098 124180 406104
rect 124034 403744 124090 403753
rect 124034 403679 124090 403688
rect 124048 403034 124076 403679
rect 124036 403028 124088 403034
rect 124036 402970 124088 402976
rect 124128 401600 124180 401606
rect 124126 401568 124128 401577
rect 124180 401568 124182 401577
rect 124126 401503 124182 401512
rect 123668 400172 123720 400178
rect 123668 400114 123720 400120
rect 123680 399401 123708 400114
rect 123666 399392 123722 399401
rect 123666 399327 123722 399336
rect 123668 396024 123720 396030
rect 123668 395966 123720 395972
rect 123680 394777 123708 395966
rect 123666 394768 123722 394777
rect 123666 394703 123722 394712
rect 123484 381540 123536 381546
rect 123484 381482 123536 381488
rect 123116 359508 123168 359514
rect 123116 359450 123168 359456
rect 122932 358896 122984 358902
rect 122932 358838 122984 358844
rect 121458 353424 121514 353433
rect 121458 353359 121514 353368
rect 122746 353424 122802 353433
rect 122746 353359 122802 353368
rect 121472 345710 121500 353359
rect 122748 348492 122800 348498
rect 122748 348434 122800 348440
rect 121460 345704 121512 345710
rect 121460 345646 121512 345652
rect 122102 328536 122158 328545
rect 122102 328471 122158 328480
rect 122116 327570 122144 328471
rect 122760 327570 122788 348434
rect 117884 327542 118312 327570
rect 118804 327542 119048 327570
rect 119448 327542 119784 327570
rect 120092 327542 120336 327570
rect 121072 327542 121408 327570
rect 121808 327542 122144 327570
rect 122544 327542 122788 327570
rect 108776 327270 108928 327298
rect 122944 327146 122972 358838
rect 123484 350600 123536 350606
rect 123484 350542 123536 350548
rect 123496 331226 123524 350542
rect 124876 345681 124904 445742
rect 124968 400246 124996 452610
rect 124956 400240 125008 400246
rect 124956 400182 125008 400188
rect 125612 396030 125640 557534
rect 126256 546446 126284 702850
rect 129004 702704 129056 702710
rect 129004 702646 129056 702652
rect 128544 593428 128596 593434
rect 128544 593370 128596 593376
rect 126980 565888 127032 565894
rect 126980 565830 127032 565836
rect 126244 546440 126296 546446
rect 126244 546382 126296 546388
rect 125692 465792 125744 465798
rect 125692 465734 125744 465740
rect 125704 439550 125732 465734
rect 126244 444508 126296 444514
rect 126244 444450 126296 444456
rect 125692 439544 125744 439550
rect 125692 439486 125744 439492
rect 125600 396024 125652 396030
rect 125600 395966 125652 395972
rect 124956 380180 125008 380186
rect 124956 380122 125008 380128
rect 124968 358834 124996 380122
rect 126256 368966 126284 444450
rect 126992 406994 127020 565830
rect 128452 454164 128504 454170
rect 128452 454106 128504 454112
rect 128360 449200 128412 449206
rect 128360 449142 128412 449148
rect 128266 446312 128322 446321
rect 128266 446247 128322 446256
rect 128280 445913 128308 446247
rect 128266 445904 128322 445913
rect 128266 445839 128322 445848
rect 126900 406966 127020 406994
rect 126900 406162 126928 406966
rect 126888 406156 126940 406162
rect 126888 406098 126940 406104
rect 125600 368960 125652 368966
rect 125600 368902 125652 368908
rect 126244 368960 126296 368966
rect 126244 368902 126296 368908
rect 124956 358828 125008 358834
rect 124956 358770 125008 358776
rect 124862 345672 124918 345681
rect 124862 345607 124918 345616
rect 123484 331220 123536 331226
rect 123484 331162 123536 331168
rect 123496 327570 123524 331162
rect 124968 328506 124996 358770
rect 125506 338192 125562 338201
rect 125506 338127 125562 338136
rect 124956 328500 125008 328506
rect 124956 328442 125008 328448
rect 124968 327570 124996 328442
rect 125520 327842 125548 338127
rect 123280 327542 123524 327570
rect 124752 327542 124996 327570
rect 125474 327814 125548 327842
rect 125474 327556 125502 327814
rect 125612 327570 125640 368902
rect 126256 368558 126284 368902
rect 126244 368552 126296 368558
rect 126244 368494 126296 368500
rect 126900 357377 126928 406098
rect 128280 363633 128308 445839
rect 128372 412622 128400 449142
rect 128360 412616 128412 412622
rect 128360 412558 128412 412564
rect 128360 365696 128412 365702
rect 128360 365638 128412 365644
rect 128372 365022 128400 365638
rect 128360 365016 128412 365022
rect 128360 364958 128412 364964
rect 128266 363624 128322 363633
rect 128266 363559 128322 363568
rect 126978 362264 127034 362273
rect 126978 362199 127034 362208
rect 125690 357368 125746 357377
rect 125690 357303 125746 357312
rect 126886 357368 126942 357377
rect 126886 357303 126942 357312
rect 125704 356153 125732 357303
rect 125690 356144 125746 356153
rect 125690 356079 125746 356088
rect 125704 345014 125732 356079
rect 126992 345014 127020 362199
rect 128360 354748 128412 354754
rect 128360 354690 128412 354696
rect 128372 345014 128400 354690
rect 128464 348430 128492 454106
rect 128556 446321 128584 593370
rect 129016 544406 129044 702646
rect 129740 571396 129792 571402
rect 129740 571338 129792 571344
rect 129004 544400 129056 544406
rect 129004 544342 129056 544348
rect 129002 536072 129058 536081
rect 129002 536007 129058 536016
rect 128542 446312 128598 446321
rect 128542 446247 128598 446256
rect 129016 365702 129044 536007
rect 129752 415206 129780 571338
rect 130396 536790 130424 703190
rect 133144 700324 133196 700330
rect 133144 700266 133196 700272
rect 133156 538218 133184 700266
rect 133880 567248 133932 567254
rect 133880 567190 133932 567196
rect 133236 563100 133288 563106
rect 133236 563042 133288 563048
rect 133144 538212 133196 538218
rect 133144 538154 133196 538160
rect 130384 536784 130436 536790
rect 130384 536726 130436 536732
rect 130384 448588 130436 448594
rect 130384 448530 130436 448536
rect 129740 415200 129792 415206
rect 129740 415142 129792 415148
rect 129752 414730 129780 415142
rect 129740 414724 129792 414730
rect 129740 414666 129792 414672
rect 129740 371340 129792 371346
rect 129740 371282 129792 371288
rect 129004 365696 129056 365702
rect 129004 365638 129056 365644
rect 128452 348424 128504 348430
rect 128450 348392 128452 348401
rect 128504 348392 128506 348401
rect 128450 348327 128506 348336
rect 125704 344986 126376 345014
rect 126992 344986 127848 345014
rect 128372 344986 128584 345014
rect 126348 327570 126376 344986
rect 127716 330404 127768 330410
rect 127716 330346 127768 330352
rect 127728 327570 127756 330346
rect 125612 327542 126040 327570
rect 126348 327542 126776 327570
rect 127512 327542 127756 327570
rect 127820 327570 127848 344986
rect 128556 327570 128584 344986
rect 129752 331498 129780 371282
rect 129830 352608 129886 352617
rect 129830 352543 129886 352552
rect 129844 351937 129872 352543
rect 129830 351928 129886 351937
rect 129830 351863 129886 351872
rect 129844 345014 129872 351863
rect 130396 349897 130424 448530
rect 130474 447264 130530 447273
rect 130474 447199 130530 447208
rect 130488 365809 130516 447199
rect 131120 414724 131172 414730
rect 131120 414666 131172 414672
rect 130474 365800 130530 365809
rect 130474 365735 130530 365744
rect 130382 349888 130438 349897
rect 130382 349823 130438 349832
rect 130488 348498 130516 365735
rect 131132 355337 131160 414666
rect 133248 401606 133276 563042
rect 133892 407794 133920 567190
rect 136652 541686 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202604 703656 202656 703662
rect 202604 703598 202656 703604
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702545 154160 703520
rect 154118 702536 154174 702545
rect 154118 702471 154174 702480
rect 170324 702434 170352 703520
rect 202616 703474 202644 703598
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234988 703588 235040 703594
rect 234988 703530 235040 703536
rect 202800 703474 202828 703520
rect 202616 703446 202828 703474
rect 169772 702406 170352 702434
rect 169772 596834 169800 702406
rect 218992 700330 219020 703520
rect 235000 703474 235028 703530
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267464 703520 267516 703526
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 703474 267688 703520
rect 267516 703468 267688 703474
rect 267464 703462 267688 703468
rect 267476 703446 267688 703462
rect 283852 703390 283880 703520
rect 300136 703458 300164 703520
rect 300124 703452 300176 703458
rect 300124 703394 300176 703400
rect 283840 703384 283892 703390
rect 283840 703326 283892 703332
rect 332520 703322 332548 703520
rect 332508 703316 332560 703322
rect 332508 703258 332560 703264
rect 348804 703186 348832 703520
rect 348792 703180 348844 703186
rect 348792 703122 348844 703128
rect 364996 702982 365024 703520
rect 397472 703118 397500 703520
rect 413664 703254 413692 703520
rect 413652 703248 413704 703254
rect 413652 703190 413704 703196
rect 397460 703112 397512 703118
rect 397460 703054 397512 703060
rect 429856 703050 429884 703520
rect 429844 703044 429896 703050
rect 429844 702986 429896 702992
rect 364984 702976 365036 702982
rect 364984 702918 365036 702924
rect 462332 702914 462360 703520
rect 462320 702908 462372 702914
rect 462320 702850 462372 702856
rect 478524 702778 478552 703520
rect 494808 702846 494836 703520
rect 494796 702840 494848 702846
rect 494796 702782 494848 702788
rect 478512 702772 478564 702778
rect 478512 702714 478564 702720
rect 527192 702642 527220 703520
rect 543476 702710 543504 703520
rect 543464 702704 543516 702710
rect 543464 702646 543516 702652
rect 527180 702636 527232 702642
rect 527180 702578 527232 702584
rect 559668 702506 559696 703520
rect 580264 702568 580316 702574
rect 580264 702510 580316 702516
rect 559656 702500 559708 702506
rect 559656 702442 559708 702448
rect 218980 700324 219032 700330
rect 218980 700266 219032 700272
rect 580276 670721 580304 702510
rect 582378 697232 582434 697241
rect 582378 697167 582434 697176
rect 580262 670712 580318 670721
rect 580262 670647 580318 670656
rect 169760 596828 169812 596834
rect 169760 596770 169812 596776
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 589937 580212 590951
rect 580170 589928 580226 589937
rect 580170 589863 580226 589872
rect 580262 577688 580318 577697
rect 580262 577623 580318 577632
rect 143448 577516 143500 577522
rect 143448 577458 143500 577464
rect 143460 576910 143488 577458
rect 142160 576904 142212 576910
rect 142160 576846 142212 576852
rect 143448 576904 143500 576910
rect 143448 576846 143500 576852
rect 136640 541680 136692 541686
rect 136640 541622 136692 541628
rect 134524 421592 134576 421598
rect 134524 421534 134576 421540
rect 133880 407788 133932 407794
rect 133880 407730 133932 407736
rect 133786 401704 133842 401713
rect 133786 401639 133842 401648
rect 133800 401606 133828 401639
rect 133236 401600 133288 401606
rect 133236 401542 133288 401548
rect 133788 401600 133840 401606
rect 133788 401542 133840 401548
rect 132500 367124 132552 367130
rect 132500 367066 132552 367072
rect 131118 355328 131174 355337
rect 131118 355263 131174 355272
rect 130476 348492 130528 348498
rect 130476 348434 130528 348440
rect 129844 344986 129964 345014
rect 129740 331492 129792 331498
rect 129740 331434 129792 331440
rect 129740 331356 129792 331362
rect 129740 331298 129792 331304
rect 129752 329225 129780 331298
rect 129738 329216 129794 329225
rect 129738 329151 129794 329160
rect 129936 327570 129964 344986
rect 132038 331528 132094 331537
rect 130108 331492 130160 331498
rect 132038 331463 132094 331472
rect 130108 331434 130160 331440
rect 127820 327542 128248 327570
rect 128556 327542 128984 327570
rect 129720 327542 129964 327570
rect 130120 327570 130148 331434
rect 131486 329896 131542 329905
rect 131486 329831 131542 329840
rect 130120 327542 130456 327570
rect 131500 327434 131528 329831
rect 132052 327570 132080 331463
rect 132512 330290 132540 367066
rect 134536 349761 134564 421534
rect 135904 409896 135956 409902
rect 135904 409838 135956 409844
rect 134616 407788 134668 407794
rect 134616 407730 134668 407736
rect 134628 353394 134656 407730
rect 135916 355609 135944 409838
rect 136652 389162 136680 541622
rect 137282 444544 137338 444553
rect 137282 444479 137338 444488
rect 136640 389156 136692 389162
rect 136640 389098 136692 389104
rect 136652 388793 136680 389098
rect 136638 388784 136694 388793
rect 136638 388719 136694 388728
rect 137296 367062 137324 444479
rect 142172 425649 142200 576846
rect 579802 537840 579858 537849
rect 579802 537775 579858 537784
rect 579816 537538 579844 537775
rect 579804 537532 579856 537538
rect 579804 537474 579856 537480
rect 580276 534070 580304 577623
rect 582392 536081 582420 697167
rect 582470 683904 582526 683913
rect 582470 683839 582526 683848
rect 582484 577522 582512 683839
rect 582562 644056 582618 644065
rect 582562 643991 582618 644000
rect 582472 577516 582524 577522
rect 582472 577458 582524 577464
rect 582472 554804 582524 554810
rect 582472 554746 582524 554752
rect 582378 536072 582434 536081
rect 582378 536007 582434 536016
rect 580264 534064 580316 534070
rect 580264 534006 580316 534012
rect 582484 524521 582512 554746
rect 582576 538286 582604 643991
rect 582654 630864 582710 630873
rect 582654 630799 582710 630808
rect 582668 540938 582696 630799
rect 582746 617536 582802 617545
rect 582746 617471 582802 617480
rect 582760 595474 582788 617471
rect 582748 595468 582800 595474
rect 582748 595410 582800 595416
rect 582748 593428 582800 593434
rect 582748 593370 582800 593376
rect 582760 564369 582788 593370
rect 582746 564360 582802 564369
rect 582746 564295 582802 564304
rect 582656 540932 582708 540938
rect 582656 540874 582708 540880
rect 582564 538280 582616 538286
rect 582564 538222 582616 538228
rect 582470 524512 582526 524521
rect 582470 524447 582526 524456
rect 580170 511320 580226 511329
rect 580170 511255 580172 511264
rect 580224 511255 580226 511264
rect 580172 511226 580224 511232
rect 582378 484664 582434 484673
rect 582378 484599 582434 484608
rect 178040 460964 178092 460970
rect 178040 460906 178092 460912
rect 152464 458856 152516 458862
rect 152464 458798 152516 458804
rect 144184 454096 144236 454102
rect 144184 454038 144236 454044
rect 142804 445868 142856 445874
rect 142804 445810 142856 445816
rect 142158 425640 142214 425649
rect 142158 425575 142214 425584
rect 142068 372632 142120 372638
rect 142068 372574 142120 372580
rect 137926 368520 137982 368529
rect 137926 368455 137982 368464
rect 137284 367056 137336 367062
rect 137284 366998 137336 367004
rect 137836 367056 137888 367062
rect 137836 366998 137888 367004
rect 137848 365838 137876 366998
rect 137836 365832 137888 365838
rect 137836 365774 137888 365780
rect 135902 355600 135958 355609
rect 135902 355535 135958 355544
rect 134616 353388 134668 353394
rect 134616 353330 134668 353336
rect 136546 350568 136602 350577
rect 136546 350503 136602 350512
rect 134522 349752 134578 349761
rect 134522 349687 134578 349696
rect 133144 347812 133196 347818
rect 133144 347754 133196 347760
rect 133156 337385 133184 347754
rect 135168 346520 135220 346526
rect 135168 346462 135220 346468
rect 134248 342372 134300 342378
rect 134248 342314 134300 342320
rect 133142 337376 133198 337385
rect 133142 337311 133198 337320
rect 132590 336968 132646 336977
rect 132590 336903 132646 336912
rect 132604 330546 132632 336903
rect 133328 332648 133380 332654
rect 133328 332590 133380 332596
rect 133420 332648 133472 332654
rect 133420 332590 133472 332596
rect 132592 330540 132644 330546
rect 132592 330482 132644 330488
rect 132512 330262 132816 330290
rect 132682 330168 132738 330177
rect 132682 330103 132738 330112
rect 132696 327570 132724 330103
rect 131744 327542 132080 327570
rect 132480 327542 132724 327570
rect 132788 327570 132816 330262
rect 133340 330154 133368 332590
rect 133432 330410 133460 332590
rect 133420 330404 133472 330410
rect 133420 330346 133472 330352
rect 134154 330304 134210 330313
rect 134154 330239 134210 330248
rect 133340 330126 133460 330154
rect 133326 330032 133382 330041
rect 133326 329967 133382 329976
rect 132788 327542 133216 327570
rect 131192 327406 131528 327434
rect 123680 327146 124016 327162
rect 122932 327140 122984 327146
rect 122932 327082 122984 327088
rect 123668 327140 124016 327146
rect 123720 327134 124016 327140
rect 123668 327082 123720 327088
rect 133340 327078 133368 329967
rect 133432 329118 133460 330126
rect 133420 329112 133472 329118
rect 133420 329054 133472 329060
rect 134168 327570 134196 330239
rect 133952 327542 134196 327570
rect 134260 327570 134288 342314
rect 135180 329798 135208 346462
rect 135168 329792 135220 329798
rect 135168 329734 135220 329740
rect 135180 328522 135208 329734
rect 135180 328494 135300 328522
rect 135272 327570 135300 328494
rect 136560 327570 136588 350503
rect 137008 338224 137060 338230
rect 137008 338166 137060 338172
rect 136916 329860 136968 329866
rect 136916 329802 136968 329808
rect 136928 327706 136956 329802
rect 134260 327542 134688 327570
rect 135272 327542 135424 327570
rect 136160 327542 136588 327570
rect 136882 327678 136956 327706
rect 136882 327556 136910 327678
rect 137020 327570 137048 338166
rect 137848 331158 137876 365774
rect 137836 331152 137888 331158
rect 137836 331094 137888 331100
rect 137940 329866 137968 368455
rect 140688 357468 140740 357474
rect 140688 357410 140740 357416
rect 138020 353388 138072 353394
rect 138020 353330 138072 353336
rect 137928 329860 137980 329866
rect 137928 329802 137980 329808
rect 138032 327570 138060 353330
rect 139398 337104 139454 337113
rect 139398 337039 139454 337048
rect 139412 336054 139440 337039
rect 139400 336048 139452 336054
rect 139400 335990 139452 335996
rect 139400 331152 139452 331158
rect 139400 331094 139452 331100
rect 139216 330404 139268 330410
rect 139216 330346 139268 330352
rect 139228 327570 139256 330346
rect 137020 327542 137448 327570
rect 138032 327542 138184 327570
rect 138920 327542 139256 327570
rect 139412 327570 139440 331094
rect 140700 327570 140728 357410
rect 141424 341080 141476 341086
rect 141424 341022 141476 341028
rect 140780 341012 140832 341018
rect 140780 340954 140832 340960
rect 140792 337414 140820 340954
rect 140780 337408 140832 337414
rect 140780 337350 140832 337356
rect 140780 336048 140832 336054
rect 140780 335990 140832 335996
rect 139412 327542 139656 327570
rect 140392 327542 140728 327570
rect 140792 327570 140820 335990
rect 141240 331356 141292 331362
rect 141240 331298 141292 331304
rect 140792 327542 141128 327570
rect 141252 327078 141280 331298
rect 141436 327078 141464 341022
rect 142080 327570 142108 372574
rect 142816 348430 142844 445810
rect 144196 351966 144224 454038
rect 145562 377360 145618 377369
rect 145562 377295 145618 377304
rect 145576 353841 145604 377295
rect 151084 369232 151136 369238
rect 151084 369174 151136 369180
rect 144918 353832 144974 353841
rect 144918 353767 144974 353776
rect 145562 353832 145618 353841
rect 145562 353767 145618 353776
rect 144826 353696 144882 353705
rect 144826 353631 144882 353640
rect 144840 352617 144868 353631
rect 144826 352608 144882 352617
rect 144826 352543 144882 352552
rect 144184 351960 144236 351966
rect 144184 351902 144236 351908
rect 142804 348424 142856 348430
rect 142804 348366 142856 348372
rect 143540 345160 143592 345166
rect 143540 345102 143592 345108
rect 143552 345014 143580 345102
rect 143552 344986 144316 345014
rect 143446 332888 143502 332897
rect 143446 332823 143502 332832
rect 143460 330410 143488 332823
rect 144184 331152 144236 331158
rect 144184 331094 144236 331100
rect 143448 330404 143500 330410
rect 143448 330346 143500 330352
rect 143448 328500 143500 328506
rect 143448 328442 143500 328448
rect 143460 327570 143488 328442
rect 144196 327570 144224 331094
rect 141864 327542 142108 327570
rect 143152 327542 143488 327570
rect 143888 327542 144224 327570
rect 144288 327570 144316 344986
rect 144826 341184 144882 341193
rect 144826 341119 144882 341128
rect 144840 331158 144868 341119
rect 144828 331152 144880 331158
rect 144828 331094 144880 331100
rect 144932 327570 144960 353767
rect 146300 351960 146352 351966
rect 146300 351902 146352 351908
rect 146312 345014 146340 351902
rect 146312 344986 146432 345014
rect 145380 340944 145432 340950
rect 146208 340944 146260 340950
rect 145380 340886 145432 340892
rect 146206 340912 146208 340921
rect 146260 340912 146262 340921
rect 145392 336025 145420 340886
rect 146206 340847 146262 340856
rect 145378 336016 145434 336025
rect 145378 335951 145434 335960
rect 146206 328536 146262 328545
rect 146206 328471 146262 328480
rect 146220 327570 146248 328471
rect 144288 327542 144624 327570
rect 144932 327542 145360 327570
rect 146096 327542 146248 327570
rect 146404 327570 146432 344986
rect 150346 340912 150402 340921
rect 150346 340847 150402 340856
rect 146944 336796 146996 336802
rect 146944 336738 146996 336744
rect 146956 336054 146984 336738
rect 146944 336048 146996 336054
rect 146944 335990 146996 335996
rect 149152 335368 149204 335374
rect 149152 335310 149204 335316
rect 147586 330032 147642 330041
rect 147586 329967 147642 329976
rect 147404 328500 147456 328506
rect 147404 328442 147456 328448
rect 146404 327542 146832 327570
rect 142600 327134 142936 327162
rect 99380 327072 99432 327078
rect 99380 327014 99432 327020
rect 100116 327072 100168 327078
rect 133328 327072 133380 327078
rect 100168 327020 100464 327026
rect 100116 327014 100464 327020
rect 133328 327014 133380 327020
rect 141240 327072 141292 327078
rect 141240 327014 141292 327020
rect 141424 327072 141476 327078
rect 142908 327049 142936 327134
rect 141424 327014 141476 327020
rect 142894 327040 142950 327049
rect 70030 326975 70032 326984
rect 70084 326975 70086 326984
rect 76564 327004 76616 327010
rect 70032 326946 70084 326952
rect 100128 326998 100464 327014
rect 147416 327010 147444 328442
rect 147600 327706 147628 329967
rect 149060 329860 149112 329866
rect 149060 329802 149112 329808
rect 149072 329089 149100 329802
rect 149058 329080 149114 329089
rect 149058 329015 149114 329024
rect 148968 328500 149020 328506
rect 148968 328442 149020 328448
rect 147554 327678 147628 327706
rect 148276 327720 148332 327729
rect 147554 327556 147582 327678
rect 148276 327655 148332 327664
rect 148290 327556 148318 327655
rect 148980 327570 149008 328442
rect 148856 327542 149008 327570
rect 149164 327570 149192 335310
rect 150360 327842 150388 340847
rect 151096 329089 151124 369174
rect 151174 356688 151230 356697
rect 151174 356623 151230 356632
rect 151082 329080 151138 329089
rect 151082 329015 151138 329024
rect 150314 327814 150388 327842
rect 149164 327542 149592 327570
rect 150314 327556 150342 327814
rect 150714 327584 150770 327593
rect 151188 327570 151216 356623
rect 152476 355473 152504 458798
rect 161480 452736 161532 452742
rect 161480 452678 161532 452684
rect 157340 439544 157392 439550
rect 157340 439486 157392 439492
rect 155316 358080 155368 358086
rect 155316 358022 155368 358028
rect 152462 355464 152518 355473
rect 152462 355399 152518 355408
rect 154672 352572 154724 352578
rect 154672 352514 154724 352520
rect 153842 347032 153898 347041
rect 153842 346967 153898 346976
rect 153856 335354 153884 346967
rect 153934 335608 153990 335617
rect 153934 335543 153990 335552
rect 153672 335326 153884 335354
rect 153672 328681 153700 335326
rect 153658 328672 153714 328681
rect 153658 328607 153714 328616
rect 151726 328536 151782 328545
rect 151726 328471 151782 328480
rect 151740 327826 151768 328471
rect 151728 327820 151780 327826
rect 151728 327762 151780 327768
rect 152830 327584 152886 327593
rect 150770 327542 151216 327570
rect 152536 327542 152830 327570
rect 150714 327519 150770 327528
rect 153672 327570 153700 328607
rect 153948 327758 153976 335543
rect 154304 329860 154356 329866
rect 154304 329802 154356 329808
rect 154580 329860 154632 329866
rect 154580 329802 154632 329808
rect 153936 327752 153988 327758
rect 153936 327694 153988 327700
rect 153272 327542 153700 327570
rect 152830 327519 152886 327528
rect 154316 327146 154344 329802
rect 154592 327842 154620 329802
rect 154546 327814 154620 327842
rect 154546 327556 154574 327814
rect 154394 327312 154450 327321
rect 154394 327247 154450 327256
rect 154408 327214 154436 327247
rect 154396 327208 154448 327214
rect 154396 327150 154448 327156
rect 154304 327140 154356 327146
rect 154304 327082 154356 327088
rect 152096 327072 152148 327078
rect 151800 327020 152096 327026
rect 154396 327072 154448 327078
rect 151800 327014 152148 327020
rect 153106 327040 153162 327049
rect 142894 326975 142950 326984
rect 147404 327004 147456 327010
rect 76564 326946 76616 326952
rect 151800 326998 152136 327014
rect 153106 326975 153162 326984
rect 154394 327040 154396 327049
rect 154448 327040 154450 327049
rect 154394 326975 154450 326984
rect 147404 326946 147456 326952
rect 153120 326942 153148 326975
rect 69572 326936 69624 326942
rect 69572 326878 69624 326884
rect 153108 326936 153160 326942
rect 154304 326936 154356 326942
rect 153108 326878 153160 326884
rect 154008 326884 154304 326890
rect 154008 326878 154356 326884
rect 154008 326862 154344 326878
rect 68650 326224 68706 326233
rect 68650 326159 68706 326168
rect 68284 320884 68336 320890
rect 68284 320826 68336 320832
rect 67744 316006 67864 316034
rect 67638 309088 67694 309097
rect 67638 309023 67694 309032
rect 67652 308446 67680 309023
rect 67640 308440 67692 308446
rect 67640 308382 67692 308388
rect 67546 298480 67602 298489
rect 67546 298415 67602 298424
rect 67546 295216 67602 295225
rect 67546 295151 67602 295160
rect 67560 294030 67588 295151
rect 67548 294024 67600 294030
rect 67548 293966 67600 293972
rect 67454 281616 67510 281625
rect 67454 281551 67510 281560
rect 67362 278352 67418 278361
rect 67362 278287 67418 278296
rect 67362 275360 67418 275369
rect 67362 275295 67418 275304
rect 67086 274272 67142 274281
rect 67086 274207 67142 274216
rect 66994 273184 67050 273193
rect 66994 273119 67050 273128
rect 67008 271998 67036 273119
rect 66996 271992 67048 271998
rect 66996 271934 67048 271940
rect 66904 267028 66956 267034
rect 66904 266970 66956 266976
rect 66810 265840 66866 265849
rect 66810 265775 66866 265784
rect 66824 264994 66852 265775
rect 66812 264988 66864 264994
rect 66812 264930 66864 264936
rect 66810 264752 66866 264761
rect 66810 264687 66866 264696
rect 66444 264240 66496 264246
rect 66444 264182 66496 264188
rect 66456 263673 66484 264182
rect 66824 263702 66852 264687
rect 66812 263696 66864 263702
rect 66442 263664 66498 263673
rect 66812 263638 66864 263644
rect 66442 263599 66498 263608
rect 66810 262576 66866 262585
rect 66810 262511 66866 262520
rect 66824 262274 66852 262511
rect 66812 262268 66864 262274
rect 66812 262210 66864 262216
rect 66810 261488 66866 261497
rect 66810 261423 66866 261432
rect 66824 260914 66852 261423
rect 66812 260908 66864 260914
rect 66812 260850 66864 260856
rect 66810 258496 66866 258505
rect 66810 258431 66866 258440
rect 66352 258188 66404 258194
rect 66352 258130 66404 258136
rect 66364 258058 66392 258130
rect 66824 258126 66852 258431
rect 66812 258120 66864 258126
rect 67100 258074 67128 274207
rect 66812 258062 66864 258068
rect 66352 258052 66404 258058
rect 66352 257994 66404 258000
rect 67008 258046 67128 258074
rect 66442 257408 66498 257417
rect 66442 257343 66498 257352
rect 66456 256766 66484 257343
rect 66444 256760 66496 256766
rect 66444 256702 66496 256708
rect 67008 256057 67036 258046
rect 66994 256048 67050 256057
rect 66994 255983 67050 255992
rect 66442 255232 66498 255241
rect 66442 255167 66498 255176
rect 66456 253978 66484 255167
rect 66444 253972 66496 253978
rect 66444 253914 66496 253920
rect 66626 253056 66682 253065
rect 66626 252991 66682 253000
rect 66640 252686 66668 252991
rect 66628 252680 66680 252686
rect 66628 252622 66680 252628
rect 66810 248976 66866 248985
rect 66810 248911 66866 248920
rect 66824 248470 66852 248911
rect 66812 248464 66864 248470
rect 66812 248406 66864 248412
rect 66810 247888 66866 247897
rect 66810 247823 66866 247832
rect 66824 247110 66852 247823
rect 66812 247104 66864 247110
rect 66812 247046 66864 247052
rect 67270 246800 67326 246809
rect 67270 246735 67326 246744
rect 67180 244928 67232 244934
rect 67180 244870 67232 244876
rect 67192 244633 67220 244870
rect 67178 244624 67234 244633
rect 67178 244559 67234 244568
rect 67178 241360 67234 241369
rect 67178 241295 67234 241304
rect 67192 204270 67220 241295
rect 67284 221513 67312 246735
rect 67376 238066 67404 275295
rect 67468 240854 67496 281551
rect 67546 260400 67602 260409
rect 67546 260335 67602 260344
rect 67456 240848 67508 240854
rect 67456 240790 67508 240796
rect 67364 238060 67416 238066
rect 67364 238002 67416 238008
rect 67270 221504 67326 221513
rect 67270 221439 67326 221448
rect 67180 204264 67232 204270
rect 67180 204206 67232 204212
rect 66166 202872 66222 202881
rect 66166 202807 66222 202816
rect 67560 189038 67588 260335
rect 67652 233209 67680 308382
rect 67744 306921 67772 316006
rect 67730 306912 67786 306921
rect 67730 306847 67786 306856
rect 154684 277001 154712 352514
rect 155224 351212 155276 351218
rect 155224 351154 155276 351160
rect 154856 327140 154908 327146
rect 154856 327082 154908 327088
rect 154868 326913 154896 327082
rect 154854 326904 154910 326913
rect 154854 326839 154910 326848
rect 154764 307760 154816 307766
rect 154764 307702 154816 307708
rect 154776 306406 154804 307702
rect 154764 306400 154816 306406
rect 154764 306342 154816 306348
rect 154670 276992 154726 277001
rect 154670 276927 154726 276936
rect 154776 264761 154804 306342
rect 155236 296714 155264 351154
rect 155328 307766 155356 358022
rect 155868 357536 155920 357542
rect 155868 357478 155920 357484
rect 155880 356697 155908 357478
rect 155866 356688 155922 356697
rect 155866 356623 155922 356632
rect 156142 349752 156198 349761
rect 156142 349687 156198 349696
rect 156052 348424 156104 348430
rect 156052 348366 156104 348372
rect 155958 345672 156014 345681
rect 155958 345607 156014 345616
rect 155868 326936 155920 326942
rect 155868 326878 155920 326884
rect 155880 320958 155908 326878
rect 155868 320952 155920 320958
rect 155868 320894 155920 320900
rect 155972 318073 156000 345607
rect 155958 318064 156014 318073
rect 155958 317999 156014 318008
rect 155316 307760 155368 307766
rect 155316 307702 155368 307708
rect 154868 296686 155264 296714
rect 154868 295633 154896 296686
rect 154854 295624 154910 295633
rect 154854 295559 154910 295568
rect 154762 264752 154818 264761
rect 154762 264687 154818 264696
rect 154868 262041 154896 295559
rect 155222 290456 155278 290465
rect 155222 290391 155278 290400
rect 154854 262032 154910 262041
rect 154854 261967 154910 261976
rect 68098 258768 68154 258777
rect 68098 258703 68154 258712
rect 68112 258058 68140 258703
rect 68100 258052 68152 258058
rect 68100 257994 68152 258000
rect 67914 250880 67970 250889
rect 67914 250815 67970 250824
rect 67730 250064 67786 250073
rect 67730 249999 67786 250008
rect 67638 233200 67694 233209
rect 67638 233135 67694 233144
rect 67744 226137 67772 249999
rect 67928 238134 67956 250815
rect 155236 242078 155264 290391
rect 155316 276684 155368 276690
rect 155316 276626 155368 276632
rect 71044 242072 71096 242078
rect 152464 242072 152516 242078
rect 135994 242040 136050 242049
rect 71044 242014 71096 242020
rect 69754 241904 69810 241913
rect 69754 241839 69756 241848
rect 69808 241839 69810 241848
rect 69756 241810 69808 241816
rect 69662 241768 69718 241777
rect 69662 241703 69718 241712
rect 68816 241590 68968 241618
rect 68940 239562 68968 241590
rect 69032 241590 69368 241618
rect 68928 239556 68980 239562
rect 68928 239498 68980 239504
rect 67916 238128 67968 238134
rect 67916 238070 67968 238076
rect 67730 226128 67786 226137
rect 67730 226063 67786 226072
rect 69032 209778 69060 241590
rect 69676 216481 69704 241703
rect 70104 241590 70256 241618
rect 70228 239494 70256 241590
rect 70412 241590 70840 241618
rect 70308 239556 70360 239562
rect 70308 239498 70360 239504
rect 70216 239488 70268 239494
rect 70216 239430 70268 239436
rect 70320 238649 70348 239498
rect 70306 238640 70362 238649
rect 70306 238575 70362 238584
rect 69662 216472 69718 216481
rect 69662 216407 69718 216416
rect 70412 210458 70440 241590
rect 71056 230450 71084 242014
rect 135272 241998 135994 242026
rect 72424 241868 72476 241874
rect 72424 241810 72476 241816
rect 71576 241590 71728 241618
rect 71700 240417 71728 241590
rect 71792 241590 72312 241618
rect 71686 240408 71742 240417
rect 71686 240343 71742 240352
rect 71792 234433 71820 241590
rect 71778 234424 71834 234433
rect 71778 234359 71834 234368
rect 71044 230444 71096 230450
rect 71044 230386 71096 230392
rect 70400 210452 70452 210458
rect 70400 210394 70452 210400
rect 69020 209772 69072 209778
rect 69020 209714 69072 209720
rect 72436 204950 72464 241810
rect 73048 241590 73108 241618
rect 72424 204944 72476 204950
rect 72424 204886 72476 204892
rect 73080 196625 73108 241590
rect 73172 241590 73784 241618
rect 74520 241590 74580 241618
rect 75072 241590 75408 241618
rect 73172 238513 73200 241590
rect 74446 239592 74502 239601
rect 74446 239527 74502 239536
rect 74460 238814 74488 239527
rect 74448 238808 74500 238814
rect 74448 238750 74500 238756
rect 73158 238504 73214 238513
rect 73158 238439 73214 238448
rect 73802 237960 73858 237969
rect 73802 237895 73858 237904
rect 73816 220697 73844 237895
rect 73802 220688 73858 220697
rect 73802 220623 73858 220632
rect 74460 197334 74488 238750
rect 74552 205601 74580 241590
rect 75380 239970 75408 241590
rect 75472 241590 75808 241618
rect 76544 241590 77156 241618
rect 77280 241590 77340 241618
rect 75368 239964 75420 239970
rect 75368 239906 75420 239912
rect 75472 238814 75500 241590
rect 75828 239964 75880 239970
rect 75828 239906 75880 239912
rect 75460 238808 75512 238814
rect 75460 238750 75512 238756
rect 75184 235340 75236 235346
rect 75184 235282 75236 235288
rect 75196 213897 75224 235282
rect 75840 220794 75868 239906
rect 75828 220788 75880 220794
rect 75828 220730 75880 220736
rect 75182 213888 75238 213897
rect 75182 213823 75238 213832
rect 77128 212401 77156 241590
rect 77206 239456 77262 239465
rect 77312 239442 77340 241590
rect 77262 239414 77340 239442
rect 77206 239391 77262 239400
rect 77312 238754 77340 239414
rect 77220 238726 77340 238754
rect 77404 241590 78016 241618
rect 78752 241590 79088 241618
rect 79488 241590 79916 241618
rect 80224 241590 80560 241618
rect 80776 241590 81388 241618
rect 81512 241590 81572 241618
rect 77114 212392 77170 212401
rect 77114 212327 77170 212336
rect 74538 205592 74594 205601
rect 74538 205527 74594 205536
rect 77220 201482 77248 238726
rect 77404 214849 77432 241590
rect 79060 239426 79088 241590
rect 79048 239420 79100 239426
rect 79048 239362 79100 239368
rect 79324 238128 79376 238134
rect 79324 238070 79376 238076
rect 79336 226001 79364 238070
rect 79888 229022 79916 241590
rect 80532 239426 80560 241590
rect 81256 240848 81308 240854
rect 81256 240790 81308 240796
rect 79968 239420 80020 239426
rect 79968 239362 80020 239368
rect 80520 239420 80572 239426
rect 80520 239362 80572 239368
rect 79876 229016 79928 229022
rect 79876 228958 79928 228964
rect 79322 225992 79378 226001
rect 79322 225927 79378 225936
rect 77390 214840 77446 214849
rect 77390 214775 77446 214784
rect 77208 201476 77260 201482
rect 77208 201418 77260 201424
rect 74448 197328 74500 197334
rect 74448 197270 74500 197276
rect 73066 196616 73122 196625
rect 73066 196551 73122 196560
rect 67548 189032 67600 189038
rect 67548 188974 67600 188980
rect 79980 185609 80008 239362
rect 81268 236706 81296 240790
rect 81256 236700 81308 236706
rect 81256 236642 81308 236648
rect 81360 188329 81388 241590
rect 81544 239562 81572 241590
rect 81636 241590 82248 241618
rect 81532 239556 81584 239562
rect 81532 239498 81584 239504
rect 81636 216646 81664 241590
rect 82970 241505 82998 241604
rect 83108 241590 83720 241618
rect 84456 241590 84792 241618
rect 85192 241590 85528 241618
rect 85928 241590 86080 241618
rect 82956 241496 83012 241505
rect 82956 241431 83012 241440
rect 82728 239556 82780 239562
rect 82728 239498 82780 239504
rect 82740 224262 82768 239498
rect 83108 238746 83136 241590
rect 84106 241496 84162 241505
rect 84106 241431 84162 241440
rect 83096 238740 83148 238746
rect 83096 238682 83148 238688
rect 84120 226273 84148 241431
rect 84764 239465 84792 241590
rect 84750 239456 84806 239465
rect 84750 239391 84806 239400
rect 84106 226264 84162 226273
rect 84106 226199 84162 226208
rect 82728 224256 82780 224262
rect 82728 224198 82780 224204
rect 81624 216640 81676 216646
rect 81624 216582 81676 216588
rect 85500 200977 85528 241590
rect 86052 240106 86080 241590
rect 86144 241590 86480 241618
rect 86972 241590 87216 241618
rect 87952 241590 88288 241618
rect 88688 241590 89024 241618
rect 89424 241590 89668 241618
rect 90160 241590 90496 241618
rect 90896 241590 91048 241618
rect 91632 241590 91968 241618
rect 92184 241590 92336 241618
rect 86040 240100 86092 240106
rect 86040 240042 86092 240048
rect 86144 238754 86172 241590
rect 86868 240100 86920 240106
rect 86868 240042 86920 240048
rect 85592 238726 86172 238754
rect 85592 207670 85620 238726
rect 85580 207664 85632 207670
rect 85580 207606 85632 207612
rect 86880 204921 86908 240042
rect 86972 223582 87000 241590
rect 86960 223576 87012 223582
rect 86960 223518 87012 223524
rect 86866 204912 86922 204921
rect 86866 204847 86922 204856
rect 85486 200968 85542 200977
rect 85486 200903 85542 200912
rect 88260 195265 88288 241590
rect 88996 239970 89024 241590
rect 88984 239964 89036 239970
rect 88984 239906 89036 239912
rect 89536 239964 89588 239970
rect 89536 239906 89588 239912
rect 88984 239420 89036 239426
rect 88984 239362 89036 239368
rect 88996 220833 89024 239362
rect 88982 220824 89038 220833
rect 88982 220759 89038 220768
rect 89548 206990 89576 239906
rect 89536 206984 89588 206990
rect 89536 206926 89588 206932
rect 88246 195256 88302 195265
rect 88246 195191 88302 195200
rect 89640 189689 89668 241590
rect 90468 239970 90496 241590
rect 90456 239964 90508 239970
rect 90456 239906 90508 239912
rect 90916 239964 90968 239970
rect 90916 239906 90968 239912
rect 90928 228313 90956 239906
rect 90914 228304 90970 228313
rect 90914 228239 90970 228248
rect 89626 189680 89682 189689
rect 89626 189615 89682 189624
rect 81346 188320 81402 188329
rect 81346 188255 81402 188264
rect 91020 185638 91048 241590
rect 91940 240106 91968 241590
rect 91928 240100 91980 240106
rect 91928 240042 91980 240048
rect 92308 217297 92336 241590
rect 92492 241590 92920 241618
rect 93656 241590 93808 241618
rect 92388 240100 92440 240106
rect 92388 240042 92440 240048
rect 92294 217288 92350 217297
rect 92294 217223 92350 217232
rect 92400 209710 92428 240042
rect 92492 231810 92520 241590
rect 92480 231804 92532 231810
rect 92480 231746 92532 231752
rect 92492 231130 92520 231746
rect 92480 231124 92532 231130
rect 92480 231066 92532 231072
rect 93124 231124 93176 231130
rect 93124 231066 93176 231072
rect 92388 209704 92440 209710
rect 92388 209646 92440 209652
rect 93136 194546 93164 231066
rect 93124 194540 93176 194546
rect 93124 194482 93176 194488
rect 93780 186969 93808 241590
rect 93872 241590 94392 241618
rect 95128 241590 95188 241618
rect 93872 231810 93900 241590
rect 93860 231804 93912 231810
rect 93860 231746 93912 231752
rect 94504 231804 94556 231810
rect 94504 231746 94556 231752
rect 94516 220726 94544 231746
rect 94504 220720 94556 220726
rect 94504 220662 94556 220668
rect 95160 199345 95188 241590
rect 95252 241590 95864 241618
rect 96600 241590 96936 241618
rect 97336 241590 97672 241618
rect 97888 241590 97948 241618
rect 98624 241590 99236 241618
rect 99360 241590 99420 241618
rect 95252 212537 95280 241590
rect 96908 240038 96936 241590
rect 96896 240032 96948 240038
rect 96896 239974 96948 239980
rect 97644 238754 97672 241590
rect 97644 238726 97856 238754
rect 97264 229764 97316 229770
rect 97264 229706 97316 229712
rect 97276 222154 97304 229706
rect 97264 222148 97316 222154
rect 97264 222090 97316 222096
rect 95238 212528 95294 212537
rect 95238 212463 95294 212472
rect 97828 202774 97856 238726
rect 97816 202768 97868 202774
rect 97816 202710 97868 202716
rect 95146 199336 95202 199345
rect 95146 199271 95202 199280
rect 97920 191146 97948 241590
rect 99208 238754 99236 241590
rect 99392 239562 99420 241590
rect 99484 241590 100096 241618
rect 100832 241590 101168 241618
rect 101568 241590 102088 241618
rect 102304 241590 102640 241618
rect 103040 241590 103468 241618
rect 99380 239556 99432 239562
rect 99380 239498 99432 239504
rect 99208 238726 99328 238754
rect 98552 238060 98604 238066
rect 98552 238002 98604 238008
rect 98564 233238 98592 238002
rect 98552 233232 98604 233238
rect 98552 233174 98604 233180
rect 99300 213353 99328 238726
rect 99484 219434 99512 241590
rect 101140 240106 101168 241590
rect 101128 240100 101180 240106
rect 101128 240042 101180 240048
rect 101956 240100 102008 240106
rect 101956 240042 102008 240048
rect 101496 240032 101548 240038
rect 101496 239974 101548 239980
rect 100668 239556 100720 239562
rect 100668 239498 100720 239504
rect 99472 219428 99524 219434
rect 99472 219370 99524 219376
rect 99286 213344 99342 213353
rect 99286 213279 99342 213288
rect 100680 193866 100708 239498
rect 101508 238678 101536 239974
rect 101496 238672 101548 238678
rect 101496 238614 101548 238620
rect 101968 207777 101996 240042
rect 101954 207768 102010 207777
rect 101954 207703 102010 207712
rect 102060 200841 102088 241590
rect 102612 239290 102640 241590
rect 102600 239284 102652 239290
rect 102600 239226 102652 239232
rect 103336 239284 103388 239290
rect 103336 239226 103388 239232
rect 103348 231849 103376 239226
rect 103334 231840 103390 231849
rect 103334 231775 103390 231784
rect 103440 216510 103468 241590
rect 103532 241590 103592 241618
rect 104328 241590 104848 241618
rect 103532 237289 103560 241590
rect 103612 240780 103664 240786
rect 103612 240722 103664 240728
rect 103518 237280 103574 237289
rect 103518 237215 103574 237224
rect 103624 235958 103652 240722
rect 103612 235952 103664 235958
rect 103612 235894 103664 235900
rect 104164 233912 104216 233918
rect 104164 233854 104216 233860
rect 104176 220114 104204 233854
rect 104164 220108 104216 220114
rect 104164 220050 104216 220056
rect 103428 216504 103480 216510
rect 103428 216446 103480 216452
rect 104820 211041 104848 241590
rect 105050 241466 105078 241604
rect 105464 241590 105800 241618
rect 106536 241590 106872 241618
rect 107272 241590 107516 241618
rect 108008 241590 108252 241618
rect 105038 241460 105090 241466
rect 105038 241402 105090 241408
rect 105464 238754 105492 241590
rect 106844 239834 106872 241590
rect 106832 239828 106884 239834
rect 106832 239770 106884 239776
rect 106922 239456 106978 239465
rect 106922 239391 106978 239400
rect 104912 238726 105492 238754
rect 104912 213217 104940 238726
rect 106936 227730 106964 239391
rect 106924 227724 106976 227730
rect 106924 227666 106976 227672
rect 107488 224777 107516 241590
rect 107568 239828 107620 239834
rect 107568 239770 107620 239776
rect 107474 224768 107530 224777
rect 107474 224703 107530 224712
rect 107580 214713 107608 239770
rect 108224 239426 108252 241590
rect 108408 241590 108744 241618
rect 109296 241590 109632 241618
rect 110032 241590 110276 241618
rect 110768 241590 111104 241618
rect 111504 241590 111656 241618
rect 112240 241590 112576 241618
rect 112976 241590 113128 241618
rect 108304 239488 108356 239494
rect 108304 239430 108356 239436
rect 108212 239420 108264 239426
rect 108212 239362 108264 239368
rect 107752 239284 107804 239290
rect 107752 239226 107804 239232
rect 107764 233918 107792 239226
rect 107752 233912 107804 233918
rect 107752 233854 107804 233860
rect 108316 230353 108344 239430
rect 108408 239290 108436 241590
rect 109604 239834 109632 241590
rect 109592 239828 109644 239834
rect 109592 239770 109644 239776
rect 110248 239494 110276 241590
rect 110328 239828 110380 239834
rect 110328 239770 110380 239776
rect 110236 239488 110288 239494
rect 110236 239430 110288 239436
rect 108396 239284 108448 239290
rect 108396 239226 108448 239232
rect 108302 230344 108358 230353
rect 108302 230279 108358 230288
rect 107566 214704 107622 214713
rect 107566 214639 107622 214648
rect 104898 213208 104954 213217
rect 104898 213143 104954 213152
rect 104806 211032 104862 211041
rect 104806 210967 104862 210976
rect 110340 206922 110368 239770
rect 111076 239290 111104 241590
rect 111064 239284 111116 239290
rect 111064 239226 111116 239232
rect 110328 206916 110380 206922
rect 110328 206858 110380 206864
rect 102046 200832 102102 200841
rect 102046 200767 102102 200776
rect 111628 199442 111656 241590
rect 112548 239465 112576 241590
rect 112534 239456 112590 239465
rect 112534 239391 112590 239400
rect 111708 239284 111760 239290
rect 111708 239226 111760 239232
rect 111616 199436 111668 199442
rect 111616 199378 111668 199384
rect 100668 193860 100720 193866
rect 100668 193802 100720 193808
rect 97908 191140 97960 191146
rect 97908 191082 97960 191088
rect 106188 190528 106240 190534
rect 106188 190470 106240 190476
rect 93766 186960 93822 186969
rect 93766 186895 93822 186904
rect 91008 185632 91060 185638
rect 79966 185600 80022 185609
rect 91008 185574 91060 185580
rect 79966 185535 80022 185544
rect 104806 183832 104862 183841
rect 104806 183767 104862 183776
rect 101954 183696 102010 183705
rect 101954 183631 102010 183640
rect 99470 182200 99526 182209
rect 99470 182135 99526 182144
rect 99484 176769 99512 182135
rect 101968 177585 101996 183631
rect 103336 182300 103388 182306
rect 103336 182242 103388 182248
rect 101954 177576 102010 177585
rect 101954 177511 102010 177520
rect 102048 176928 102100 176934
rect 102048 176870 102100 176876
rect 102060 176769 102088 176870
rect 103348 176769 103376 182242
rect 104820 177585 104848 183767
rect 105450 179480 105506 179489
rect 105450 179415 105506 179424
rect 104806 177576 104862 177585
rect 104806 177511 104862 177520
rect 105464 176934 105492 179415
rect 106200 177585 106228 190470
rect 111720 188465 111748 239226
rect 113100 211886 113128 241590
rect 113192 241590 113712 241618
rect 114448 241590 114508 241618
rect 115000 241590 115336 241618
rect 113192 232937 113220 241590
rect 113178 232928 113234 232937
rect 113178 232863 113234 232872
rect 113088 211880 113140 211886
rect 113088 211822 113140 211828
rect 114480 204105 114508 241590
rect 115308 240106 115336 241590
rect 115400 241590 115736 241618
rect 116472 241590 116808 241618
rect 117208 241590 117268 241618
rect 117944 241590 118372 241618
rect 118680 241590 118832 241618
rect 115296 240100 115348 240106
rect 115296 240042 115348 240048
rect 115400 240038 115428 241590
rect 115848 240100 115900 240106
rect 115848 240042 115900 240048
rect 114652 240032 114704 240038
rect 114652 239974 114704 239980
rect 115388 240032 115440 240038
rect 115388 239974 115440 239980
rect 114664 233986 114692 239974
rect 115204 239488 115256 239494
rect 115204 239430 115256 239436
rect 114652 233980 114704 233986
rect 114652 233922 114704 233928
rect 114466 204096 114522 204105
rect 114466 204031 114522 204040
rect 115216 198694 115244 239430
rect 115204 198688 115256 198694
rect 115204 198630 115256 198636
rect 111706 188456 111762 188465
rect 111706 188391 111762 188400
rect 115860 186998 115888 240042
rect 116780 240038 116808 241590
rect 116768 240032 116820 240038
rect 116768 239974 116820 239980
rect 117240 239873 117268 241590
rect 117226 239864 117282 239873
rect 117226 239799 117282 239808
rect 118344 238754 118372 241590
rect 118804 240106 118832 241590
rect 118896 241590 119416 241618
rect 120092 241590 120152 241618
rect 120704 241590 121040 241618
rect 121440 241590 121776 241618
rect 122176 241590 122696 241618
rect 118792 240100 118844 240106
rect 118792 240042 118844 240048
rect 118344 238726 118648 238754
rect 118620 202201 118648 238726
rect 118896 227662 118924 241590
rect 119988 240100 120040 240106
rect 119988 240042 120040 240048
rect 118884 227656 118936 227662
rect 118884 227598 118936 227604
rect 118896 222057 118924 227598
rect 120000 223514 120028 240042
rect 120092 235793 120120 241590
rect 121012 240786 121040 241590
rect 121000 240780 121052 240786
rect 121000 240722 121052 240728
rect 121748 240106 121776 241590
rect 121736 240100 121788 240106
rect 121736 240042 121788 240048
rect 120078 235784 120134 235793
rect 120078 235719 120134 235728
rect 119988 223508 120040 223514
rect 119988 223450 120040 223456
rect 118882 222048 118938 222057
rect 118882 221983 118938 221992
rect 122668 218754 122696 241590
rect 122852 241590 122912 241618
rect 123036 241590 123648 241618
rect 124384 241590 124720 241618
rect 125120 241590 125456 241618
rect 125856 241590 126192 241618
rect 126408 241590 126928 241618
rect 122748 240100 122800 240106
rect 122748 240042 122800 240048
rect 122656 218748 122708 218754
rect 122656 218690 122708 218696
rect 118606 202192 118662 202201
rect 118606 202127 118662 202136
rect 122760 195294 122788 240042
rect 122852 217938 122880 241590
rect 123036 226302 123064 241590
rect 124692 240106 124720 241590
rect 124680 240100 124732 240106
rect 124680 240042 124732 240048
rect 124312 240032 124364 240038
rect 124312 239974 124364 239980
rect 124324 238377 124352 239974
rect 124310 238368 124366 238377
rect 124310 238303 124366 238312
rect 124588 235272 124640 235278
rect 124588 235214 124640 235220
rect 124600 233170 124628 235214
rect 124588 233164 124640 233170
rect 124588 233106 124640 233112
rect 123484 232552 123536 232558
rect 123484 232494 123536 232500
rect 123496 228993 123524 232494
rect 123482 228984 123538 228993
rect 123482 228919 123538 228928
rect 123024 226296 123076 226302
rect 123024 226238 123076 226244
rect 122840 217932 122892 217938
rect 122840 217874 122892 217880
rect 125428 205630 125456 241590
rect 125508 240100 125560 240106
rect 125508 240042 125560 240048
rect 125416 205624 125468 205630
rect 125416 205566 125468 205572
rect 125520 205465 125548 240042
rect 126164 240009 126192 241590
rect 126150 240000 126206 240009
rect 126150 239935 126206 239944
rect 126796 235272 126848 235278
rect 126796 235214 126848 235220
rect 126808 209681 126836 235214
rect 126900 210905 126928 241590
rect 127084 241590 127144 241618
rect 127880 241590 128308 241618
rect 128616 241590 128952 241618
rect 129352 241590 129596 241618
rect 130088 241590 130424 241618
rect 130824 241590 131068 241618
rect 131560 241590 131896 241618
rect 132112 241590 132448 241618
rect 132848 241590 133184 241618
rect 133584 241590 133828 241618
rect 134320 241590 134656 241618
rect 127084 237153 127112 241590
rect 127070 237144 127126 237153
rect 127070 237079 127126 237088
rect 126886 210896 126942 210905
rect 126886 210831 126942 210840
rect 126794 209672 126850 209681
rect 126794 209607 126850 209616
rect 125506 205456 125562 205465
rect 125506 205391 125562 205400
rect 126808 202842 126836 209607
rect 128280 206961 128308 241590
rect 128924 240106 128952 241590
rect 128912 240100 128964 240106
rect 128912 240042 128964 240048
rect 128358 236600 128414 236609
rect 128358 236535 128414 236544
rect 128372 231674 128400 236535
rect 128360 231668 128412 231674
rect 128360 231610 128412 231616
rect 129568 227361 129596 241590
rect 130396 240106 130424 241590
rect 129648 240100 129700 240106
rect 129648 240042 129700 240048
rect 130384 240100 130436 240106
rect 130384 240042 130436 240048
rect 130936 240100 130988 240106
rect 130936 240042 130988 240048
rect 129554 227352 129610 227361
rect 129554 227287 129610 227296
rect 128266 206952 128322 206961
rect 128266 206887 128322 206896
rect 126796 202836 126848 202842
rect 126796 202778 126848 202784
rect 129660 202337 129688 240042
rect 130948 224942 130976 240042
rect 130936 224936 130988 224942
rect 130936 224878 130988 224884
rect 131040 210526 131068 241590
rect 131868 239290 131896 241590
rect 131856 239284 131908 239290
rect 131856 239226 131908 239232
rect 132316 239284 132368 239290
rect 132316 239226 132368 239232
rect 132328 215286 132356 239226
rect 132316 215280 132368 215286
rect 132316 215222 132368 215228
rect 131028 210520 131080 210526
rect 131028 210462 131080 210468
rect 129646 202328 129702 202337
rect 129646 202263 129702 202272
rect 122748 195288 122800 195294
rect 122748 195230 122800 195236
rect 132420 192506 132448 241590
rect 133156 239018 133184 241590
rect 133144 239012 133196 239018
rect 133144 238954 133196 238960
rect 133696 239012 133748 239018
rect 133696 238954 133748 238960
rect 133708 198121 133736 238954
rect 133694 198112 133750 198121
rect 133694 198047 133750 198056
rect 133800 193905 133828 241590
rect 134628 239018 134656 241590
rect 134720 241590 135056 241618
rect 134616 239012 134668 239018
rect 134616 238954 134668 238960
rect 134720 238754 134748 241590
rect 135168 239012 135220 239018
rect 135168 238954 135220 238960
rect 133892 238726 134748 238754
rect 133892 221474 133920 238726
rect 135180 230217 135208 238954
rect 135272 235278 135300 241998
rect 135994 241975 136050 241984
rect 138202 242040 138258 242049
rect 150254 242040 150310 242049
rect 138258 241998 138552 242026
rect 149960 241998 150254 242026
rect 138202 241975 138258 241984
rect 152464 242014 152516 242020
rect 155224 242072 155276 242078
rect 155224 242014 155276 242020
rect 150254 241975 150310 241984
rect 136528 241590 136588 241618
rect 135260 235272 135312 235278
rect 135260 235214 135312 235220
rect 135994 234696 136050 234705
rect 135994 234631 136050 234640
rect 136008 231810 136036 234631
rect 135996 231804 136048 231810
rect 135996 231746 136048 231752
rect 136560 231742 136588 241590
rect 136652 241590 137264 241618
rect 137816 241590 137968 241618
rect 136652 237386 136680 241590
rect 136640 237380 136692 237386
rect 136640 237322 136692 237328
rect 136652 236026 136680 237322
rect 136640 236020 136692 236026
rect 136640 235962 136692 235968
rect 137284 236020 137336 236026
rect 137284 235962 137336 235968
rect 136548 231736 136600 231742
rect 136548 231678 136600 231684
rect 135166 230208 135222 230217
rect 135166 230143 135222 230152
rect 137296 223417 137324 235962
rect 137940 230382 137968 241590
rect 138216 238754 138244 241975
rect 139288 241590 139348 241618
rect 140024 241590 140544 241618
rect 140760 241590 140820 241618
rect 141496 241590 142108 241618
rect 138124 238726 138244 238754
rect 138124 237386 138152 238726
rect 138112 237380 138164 237386
rect 138112 237322 138164 237328
rect 139214 234016 139270 234025
rect 139214 233951 139216 233960
rect 139268 233951 139270 233960
rect 139216 233922 139268 233928
rect 137928 230376 137980 230382
rect 137928 230318 137980 230324
rect 137282 223408 137338 223417
rect 137282 223343 137338 223352
rect 133880 221468 133932 221474
rect 133880 221410 133932 221416
rect 139228 195945 139256 233922
rect 139320 200122 139348 241590
rect 140516 238754 140544 241590
rect 140516 238726 140728 238754
rect 139400 233980 139452 233986
rect 139400 233922 139452 233928
rect 139412 233170 139440 233922
rect 139400 233164 139452 233170
rect 139400 233106 139452 233112
rect 140700 207641 140728 238726
rect 140792 233073 140820 241590
rect 140778 233064 140834 233073
rect 140778 232999 140834 233008
rect 142080 227662 142108 241590
rect 142172 241590 142232 241618
rect 142968 241590 143488 241618
rect 143704 241590 144040 241618
rect 144256 241590 144868 241618
rect 144992 241590 145328 241618
rect 145728 241590 146248 241618
rect 142068 227656 142120 227662
rect 142068 227598 142120 227604
rect 142172 220561 142200 241590
rect 143460 231713 143488 241590
rect 144012 239290 144040 241590
rect 144000 239284 144052 239290
rect 144000 239226 144052 239232
rect 144736 239284 144788 239290
rect 144736 239226 144788 239232
rect 143446 231704 143502 231713
rect 143446 231639 143502 231648
rect 142158 220552 142214 220561
rect 142158 220487 142214 220496
rect 144748 215218 144776 239226
rect 144736 215212 144788 215218
rect 144736 215154 144788 215160
rect 140686 207632 140742 207641
rect 140686 207567 140742 207576
rect 144840 201414 144868 241590
rect 145300 239154 145328 241590
rect 145288 239148 145340 239154
rect 145288 239090 145340 239096
rect 145932 239148 145984 239154
rect 145932 239090 145984 239096
rect 145944 231577 145972 239090
rect 146024 235476 146076 235482
rect 146024 235418 146076 235424
rect 146036 231674 146064 235418
rect 146220 231826 146248 241590
rect 146404 241590 146464 241618
rect 147200 241590 147628 241618
rect 147936 241590 148272 241618
rect 146404 234297 146432 241590
rect 146390 234288 146446 234297
rect 146390 234223 146446 234232
rect 146944 233912 146996 233918
rect 146944 233854 146996 233860
rect 146956 233170 146984 233854
rect 146944 233164 146996 233170
rect 146944 233106 146996 233112
rect 146128 231798 146248 231826
rect 147600 231810 147628 241590
rect 148138 241496 148194 241505
rect 148138 241431 148194 241440
rect 148152 240553 148180 241431
rect 148138 240544 148194 240553
rect 148138 240479 148194 240488
rect 147772 239964 147824 239970
rect 147772 239906 147824 239912
rect 147678 237688 147734 237697
rect 147678 237623 147734 237632
rect 147692 233986 147720 237623
rect 147680 233980 147732 233986
rect 147680 233922 147732 233928
rect 147784 233918 147812 239906
rect 148152 238377 148180 240479
rect 148244 239154 148272 241590
rect 148336 241590 148672 241618
rect 149408 241590 149744 241618
rect 148336 239970 148364 241590
rect 148324 239964 148376 239970
rect 148324 239906 148376 239912
rect 149716 239494 149744 241590
rect 150682 241505 150710 241604
rect 151432 241590 151768 241618
rect 150668 241496 150724 241505
rect 150668 241431 150724 241440
rect 149704 239488 149756 239494
rect 149704 239430 149756 239436
rect 148232 239148 148284 239154
rect 148232 239090 148284 239096
rect 148968 239148 149020 239154
rect 148968 239090 149020 239096
rect 148138 238368 148194 238377
rect 148138 238303 148194 238312
rect 147772 233912 147824 233918
rect 147772 233854 147824 233860
rect 147588 231804 147640 231810
rect 146024 231668 146076 231674
rect 146024 231610 146076 231616
rect 145930 231568 145986 231577
rect 145930 231503 145986 231512
rect 146128 225622 146156 231798
rect 147588 231746 147640 231752
rect 146206 231160 146262 231169
rect 146206 231095 146262 231104
rect 146220 228857 146248 231095
rect 146206 228848 146262 228857
rect 146206 228783 146262 228792
rect 146116 225616 146168 225622
rect 146116 225558 146168 225564
rect 144828 201408 144880 201414
rect 144828 201350 144880 201356
rect 139308 200116 139360 200122
rect 139308 200058 139360 200064
rect 148980 196654 149008 239090
rect 151082 228304 151138 228313
rect 151082 228239 151138 228248
rect 151096 210594 151124 228239
rect 151084 210588 151136 210594
rect 151084 210530 151136 210536
rect 150440 210452 150492 210458
rect 150440 210394 150492 210400
rect 150452 204202 150480 210394
rect 150440 204196 150492 204202
rect 150440 204138 150492 204144
rect 148968 196648 149020 196654
rect 148968 196590 149020 196596
rect 139214 195936 139270 195945
rect 139214 195871 139270 195880
rect 133786 193896 133842 193905
rect 133786 193831 133842 193840
rect 132408 192500 132460 192506
rect 132408 192442 132460 192448
rect 151740 191049 151768 241590
rect 151832 241590 152168 241618
rect 151832 235657 151860 241590
rect 152476 237697 152504 242014
rect 152554 241904 152610 241913
rect 152610 241862 153148 241890
rect 152554 241839 152610 241848
rect 152462 237688 152518 237697
rect 152462 237623 152518 237632
rect 151818 235648 151874 235657
rect 151818 235583 151874 235592
rect 153014 234696 153070 234705
rect 153014 234631 153070 234640
rect 153028 234598 153056 234631
rect 153016 234592 153068 234598
rect 153016 234534 153068 234540
rect 153120 216345 153148 241862
rect 153640 241590 153976 241618
rect 154376 241590 154436 241618
rect 153844 241528 153896 241534
rect 153844 241470 153896 241476
rect 153856 235482 153884 241470
rect 153948 239290 153976 241590
rect 153936 239284 153988 239290
rect 153936 239226 153988 239232
rect 153844 235476 153896 235482
rect 153844 235418 153896 235424
rect 153106 216336 153162 216345
rect 153106 216271 153162 216280
rect 154408 214849 154436 241590
rect 154488 239284 154540 239290
rect 154488 239226 154540 239232
rect 152462 214840 152518 214849
rect 152462 214775 152518 214784
rect 154394 214840 154450 214849
rect 154394 214775 154450 214784
rect 152476 206825 152504 214775
rect 152462 206816 152518 206825
rect 152462 206751 152518 206760
rect 154500 202230 154528 239226
rect 155328 231810 155356 276626
rect 155408 259480 155460 259486
rect 155408 259422 155460 259428
rect 155420 241466 155448 259422
rect 155590 245848 155646 245857
rect 155590 245783 155646 245792
rect 155498 241768 155554 241777
rect 155498 241703 155554 241712
rect 155408 241460 155460 241466
rect 155408 241402 155460 241408
rect 155316 231804 155368 231810
rect 155316 231746 155368 231752
rect 155512 227662 155540 241703
rect 155604 233238 155632 245783
rect 155592 233232 155644 233238
rect 155592 233174 155644 233180
rect 155868 231804 155920 231810
rect 155868 231746 155920 231752
rect 155880 231441 155908 231746
rect 155866 231432 155922 231441
rect 155866 231367 155922 231376
rect 155500 227656 155552 227662
rect 155500 227598 155552 227604
rect 155972 223530 156000 317999
rect 156064 254697 156092 348366
rect 156156 325694 156184 349687
rect 157246 326904 157302 326913
rect 157246 326839 157302 326848
rect 156418 326496 156474 326505
rect 156418 326431 156474 326440
rect 156432 325718 156460 326431
rect 156420 325712 156472 325718
rect 156156 325666 156276 325694
rect 156142 310448 156198 310457
rect 156142 310383 156198 310392
rect 156156 309330 156184 310383
rect 156144 309324 156196 309330
rect 156144 309266 156196 309272
rect 156248 308553 156276 325666
rect 156420 325654 156472 325660
rect 157154 325408 157210 325417
rect 157154 325343 157156 325352
rect 157208 325343 157210 325352
rect 157156 325314 157208 325320
rect 157260 324970 157288 326839
rect 157248 324964 157300 324970
rect 157248 324906 157300 324912
rect 156878 324320 156934 324329
rect 156878 324255 156934 324264
rect 156892 322998 156920 324255
rect 156880 322992 156932 322998
rect 156880 322934 156932 322940
rect 157246 322144 157302 322153
rect 157246 322079 157302 322088
rect 157260 321638 157288 322079
rect 157248 321632 157300 321638
rect 157248 321574 157300 321580
rect 157246 318880 157302 318889
rect 157246 318815 157248 318824
rect 157300 318815 157302 318824
rect 157248 318786 157300 318792
rect 156602 318744 156658 318753
rect 156602 318679 156658 318688
rect 156616 317529 156644 318679
rect 156602 317520 156658 317529
rect 156602 317455 156658 317464
rect 156418 312624 156474 312633
rect 156418 312559 156474 312568
rect 156432 311914 156460 312559
rect 156420 311908 156472 311914
rect 156420 311850 156472 311856
rect 156234 308544 156290 308553
rect 156234 308479 156290 308488
rect 156616 296857 156644 317455
rect 157248 317416 157300 317422
rect 157248 317358 157300 317364
rect 157260 316985 157288 317358
rect 157246 316976 157302 316985
rect 157246 316911 157302 316920
rect 156786 315888 156842 315897
rect 156786 315823 156842 315832
rect 156800 314702 156828 315823
rect 157248 315376 157300 315382
rect 157248 315318 157300 315324
rect 157260 314809 157288 315318
rect 157246 314800 157302 314809
rect 157246 314735 157302 314744
rect 156788 314696 156840 314702
rect 156788 314638 156840 314644
rect 157246 311536 157302 311545
rect 157246 311471 157302 311480
rect 157260 310554 157288 311471
rect 157248 310548 157300 310554
rect 157248 310490 157300 310496
rect 157246 309632 157302 309641
rect 157246 309567 157302 309576
rect 157260 309262 157288 309567
rect 157248 309256 157300 309262
rect 157248 309198 157300 309204
rect 156694 308544 156750 308553
rect 156694 308479 156696 308488
rect 156748 308479 156750 308488
rect 156696 308450 156748 308456
rect 157246 306368 157302 306377
rect 157246 306303 157248 306312
rect 157300 306303 157302 306312
rect 157248 306274 157300 306280
rect 157246 305280 157302 305289
rect 157246 305215 157302 305224
rect 157260 304298 157288 305215
rect 157248 304292 157300 304298
rect 157248 304234 157300 304240
rect 157246 304192 157302 304201
rect 157246 304127 157302 304136
rect 157260 303754 157288 304127
rect 157248 303748 157300 303754
rect 157248 303690 157300 303696
rect 157246 303104 157302 303113
rect 157246 303039 157302 303048
rect 157260 302258 157288 303039
rect 157248 302252 157300 302258
rect 157248 302194 157300 302200
rect 157246 300112 157302 300121
rect 157246 300047 157302 300056
rect 157260 299606 157288 300047
rect 157248 299600 157300 299606
rect 157248 299542 157300 299548
rect 157248 299464 157300 299470
rect 157248 299406 157300 299412
rect 157260 299033 157288 299406
rect 157246 299024 157302 299033
rect 157246 298959 157302 298968
rect 156786 297936 156842 297945
rect 156786 297871 156842 297880
rect 156602 296848 156658 296857
rect 156800 296818 156828 297871
rect 156602 296783 156658 296792
rect 156788 296812 156840 296818
rect 156788 296754 156840 296760
rect 157248 295996 157300 296002
rect 157248 295938 157300 295944
rect 157260 295769 157288 295938
rect 157246 295760 157302 295769
rect 157246 295695 157302 295704
rect 156420 295316 156472 295322
rect 156420 295258 156472 295264
rect 156432 294681 156460 295258
rect 156418 294672 156474 294681
rect 156418 294607 156474 294616
rect 157246 292768 157302 292777
rect 157246 292703 157302 292712
rect 157260 292602 157288 292703
rect 157248 292596 157300 292602
rect 157248 292538 157300 292544
rect 157246 291680 157302 291689
rect 157246 291615 157302 291624
rect 157260 291310 157288 291615
rect 157248 291304 157300 291310
rect 157248 291246 157300 291252
rect 157246 290592 157302 290601
rect 157246 290527 157302 290536
rect 157260 289882 157288 290527
rect 157248 289876 157300 289882
rect 157248 289818 157300 289824
rect 157246 289504 157302 289513
rect 157246 289439 157302 289448
rect 157260 288522 157288 289439
rect 157248 288516 157300 288522
rect 157248 288458 157300 288464
rect 156142 286240 156198 286249
rect 156142 286175 156198 286184
rect 156156 285938 156184 286175
rect 156144 285932 156196 285938
rect 156144 285874 156196 285880
rect 156788 285660 156840 285666
rect 156788 285602 156840 285608
rect 156800 284345 156828 285602
rect 157246 285152 157302 285161
rect 157246 285087 157302 285096
rect 156786 284336 156842 284345
rect 157260 284306 157288 285087
rect 156786 284271 156842 284280
rect 157248 284300 157300 284306
rect 157248 284242 157300 284248
rect 157154 283248 157210 283257
rect 157154 283183 157210 283192
rect 157168 282198 157196 283183
rect 157248 282668 157300 282674
rect 157248 282610 157300 282616
rect 157156 282192 157208 282198
rect 157260 282169 157288 282610
rect 157156 282134 157208 282140
rect 157246 282160 157302 282169
rect 157246 282095 157302 282104
rect 157248 281512 157300 281518
rect 157248 281454 157300 281460
rect 157260 281081 157288 281454
rect 157246 281072 157302 281081
rect 157246 281007 157302 281016
rect 157062 279984 157118 279993
rect 157062 279919 157118 279928
rect 156972 279676 157024 279682
rect 156972 279618 157024 279624
rect 156984 278905 157012 279618
rect 156970 278896 157026 278905
rect 156970 278831 157026 278840
rect 157076 278798 157104 279919
rect 157064 278792 157116 278798
rect 157064 278734 157116 278740
rect 156510 277808 156566 277817
rect 156510 277743 156566 277752
rect 156524 277438 156552 277743
rect 156512 277432 156564 277438
rect 156512 277374 156564 277380
rect 157248 276004 157300 276010
rect 157248 275946 157300 275952
rect 157260 275913 157288 275946
rect 157246 275904 157302 275913
rect 157246 275839 157302 275848
rect 157246 274816 157302 274825
rect 157246 274751 157302 274760
rect 157260 274718 157288 274751
rect 157248 274712 157300 274718
rect 157248 274654 157300 274660
rect 157246 273728 157302 273737
rect 157246 273663 157302 273672
rect 157260 273290 157288 273663
rect 157248 273284 157300 273290
rect 157248 273226 157300 273232
rect 157246 272640 157302 272649
rect 157246 272575 157302 272584
rect 157260 271930 157288 272575
rect 157248 271924 157300 271930
rect 157248 271866 157300 271872
rect 157246 271552 157302 271561
rect 157246 271487 157302 271496
rect 157260 270570 157288 271487
rect 157248 270564 157300 270570
rect 157248 270506 157300 270512
rect 156786 270464 156842 270473
rect 156786 270399 156842 270408
rect 156800 269142 156828 270399
rect 157246 269376 157302 269385
rect 157246 269311 157302 269320
rect 157260 269210 157288 269311
rect 157248 269204 157300 269210
rect 157248 269146 157300 269152
rect 156788 269136 156840 269142
rect 156788 269078 156840 269084
rect 156512 269068 156564 269074
rect 156512 269010 156564 269016
rect 156524 268297 156552 269010
rect 156510 268288 156566 268297
rect 156510 268223 156566 268232
rect 157248 267708 157300 267714
rect 157248 267650 157300 267656
rect 157260 267481 157288 267650
rect 157246 267472 157302 267481
rect 157246 267407 157302 267416
rect 157246 265296 157302 265305
rect 157246 265231 157302 265240
rect 157260 264994 157288 265231
rect 157248 264988 157300 264994
rect 157248 264930 157300 264936
rect 157246 263120 157302 263129
rect 157246 263055 157302 263064
rect 157260 262274 157288 263055
rect 157248 262268 157300 262274
rect 157248 262210 157300 262216
rect 156788 262200 156840 262206
rect 156788 262142 156840 262148
rect 156800 260953 156828 262142
rect 156786 260944 156842 260953
rect 156786 260879 156842 260888
rect 156694 259856 156750 259865
rect 156694 259791 156750 259800
rect 156602 259040 156658 259049
rect 156602 258975 156658 258984
rect 156616 258126 156644 258975
rect 156604 258120 156656 258126
rect 156604 258062 156656 258068
rect 156050 254688 156106 254697
rect 156050 254623 156106 254632
rect 156142 252512 156198 252521
rect 156142 252447 156198 252456
rect 156156 250510 156184 252447
rect 156144 250504 156196 250510
rect 156144 250446 156196 250452
rect 156602 245168 156658 245177
rect 156602 245103 156658 245112
rect 156144 243024 156196 243030
rect 156142 242992 156144 243001
rect 156196 242992 156198 243001
rect 156142 242927 156198 242936
rect 155880 223502 156000 223530
rect 155880 222329 155908 223502
rect 155866 222320 155922 222329
rect 155866 222255 155922 222264
rect 155880 217841 155908 222255
rect 155866 217832 155922 217841
rect 155866 217767 155922 217776
rect 154488 202224 154540 202230
rect 154488 202166 154540 202172
rect 156616 192574 156644 245103
rect 156708 222873 156736 259791
rect 157248 257984 157300 257990
rect 157246 257952 157248 257961
rect 157300 257952 157302 257961
rect 157246 257887 157302 257896
rect 157246 256864 157302 256873
rect 157246 256799 157302 256808
rect 157260 256766 157288 256799
rect 157248 256760 157300 256766
rect 157248 256702 157300 256708
rect 157246 255776 157302 255785
rect 157246 255711 157302 255720
rect 157260 255338 157288 255711
rect 157248 255332 157300 255338
rect 157248 255274 157300 255280
rect 157246 254688 157302 254697
rect 157246 254623 157302 254632
rect 157260 254590 157288 254623
rect 157248 254584 157300 254590
rect 157248 254526 157300 254532
rect 157248 253904 157300 253910
rect 157248 253846 157300 253852
rect 157260 253609 157288 253846
rect 157246 253600 157302 253609
rect 157246 253535 157302 253544
rect 156786 253192 156842 253201
rect 156786 253127 156842 253136
rect 156800 242185 156828 253127
rect 157246 251424 157302 251433
rect 157246 251359 157302 251368
rect 157260 251258 157288 251359
rect 157248 251252 157300 251258
rect 157248 251194 157300 251200
rect 157246 250608 157302 250617
rect 157246 250543 157302 250552
rect 157260 249830 157288 250543
rect 157248 249824 157300 249830
rect 157248 249766 157300 249772
rect 157154 249520 157210 249529
rect 157154 249455 157210 249464
rect 157248 249484 157300 249490
rect 157168 248470 157196 249455
rect 157248 249426 157300 249432
rect 157156 248464 157208 248470
rect 157260 248441 157288 249426
rect 157156 248406 157208 248412
rect 157246 248432 157302 248441
rect 157246 248367 157302 248376
rect 157248 247784 157300 247790
rect 157248 247726 157300 247732
rect 157260 247353 157288 247726
rect 157246 247344 157302 247353
rect 157246 247279 157302 247288
rect 157246 246256 157302 246265
rect 157246 246191 157302 246200
rect 157260 245682 157288 246191
rect 157248 245676 157300 245682
rect 157248 245618 157300 245624
rect 157246 244080 157302 244089
rect 157246 244015 157302 244024
rect 157260 242962 157288 244015
rect 157248 242956 157300 242962
rect 157248 242898 157300 242904
rect 156786 242176 156842 242185
rect 156786 242111 156842 242120
rect 157352 235793 157380 439486
rect 157984 438184 158036 438190
rect 157984 438126 158036 438132
rect 157432 331356 157484 331362
rect 157432 331298 157484 331304
rect 157444 330546 157472 331298
rect 157432 330540 157484 330546
rect 157432 330482 157484 330488
rect 157430 329080 157486 329089
rect 157430 329015 157486 329024
rect 157444 323241 157472 329015
rect 157430 323232 157486 323241
rect 157430 323167 157486 323176
rect 157996 244322 158024 438126
rect 160100 382968 160152 382974
rect 160100 382910 160152 382916
rect 158720 380248 158772 380254
rect 158720 380190 158772 380196
rect 158074 337104 158130 337113
rect 158074 337039 158130 337048
rect 158088 313954 158116 337039
rect 158732 325378 158760 380190
rect 158810 363624 158866 363633
rect 158810 363559 158866 363568
rect 158720 325372 158772 325378
rect 158720 325314 158772 325320
rect 158732 322250 158760 325314
rect 158720 322244 158772 322250
rect 158720 322186 158772 322192
rect 158824 319433 158852 363559
rect 159456 339584 159508 339590
rect 159456 339526 159508 339532
rect 159364 329860 159416 329866
rect 159364 329802 159416 329808
rect 158810 319424 158866 319433
rect 158810 319359 158866 319368
rect 158076 313948 158128 313954
rect 158076 313890 158128 313896
rect 158076 309324 158128 309330
rect 158076 309266 158128 309272
rect 158088 291174 158116 309266
rect 159376 297401 159404 329802
rect 159468 308417 159496 339526
rect 159548 308508 159600 308514
rect 159548 308450 159600 308456
rect 159454 308408 159510 308417
rect 159454 308343 159510 308352
rect 159362 297392 159418 297401
rect 159362 297327 159418 297336
rect 158076 291168 158128 291174
rect 158076 291110 158128 291116
rect 159456 286340 159508 286346
rect 159456 286282 159508 286288
rect 158076 285932 158128 285938
rect 158076 285874 158128 285880
rect 158088 247722 158116 285874
rect 159362 284336 159418 284345
rect 159362 284271 159418 284280
rect 158168 268388 158220 268394
rect 158168 268330 158220 268336
rect 158076 247716 158128 247722
rect 158076 247658 158128 247664
rect 157984 244316 158036 244322
rect 157984 244258 158036 244264
rect 157338 235784 157394 235793
rect 157338 235719 157394 235728
rect 156694 222864 156750 222873
rect 156694 222799 156750 222808
rect 157996 202774 158024 244258
rect 158076 243024 158128 243030
rect 158076 242966 158128 242972
rect 158088 213926 158116 242966
rect 158180 231577 158208 268330
rect 159376 234598 159404 284271
rect 159468 243545 159496 286282
rect 159560 284986 159588 308450
rect 159548 284980 159600 284986
rect 159548 284922 159600 284928
rect 159548 264240 159600 264246
rect 159548 264182 159600 264188
rect 159454 243536 159510 243545
rect 159454 243471 159510 243480
rect 159364 234592 159416 234598
rect 159364 234534 159416 234540
rect 159456 233300 159508 233306
rect 159456 233242 159508 233248
rect 158166 231568 158222 231577
rect 158166 231503 158222 231512
rect 159468 218006 159496 233242
rect 159560 233170 159588 264182
rect 159640 256012 159692 256018
rect 159640 255954 159692 255960
rect 159548 233164 159600 233170
rect 159548 233106 159600 233112
rect 159652 226137 159680 255954
rect 159730 243128 159786 243137
rect 159730 243063 159786 243072
rect 159638 226128 159694 226137
rect 159638 226063 159694 226072
rect 159744 219201 159772 243063
rect 160112 237153 160140 382910
rect 160190 358048 160246 358057
rect 160190 357983 160246 357992
rect 160204 306338 160232 357983
rect 160836 332716 160888 332722
rect 160836 332658 160888 332664
rect 160848 315353 160876 332658
rect 160928 318844 160980 318850
rect 160928 318786 160980 318792
rect 160834 315344 160890 315353
rect 160940 315314 160968 318786
rect 160834 315279 160890 315288
rect 160928 315308 160980 315314
rect 160928 315250 160980 315256
rect 160744 314696 160796 314702
rect 160744 314638 160796 314644
rect 160192 306332 160244 306338
rect 160192 306274 160244 306280
rect 160204 305726 160232 306274
rect 160192 305720 160244 305726
rect 160192 305662 160244 305668
rect 160756 294545 160784 314638
rect 160926 303784 160982 303793
rect 160926 303719 160982 303728
rect 160742 294536 160798 294545
rect 160742 294471 160798 294480
rect 160744 291168 160796 291174
rect 160744 291110 160796 291116
rect 160098 237144 160154 237153
rect 160098 237079 160154 237088
rect 159730 219192 159786 219201
rect 159730 219127 159786 219136
rect 159456 218000 159508 218006
rect 159456 217942 159508 217948
rect 158076 213920 158128 213926
rect 158076 213862 158128 213868
rect 157984 202768 158036 202774
rect 157984 202710 158036 202716
rect 156604 192568 156656 192574
rect 156604 192510 156656 192516
rect 151726 191040 151782 191049
rect 151726 190975 151782 190984
rect 160756 187105 160784 291110
rect 160834 283520 160890 283529
rect 160834 283455 160890 283464
rect 160848 234433 160876 283455
rect 160940 279682 160968 303719
rect 161492 296002 161520 452678
rect 173808 451240 173860 451246
rect 173808 451182 173860 451188
rect 167000 450016 167052 450022
rect 167000 449958 167052 449964
rect 172518 449984 172574 449993
rect 163504 403640 163556 403646
rect 163504 403582 163556 403588
rect 163516 403034 163544 403582
rect 163504 403028 163556 403034
rect 163504 402970 163556 402976
rect 161572 370524 161624 370530
rect 161572 370466 161624 370472
rect 161584 317422 161612 370466
rect 162124 365832 162176 365838
rect 162124 365774 162176 365780
rect 161572 317416 161624 317422
rect 161572 317358 161624 317364
rect 161480 295996 161532 296002
rect 161480 295938 161532 295944
rect 160928 279676 160980 279682
rect 160928 279618 160980 279624
rect 160926 275360 160982 275369
rect 160926 275295 160982 275304
rect 160940 237386 160968 275295
rect 162136 269113 162164 365774
rect 162216 327820 162268 327826
rect 162216 327762 162268 327768
rect 162122 269104 162178 269113
rect 162122 269039 162178 269048
rect 162228 260166 162256 327762
rect 162768 317416 162820 317422
rect 162768 317358 162820 317364
rect 162780 316810 162808 317358
rect 162768 316804 162820 316810
rect 162768 316746 162820 316752
rect 162400 299532 162452 299538
rect 162400 299474 162452 299480
rect 162308 285728 162360 285734
rect 162308 285670 162360 285676
rect 162216 260160 162268 260166
rect 162216 260102 162268 260108
rect 162124 258120 162176 258126
rect 162124 258062 162176 258068
rect 160928 237380 160980 237386
rect 160928 237322 160980 237328
rect 160834 234424 160890 234433
rect 160834 234359 160890 234368
rect 162136 200705 162164 258062
rect 162320 234297 162348 285670
rect 162412 282674 162440 299474
rect 162766 296032 162822 296041
rect 162766 295967 162768 295976
rect 162820 295967 162822 295976
rect 162768 295938 162820 295944
rect 162400 282668 162452 282674
rect 162400 282610 162452 282616
rect 162492 271176 162544 271182
rect 162492 271118 162544 271124
rect 162400 265668 162452 265674
rect 162400 265610 162452 265616
rect 162306 234288 162362 234297
rect 162306 234223 162362 234232
rect 162412 228857 162440 265610
rect 162504 257990 162532 271118
rect 162492 257984 162544 257990
rect 162492 257926 162544 257932
rect 162398 228848 162454 228857
rect 162398 228783 162454 228792
rect 163516 227361 163544 402970
rect 165620 389224 165672 389230
rect 165620 389166 165672 389172
rect 163596 376032 163648 376038
rect 163596 375974 163648 375980
rect 163608 298217 163636 375974
rect 164332 374672 164384 374678
rect 164332 374614 164384 374620
rect 164238 355464 164294 355473
rect 164238 355399 164294 355408
rect 163778 332888 163834 332897
rect 163778 332823 163834 332832
rect 163688 321632 163740 321638
rect 163688 321574 163740 321580
rect 163700 305658 163728 321574
rect 163792 316742 163820 332823
rect 163780 316736 163832 316742
rect 163780 316678 163832 316684
rect 163688 305652 163740 305658
rect 163688 305594 163740 305600
rect 163594 298208 163650 298217
rect 163594 298143 163650 298152
rect 163608 231713 163636 298143
rect 163688 288448 163740 288454
rect 163688 288390 163740 288396
rect 163700 269074 163728 288390
rect 164252 286385 164280 355399
rect 164344 315382 164372 374614
rect 164884 338224 164936 338230
rect 164884 338166 164936 338172
rect 164896 319462 164924 338166
rect 164976 327752 165028 327758
rect 164976 327694 165028 327700
rect 164884 319456 164936 319462
rect 164884 319398 164936 319404
rect 164988 318102 165016 327694
rect 164976 318096 165028 318102
rect 164976 318038 165028 318044
rect 164332 315376 164384 315382
rect 164332 315318 164384 315324
rect 164344 314702 164372 315318
rect 164332 314696 164384 314702
rect 164332 314638 164384 314644
rect 165068 314696 165120 314702
rect 165068 314638 165120 314644
rect 164974 289096 165030 289105
rect 164974 289031 165030 289040
rect 164884 287088 164936 287094
rect 164884 287030 164936 287036
rect 164238 286376 164294 286385
rect 164238 286311 164294 286320
rect 164252 285734 164280 286311
rect 164240 285728 164292 285734
rect 164240 285670 164292 285676
rect 164238 269104 164294 269113
rect 163688 269068 163740 269074
rect 164238 269039 164294 269048
rect 163688 269010 163740 269016
rect 163688 263628 163740 263634
rect 163688 263570 163740 263576
rect 163700 249490 163728 263570
rect 163688 249484 163740 249490
rect 163688 249426 163740 249432
rect 163594 231704 163650 231713
rect 163594 231639 163650 231648
rect 163502 227352 163558 227361
rect 163502 227287 163558 227296
rect 164252 211818 164280 269039
rect 164896 223582 164924 287030
rect 164988 242049 165016 289031
rect 165080 269074 165108 314638
rect 165068 269068 165120 269074
rect 165068 269010 165120 269016
rect 165632 262206 165660 389166
rect 165712 374740 165764 374746
rect 165712 374682 165764 374688
rect 165724 299470 165752 374682
rect 165712 299464 165764 299470
rect 165712 299406 165764 299412
rect 166080 299464 166132 299470
rect 166080 299406 166132 299412
rect 166092 298790 166120 299406
rect 166080 298784 166132 298790
rect 166080 298726 166132 298732
rect 166448 273284 166500 273290
rect 166448 273226 166500 273232
rect 166264 269204 166316 269210
rect 166264 269146 166316 269152
rect 165620 262200 165672 262206
rect 165620 262142 165672 262148
rect 165528 255332 165580 255338
rect 165528 255274 165580 255280
rect 165540 251870 165568 255274
rect 165528 251864 165580 251870
rect 165528 251806 165580 251812
rect 165528 247784 165580 247790
rect 165528 247726 165580 247732
rect 165540 247081 165568 247726
rect 165526 247072 165582 247081
rect 165526 247007 165582 247016
rect 164974 242040 165030 242049
rect 164974 241975 165030 241984
rect 164884 223576 164936 223582
rect 164884 223518 164936 223524
rect 166276 211857 166304 269146
rect 166356 247104 166408 247110
rect 166356 247046 166408 247052
rect 166262 211848 166318 211857
rect 164240 211812 164292 211818
rect 166262 211783 166318 211792
rect 164240 211754 164292 211760
rect 162122 200696 162178 200705
rect 162122 200631 162178 200640
rect 166264 200116 166316 200122
rect 166368 200114 166396 247046
rect 166460 242214 166488 273226
rect 166540 245744 166592 245750
rect 166540 245686 166592 245692
rect 166448 242208 166500 242214
rect 166448 242150 166500 242156
rect 166552 226001 166580 245686
rect 167012 231849 167040 449958
rect 173820 449954 173848 451182
rect 172518 449919 172520 449928
rect 172572 449919 172574 449928
rect 173808 449948 173860 449954
rect 172520 449890 172572 449896
rect 173808 449890 173860 449896
rect 168470 447400 168526 447409
rect 168470 447335 168526 447344
rect 167644 343732 167696 343738
rect 167644 343674 167696 343680
rect 167656 253230 167684 343674
rect 167736 342304 167788 342310
rect 167736 342246 167788 342252
rect 167748 319530 167776 342246
rect 167826 325272 167882 325281
rect 167826 325207 167882 325216
rect 167736 319524 167788 319530
rect 167736 319466 167788 319472
rect 167840 309126 167868 325207
rect 167828 309120 167880 309126
rect 167828 309062 167880 309068
rect 168288 309120 168340 309126
rect 168288 309062 168340 309068
rect 167734 278080 167790 278089
rect 167734 278015 167790 278024
rect 167644 253224 167696 253230
rect 167644 253166 167696 253172
rect 167748 247110 167776 278015
rect 168300 274650 168328 309062
rect 168288 274644 168340 274650
rect 168288 274586 168340 274592
rect 168380 251252 168432 251258
rect 168380 251194 168432 251200
rect 167736 247104 167788 247110
rect 167736 247046 167788 247052
rect 167642 237416 167698 237425
rect 167642 237351 167698 237360
rect 166998 231840 167054 231849
rect 166998 231775 167054 231784
rect 167656 230217 167684 237351
rect 167642 230208 167698 230217
rect 167642 230143 167698 230152
rect 167656 226137 167684 230143
rect 167642 226128 167698 226137
rect 167642 226063 167698 226072
rect 166538 225992 166594 226001
rect 166538 225927 166594 225936
rect 167826 200968 167882 200977
rect 167826 200903 167882 200912
rect 166316 200086 166396 200114
rect 166264 200058 166316 200064
rect 160742 187096 160798 187105
rect 160742 187031 160798 187040
rect 115848 186992 115900 186998
rect 115848 186934 115900 186940
rect 119988 186380 120040 186386
rect 119988 186322 120040 186328
rect 164884 186380 164936 186386
rect 164884 186322 164936 186328
rect 113732 182232 113784 182238
rect 113732 182174 113784 182180
rect 107474 180976 107530 180985
rect 107474 180911 107530 180920
rect 107488 177585 107516 180911
rect 112258 179616 112314 179625
rect 112258 179551 112314 179560
rect 106186 177576 106242 177585
rect 106186 177511 106242 177520
rect 107474 177576 107530 177585
rect 107474 177511 107530 177520
rect 112272 177177 112300 179551
rect 113744 177585 113772 182174
rect 116950 180840 117006 180849
rect 116950 180775 117006 180784
rect 115848 178084 115900 178090
rect 115848 178026 115900 178032
rect 113730 177576 113786 177585
rect 113730 177511 113786 177520
rect 112258 177168 112314 177177
rect 112258 177103 112314 177112
rect 105452 176928 105504 176934
rect 105452 176870 105504 176876
rect 115860 176769 115888 178026
rect 116964 177585 116992 180775
rect 118516 179512 118568 179518
rect 118516 179454 118568 179460
rect 116950 177576 117006 177585
rect 116950 177511 117006 177520
rect 118528 177177 118556 179454
rect 120000 177585 120028 186322
rect 121368 184952 121420 184958
rect 121368 184894 121420 184900
rect 121380 177585 121408 184894
rect 148968 183660 149020 183666
rect 148968 183602 149020 183608
rect 129648 183592 129700 183598
rect 129648 183534 129700 183540
rect 126060 180872 126112 180878
rect 126060 180814 126112 180820
rect 124496 178152 124548 178158
rect 124496 178094 124548 178100
rect 119986 177576 120042 177585
rect 119986 177511 120042 177520
rect 121366 177576 121422 177585
rect 121366 177511 121422 177520
rect 118514 177168 118570 177177
rect 118514 177103 118570 177112
rect 124508 176769 124536 178094
rect 126072 177585 126100 180814
rect 127624 177744 127676 177750
rect 127624 177686 127676 177692
rect 126058 177576 126114 177585
rect 126058 177511 126114 177520
rect 127636 176769 127664 177686
rect 129660 177585 129688 183534
rect 132500 180940 132552 180946
rect 132500 180882 132552 180888
rect 132408 179444 132460 179450
rect 132408 179386 132460 179392
rect 129646 177576 129702 177585
rect 129646 177511 129702 177520
rect 132420 176769 132448 179386
rect 132512 177750 132540 180882
rect 132500 177744 132552 177750
rect 132500 177686 132552 177692
rect 148980 177585 149008 183602
rect 148966 177576 149022 177585
rect 148966 177511 149022 177520
rect 134432 176792 134484 176798
rect 99470 176760 99526 176769
rect 99470 176695 99526 176704
rect 102046 176760 102102 176769
rect 102046 176695 102102 176704
rect 103334 176760 103390 176769
rect 103334 176695 103390 176704
rect 115846 176760 115902 176769
rect 115846 176695 115902 176704
rect 124494 176760 124550 176769
rect 124494 176695 124550 176704
rect 127622 176760 127678 176769
rect 127622 176695 127678 176704
rect 132406 176760 132462 176769
rect 132406 176695 132462 176704
rect 134430 176760 134432 176769
rect 143448 176792 143500 176798
rect 134484 176760 134486 176769
rect 134430 176695 134486 176704
rect 136086 176760 136142 176769
rect 158996 176792 159048 176798
rect 143448 176734 143500 176740
rect 158994 176760 158996 176769
rect 159048 176760 159050 176769
rect 136086 176695 136088 176704
rect 136140 176695 136142 176704
rect 136088 176666 136140 176672
rect 130752 176044 130804 176050
rect 130752 175986 130804 175992
rect 123116 175976 123168 175982
rect 123116 175918 123168 175924
rect 123128 175001 123156 175918
rect 130764 175817 130792 175986
rect 130750 175808 130806 175817
rect 130750 175743 130806 175752
rect 143460 175234 143488 176734
rect 158994 176695 159050 176704
rect 143448 175228 143500 175234
rect 143448 175170 143500 175176
rect 123114 174992 123170 175001
rect 123114 174927 123170 174936
rect 164896 167006 164924 186322
rect 164976 178152 165028 178158
rect 164976 178094 165028 178100
rect 164988 169726 165016 178094
rect 165528 176044 165580 176050
rect 165528 175986 165580 175992
rect 165540 173874 165568 175986
rect 165528 173868 165580 173874
rect 165528 173810 165580 173816
rect 164976 169720 165028 169726
rect 166276 169697 166304 200058
rect 167644 183660 167696 183666
rect 167644 183602 167696 183608
rect 166448 180872 166500 180878
rect 166448 180814 166500 180820
rect 166354 176896 166410 176905
rect 166354 176831 166410 176840
rect 164976 169662 165028 169668
rect 166262 169688 166318 169697
rect 166262 169623 166318 169632
rect 164884 167000 164936 167006
rect 164884 166942 164936 166948
rect 166368 155922 166396 176831
rect 166460 171086 166488 180814
rect 166448 171080 166500 171086
rect 166448 171022 166500 171028
rect 166356 155916 166408 155922
rect 166356 155858 166408 155864
rect 167656 150414 167684 183602
rect 167840 181490 167868 200903
rect 167920 184952 167972 184958
rect 167920 184894 167972 184900
rect 167828 181484 167880 181490
rect 167828 181426 167880 181432
rect 167734 180976 167790 180985
rect 167734 180911 167790 180920
rect 167748 161430 167776 180911
rect 167932 168366 167960 184894
rect 167920 168360 167972 168366
rect 167920 168302 167972 168308
rect 167736 161424 167788 161430
rect 167736 161366 167788 161372
rect 167644 150408 167696 150414
rect 167644 150350 167696 150356
rect 167736 137284 167788 137290
rect 167736 137226 167788 137232
rect 167644 135312 167696 135318
rect 167644 135254 167696 135260
rect 67362 129296 67418 129305
rect 67362 129231 67418 129240
rect 66166 126304 66222 126313
rect 66166 126239 66222 126248
rect 66074 123584 66130 123593
rect 66074 123519 66130 123528
rect 65982 120864 66038 120873
rect 65982 120799 66038 120808
rect 65996 90370 66024 120799
rect 66088 93158 66116 123519
rect 66076 93152 66128 93158
rect 66076 93094 66128 93100
rect 65984 90364 66036 90370
rect 65984 90306 66036 90312
rect 66180 86290 66208 126239
rect 67270 102368 67326 102377
rect 67270 102303 67326 102312
rect 67284 95169 67312 102303
rect 67270 95160 67326 95169
rect 67270 95095 67326 95104
rect 67376 93226 67404 129231
rect 67730 128072 67786 128081
rect 67730 128007 67786 128016
rect 67454 125216 67510 125225
rect 67454 125151 67510 125160
rect 67364 93220 67416 93226
rect 67364 93162 67416 93168
rect 66168 86284 66220 86290
rect 66168 86226 66220 86232
rect 67468 81433 67496 125151
rect 67546 122632 67602 122641
rect 67546 122567 67602 122576
rect 67454 81424 67510 81433
rect 67454 81359 67510 81368
rect 64418 68368 64474 68377
rect 64418 68303 64474 68312
rect 67560 66201 67588 122567
rect 67638 100736 67694 100745
rect 67638 100671 67694 100680
rect 67546 66192 67602 66201
rect 67546 66127 67602 66136
rect 67652 63481 67680 100671
rect 67744 94518 67772 128007
rect 164884 123480 164936 123486
rect 164884 123422 164936 123428
rect 124034 94752 124090 94761
rect 124034 94687 124090 94696
rect 67732 94512 67784 94518
rect 67732 94454 67784 94460
rect 100024 94512 100076 94518
rect 100024 94454 100076 94460
rect 88984 93220 89036 93226
rect 88984 93162 89036 93168
rect 86866 92440 86922 92449
rect 86866 92375 86922 92384
rect 75826 91216 75882 91225
rect 86774 91216 86830 91225
rect 75882 91174 75960 91202
rect 75826 91151 75882 91160
rect 75932 86970 75960 91174
rect 86880 91186 86908 92375
rect 88154 91216 88210 91225
rect 86774 91151 86830 91160
rect 86868 91180 86920 91186
rect 75920 86964 75972 86970
rect 75920 86906 75972 86912
rect 70214 76664 70270 76673
rect 70214 76599 70270 76608
rect 67638 63472 67694 63481
rect 67638 63407 67694 63416
rect 66166 60072 66222 60081
rect 66166 60007 66222 60016
rect 64786 51776 64842 51785
rect 64786 51711 64842 51720
rect 63408 14476 63460 14482
rect 63408 14418 63460 14424
rect 62028 3596 62080 3602
rect 62028 3538 62080 3544
rect 63224 3528 63276 3534
rect 61948 3454 62068 3482
rect 63224 3470 63276 3476
rect 62040 480 62068 3454
rect 63236 480 63264 3470
rect 64800 3466 64828 51711
rect 66180 3466 66208 60007
rect 70228 16574 70256 76599
rect 86788 73846 86816 91151
rect 88154 91151 88210 91160
rect 86868 91122 86920 91128
rect 86776 73840 86828 73846
rect 86776 73782 86828 73788
rect 79966 71088 80022 71097
rect 79966 71023 80022 71032
rect 71044 66904 71096 66910
rect 71044 66846 71096 66852
rect 70228 16546 70348 16574
rect 68928 15972 68980 15978
rect 68928 15914 68980 15920
rect 66720 8968 66772 8974
rect 66720 8910 66772 8916
rect 64328 3460 64380 3466
rect 64328 3402 64380 3408
rect 64788 3460 64840 3466
rect 64788 3402 64840 3408
rect 65524 3460 65576 3466
rect 65524 3402 65576 3408
rect 66168 3460 66220 3466
rect 66168 3402 66220 3408
rect 64340 480 64368 3402
rect 65536 480 65564 3402
rect 66732 480 66760 8910
rect 68940 3466 68968 15914
rect 69112 4888 69164 4894
rect 69112 4830 69164 4836
rect 67916 3460 67968 3466
rect 67916 3402 67968 3408
rect 68928 3460 68980 3466
rect 68928 3402 68980 3408
rect 67928 480 67956 3402
rect 69124 480 69152 4830
rect 70320 480 70348 16546
rect 71056 7682 71084 66846
rect 78586 61432 78642 61441
rect 78586 61367 78642 61376
rect 73066 58576 73122 58585
rect 73066 58511 73122 58520
rect 71688 47660 71740 47666
rect 71688 47602 71740 47608
rect 71044 7676 71096 7682
rect 71044 7618 71096 7624
rect 71700 6914 71728 47602
rect 71516 6886 71728 6914
rect 71516 480 71544 6886
rect 73080 3466 73108 58511
rect 77208 57248 77260 57254
rect 77208 57190 77260 57196
rect 75828 43444 75880 43450
rect 75828 43386 75880 43392
rect 74448 39432 74500 39438
rect 74448 39374 74500 39380
rect 74460 3466 74488 39374
rect 75840 3466 75868 43386
rect 77220 3466 77248 57190
rect 72608 3460 72660 3466
rect 72608 3402 72660 3408
rect 73068 3460 73120 3466
rect 73068 3402 73120 3408
rect 73804 3460 73856 3466
rect 73804 3402 73856 3408
rect 74448 3460 74500 3466
rect 74448 3402 74500 3408
rect 75000 3460 75052 3466
rect 75000 3402 75052 3408
rect 75828 3460 75880 3466
rect 75828 3402 75880 3408
rect 76196 3460 76248 3466
rect 76196 3402 76248 3408
rect 77208 3460 77260 3466
rect 77208 3402 77260 3408
rect 72620 480 72648 3402
rect 73816 480 73844 3402
rect 75012 480 75040 3402
rect 76208 480 76236 3402
rect 77392 3392 77444 3398
rect 77392 3334 77444 3340
rect 77404 480 77432 3334
rect 78600 480 78628 61367
rect 79324 36644 79376 36650
rect 79324 36586 79376 36592
rect 79336 15910 79364 36586
rect 79324 15904 79376 15910
rect 79324 15846 79376 15852
rect 79980 6914 80008 71023
rect 88168 64870 88196 91151
rect 88996 78674 89024 93162
rect 89074 92440 89130 92449
rect 89074 92375 89130 92384
rect 89088 91118 89116 92375
rect 98734 91488 98790 91497
rect 98734 91423 98790 91432
rect 95054 91352 95110 91361
rect 95054 91287 95110 91296
rect 91006 91216 91062 91225
rect 91006 91151 91062 91160
rect 91926 91216 91982 91225
rect 91926 91151 91982 91160
rect 93214 91216 93270 91225
rect 93214 91151 93270 91160
rect 89076 91112 89128 91118
rect 89076 91054 89128 91060
rect 88984 78668 89036 78674
rect 88984 78610 89036 78616
rect 91020 77246 91048 91151
rect 91940 88233 91968 91151
rect 91926 88224 91982 88233
rect 91926 88159 91982 88168
rect 93228 85513 93256 91151
rect 93214 85504 93270 85513
rect 93214 85439 93270 85448
rect 95068 84182 95096 91287
rect 95146 91216 95202 91225
rect 95146 91151 95202 91160
rect 96526 91216 96582 91225
rect 96526 91151 96582 91160
rect 97906 91216 97962 91225
rect 97906 91151 97962 91160
rect 95056 84176 95108 84182
rect 95056 84118 95108 84124
rect 95160 81394 95188 91151
rect 96540 82822 96568 91151
rect 97920 84114 97948 91151
rect 98748 89010 98776 91423
rect 99194 91216 99250 91225
rect 99194 91151 99250 91160
rect 98736 89004 98788 89010
rect 98736 88946 98788 88952
rect 97908 84108 97960 84114
rect 97908 84050 97960 84056
rect 96528 82816 96580 82822
rect 96528 82758 96580 82764
rect 95148 81388 95200 81394
rect 95148 81330 95200 81336
rect 99208 80073 99236 91151
rect 99286 80744 99342 80753
rect 99286 80679 99342 80688
rect 99194 80064 99250 80073
rect 99194 79999 99250 80008
rect 91008 77240 91060 77246
rect 91008 77182 91060 77188
rect 97908 75200 97960 75206
rect 88246 75168 88302 75177
rect 97908 75142 97960 75148
rect 88246 75103 88302 75112
rect 88156 64864 88208 64870
rect 88156 64806 88208 64812
rect 86868 50380 86920 50386
rect 86868 50322 86920 50328
rect 84108 43512 84160 43518
rect 84108 43454 84160 43460
rect 81348 24132 81400 24138
rect 81348 24074 81400 24080
rect 79704 6886 80008 6914
rect 79704 480 79732 6886
rect 81360 3466 81388 24074
rect 82082 3632 82138 3641
rect 82082 3567 82138 3576
rect 80888 3460 80940 3466
rect 80888 3402 80940 3408
rect 81348 3460 81400 3466
rect 81348 3402 81400 3408
rect 80900 480 80928 3402
rect 82096 480 82124 3567
rect 84120 3466 84148 43454
rect 86774 17232 86830 17241
rect 86774 17167 86830 17176
rect 86788 3466 86816 17167
rect 83280 3460 83332 3466
rect 83280 3402 83332 3408
rect 84108 3460 84160 3466
rect 84108 3402 84160 3408
rect 85672 3460 85724 3466
rect 85672 3402 85724 3408
rect 86776 3460 86828 3466
rect 86776 3402 86828 3408
rect 83292 480 83320 3402
rect 84476 2168 84528 2174
rect 84476 2110 84528 2116
rect 84488 480 84516 2110
rect 85684 480 85712 3402
rect 86880 480 86908 50322
rect 88260 6914 88288 75103
rect 95146 72584 95202 72593
rect 95146 72519 95202 72528
rect 91008 55888 91060 55894
rect 91008 55830 91060 55836
rect 88984 15904 89036 15910
rect 88984 15846 89036 15852
rect 87984 6886 88288 6914
rect 87984 480 88012 6886
rect 88996 3398 89024 15846
rect 89168 6248 89220 6254
rect 89168 6190 89220 6196
rect 88984 3392 89036 3398
rect 88984 3334 89036 3340
rect 89180 480 89208 6190
rect 91020 3058 91048 55830
rect 95056 54528 95108 54534
rect 95056 54470 95108 54476
rect 92388 13184 92440 13190
rect 92388 13126 92440 13132
rect 92400 3466 92428 13126
rect 92756 7676 92808 7682
rect 92756 7618 92808 7624
rect 91560 3460 91612 3466
rect 91560 3402 91612 3408
rect 92388 3460 92440 3466
rect 92388 3402 92440 3408
rect 90364 3052 90416 3058
rect 90364 2994 90416 3000
rect 91008 3052 91060 3058
rect 91008 2994 91060 3000
rect 90376 480 90404 2994
rect 91572 480 91600 3402
rect 92768 480 92796 7618
rect 95068 3058 95096 54470
rect 93952 3052 94004 3058
rect 93952 2994 94004 3000
rect 95056 3052 95108 3058
rect 95056 2994 95108 3000
rect 93964 480 93992 2994
rect 95160 480 95188 72519
rect 96528 25560 96580 25566
rect 96528 25502 96580 25508
rect 96540 6914 96568 25502
rect 96264 6886 96568 6914
rect 96264 480 96292 6886
rect 97920 3534 97948 75142
rect 99300 3534 99328 80679
rect 100036 73166 100064 94454
rect 124048 93906 124076 94687
rect 162860 94444 162912 94450
rect 162860 94386 162912 94392
rect 124036 93900 124088 93906
rect 124036 93842 124088 93848
rect 119710 93528 119766 93537
rect 119710 93463 119766 93472
rect 121734 93528 121790 93537
rect 121734 93463 121790 93472
rect 110142 93256 110198 93265
rect 119724 93226 119752 93463
rect 110142 93191 110198 93200
rect 119712 93220 119764 93226
rect 106188 93152 106240 93158
rect 106188 93094 106240 93100
rect 105542 91760 105598 91769
rect 105542 91695 105598 91704
rect 101862 91488 101918 91497
rect 101862 91423 101918 91432
rect 100666 91216 100722 91225
rect 100666 91151 100722 91160
rect 100680 74361 100708 91151
rect 101876 86873 101904 91423
rect 102046 91352 102102 91361
rect 102046 91287 102102 91296
rect 101954 91216 102010 91225
rect 101954 91151 102010 91160
rect 101862 86864 101918 86873
rect 101862 86799 101918 86808
rect 100666 74352 100722 74361
rect 100666 74287 100722 74296
rect 100024 73160 100076 73166
rect 100024 73102 100076 73108
rect 100666 58712 100722 58721
rect 100666 58647 100722 58656
rect 100680 3534 100708 58647
rect 101968 57934 101996 91151
rect 101956 57928 102008 57934
rect 101956 57870 102008 57876
rect 102060 55214 102088 91287
rect 102598 91216 102654 91225
rect 102598 91151 102654 91160
rect 103426 91216 103482 91225
rect 103426 91151 103482 91160
rect 104254 91216 104310 91225
rect 104254 91151 104310 91160
rect 104806 91216 104862 91225
rect 104806 91151 104862 91160
rect 102612 88330 102640 91151
rect 102600 88324 102652 88330
rect 102600 88266 102652 88272
rect 103440 64802 103468 91151
rect 104268 85241 104296 91151
rect 104254 85232 104310 85241
rect 104254 85167 104310 85176
rect 103428 64796 103480 64802
rect 103428 64738 103480 64744
rect 104820 63442 104848 91151
rect 105556 81297 105584 91695
rect 106200 85377 106228 93094
rect 109958 92440 110014 92449
rect 109958 92375 110014 92384
rect 107474 91760 107530 91769
rect 107474 91695 107530 91704
rect 106924 91180 106976 91186
rect 106924 91122 106976 91128
rect 106186 85368 106242 85377
rect 106186 85303 106242 85312
rect 105542 81288 105598 81297
rect 105542 81223 105598 81232
rect 105544 73840 105596 73846
rect 105544 73782 105596 73788
rect 104808 63436 104860 63442
rect 104808 63378 104860 63384
rect 105556 60722 105584 73782
rect 106936 66162 106964 91122
rect 107488 89622 107516 91695
rect 108854 91352 108910 91361
rect 108854 91287 108910 91296
rect 107476 89616 107528 89622
rect 107476 89558 107528 89564
rect 107016 86284 107068 86290
rect 107016 86226 107068 86232
rect 107028 74497 107056 86226
rect 107014 74488 107070 74497
rect 107014 74423 107070 74432
rect 108868 69018 108896 91287
rect 108946 91216 109002 91225
rect 108946 91151 109002 91160
rect 108856 69012 108908 69018
rect 108856 68954 108908 68960
rect 106924 66156 106976 66162
rect 106924 66098 106976 66104
rect 105544 60716 105596 60722
rect 105544 60658 105596 60664
rect 108960 59362 108988 91151
rect 109972 91050 110000 92375
rect 109960 91044 110012 91050
rect 109960 90986 110012 90992
rect 110156 89593 110184 93191
rect 119712 93162 119764 93168
rect 121748 93158 121776 93463
rect 121736 93152 121788 93158
rect 121736 93094 121788 93100
rect 158718 93120 158774 93129
rect 158718 93055 158774 93064
rect 136088 92472 136140 92478
rect 111614 92440 111670 92449
rect 111614 92375 111670 92384
rect 114466 92440 114522 92449
rect 114466 92375 114522 92384
rect 136086 92440 136088 92449
rect 136140 92440 136142 92449
rect 136086 92375 136142 92384
rect 151358 92440 151414 92449
rect 151358 92375 151360 92384
rect 110326 91216 110382 91225
rect 110326 91151 110382 91160
rect 111154 91216 111210 91225
rect 111154 91151 111210 91160
rect 110142 89584 110198 89593
rect 110142 89519 110198 89528
rect 110340 67590 110368 91151
rect 111064 90364 111116 90370
rect 111064 90306 111116 90312
rect 111076 82793 111104 90306
rect 111168 88097 111196 91151
rect 111628 90982 111656 92375
rect 112074 91216 112130 91225
rect 112074 91151 112130 91160
rect 112994 91216 113050 91225
rect 112994 91151 113050 91160
rect 113454 91216 113510 91225
rect 113454 91151 113510 91160
rect 114282 91216 114338 91225
rect 114480 91186 114508 92375
rect 151412 92375 151414 92384
rect 151360 92346 151412 92352
rect 126886 92304 126942 92313
rect 126886 92239 126942 92248
rect 126610 91896 126666 91905
rect 126610 91831 126666 91840
rect 117228 91792 117280 91798
rect 114926 91760 114982 91769
rect 117228 91734 117280 91740
rect 114926 91695 114982 91704
rect 114282 91151 114338 91160
rect 114468 91180 114520 91186
rect 111616 90976 111668 90982
rect 111616 90918 111668 90924
rect 111154 88088 111210 88097
rect 111154 88023 111210 88032
rect 112088 86737 112116 91151
rect 112074 86728 112130 86737
rect 112074 86663 112130 86672
rect 111062 82784 111118 82793
rect 111062 82719 111118 82728
rect 110328 67584 110380 67590
rect 110328 67526 110380 67532
rect 113008 66230 113036 91151
rect 113468 86902 113496 91151
rect 113456 86896 113508 86902
rect 113456 86838 113508 86844
rect 114296 82754 114324 91151
rect 114468 91122 114520 91128
rect 114940 89729 114968 91695
rect 117240 91633 117268 91734
rect 117226 91624 117282 91633
rect 117226 91559 117282 91568
rect 115754 91352 115810 91361
rect 115754 91287 115810 91296
rect 118514 91352 118570 91361
rect 118514 91287 118570 91296
rect 122838 91352 122894 91361
rect 122838 91287 122894 91296
rect 125414 91352 125470 91361
rect 125414 91287 125470 91296
rect 114926 89720 114982 89729
rect 114926 89655 114982 89664
rect 115768 84153 115796 91287
rect 115846 91216 115902 91225
rect 115846 91151 115902 91160
rect 117226 91216 117282 91225
rect 117226 91151 117282 91160
rect 115754 84144 115810 84153
rect 115754 84079 115810 84088
rect 114284 82748 114336 82754
rect 114284 82690 114336 82696
rect 113088 71052 113140 71058
rect 113088 70994 113140 71000
rect 112996 66224 113048 66230
rect 112996 66166 113048 66172
rect 108948 59356 109000 59362
rect 108948 59298 109000 59304
rect 103426 57216 103482 57225
rect 103426 57151 103482 57160
rect 102048 55208 102100 55214
rect 102048 55150 102100 55156
rect 102048 53100 102100 53106
rect 102048 53042 102100 53048
rect 102060 3534 102088 53042
rect 103440 6914 103468 57151
rect 111706 55856 111762 55865
rect 111706 55791 111762 55800
rect 106922 54496 106978 54505
rect 106922 54431 106978 54440
rect 108302 54496 108358 54505
rect 108302 54431 108358 54440
rect 104808 51740 104860 51746
rect 104808 51682 104860 51688
rect 104162 28248 104218 28257
rect 104162 28183 104218 28192
rect 104176 15978 104204 28183
rect 104164 15972 104216 15978
rect 104164 15914 104216 15920
rect 104820 6914 104848 51682
rect 106936 17270 106964 54431
rect 107568 49088 107620 49094
rect 107568 49030 107620 49036
rect 106924 17264 106976 17270
rect 106924 17206 106976 17212
rect 105542 15872 105598 15881
rect 105542 15807 105598 15816
rect 103348 6886 103468 6914
rect 104544 6886 104848 6914
rect 102232 3596 102284 3602
rect 102232 3538 102284 3544
rect 97448 3528 97500 3534
rect 97448 3470 97500 3476
rect 97908 3528 97960 3534
rect 97908 3470 97960 3476
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 99288 3528 99340 3534
rect 99288 3470 99340 3476
rect 99840 3528 99892 3534
rect 99840 3470 99892 3476
rect 100668 3528 100720 3534
rect 100668 3470 100720 3476
rect 101036 3528 101088 3534
rect 101036 3470 101088 3476
rect 102048 3528 102100 3534
rect 102048 3470 102100 3476
rect 97460 480 97488 3470
rect 98656 480 98684 3470
rect 99852 480 99880 3470
rect 101048 480 101076 3470
rect 102244 480 102272 3538
rect 103348 480 103376 6886
rect 104544 480 104572 6886
rect 105556 3466 105584 15807
rect 107580 3534 107608 49030
rect 106924 3528 106976 3534
rect 106924 3470 106976 3476
rect 107568 3528 107620 3534
rect 107568 3470 107620 3476
rect 108120 3528 108172 3534
rect 108120 3470 108172 3476
rect 105544 3460 105596 3466
rect 105544 3402 105596 3408
rect 105728 3460 105780 3466
rect 105728 3402 105780 3408
rect 105740 480 105768 3402
rect 106936 480 106964 3470
rect 108132 480 108160 3470
rect 108316 3369 108344 54431
rect 111616 22840 111668 22846
rect 111616 22782 111668 22788
rect 110328 11824 110380 11830
rect 110328 11766 110380 11772
rect 108948 10396 109000 10402
rect 108948 10338 109000 10344
rect 108960 3534 108988 10338
rect 110340 3534 110368 11766
rect 108948 3528 109000 3534
rect 108948 3470 109000 3476
rect 109316 3528 109368 3534
rect 109316 3470 109368 3476
rect 110328 3528 110380 3534
rect 110328 3470 110380 3476
rect 110512 3528 110564 3534
rect 110512 3470 110564 3476
rect 108302 3360 108358 3369
rect 108302 3295 108358 3304
rect 109328 480 109356 3470
rect 110524 480 110552 3470
rect 111628 480 111656 22782
rect 111720 3534 111748 55791
rect 112444 20188 112496 20194
rect 112444 20130 112496 20136
rect 112456 6254 112484 20130
rect 113100 6914 113128 70994
rect 115860 62082 115888 91151
rect 116584 91112 116636 91118
rect 116584 91054 116636 91060
rect 116596 74526 116624 91054
rect 116584 74520 116636 74526
rect 116584 74462 116636 74468
rect 116582 64288 116638 64297
rect 116582 64223 116638 64232
rect 115848 62076 115900 62082
rect 115848 62018 115900 62024
rect 115848 44872 115900 44878
rect 115848 44814 115900 44820
rect 114560 26988 114612 26994
rect 114560 26930 114612 26936
rect 114572 20194 114600 26930
rect 114560 20188 114612 20194
rect 114560 20130 114612 20136
rect 112824 6886 113128 6914
rect 112444 6248 112496 6254
rect 112444 6190 112496 6196
rect 111708 3528 111760 3534
rect 111708 3470 111760 3476
rect 112824 480 112852 6886
rect 114008 6248 114060 6254
rect 114008 6190 114060 6196
rect 114020 480 114048 6190
rect 115860 3534 115888 44814
rect 116596 17338 116624 64223
rect 117240 52426 117268 91151
rect 118528 77178 118556 91287
rect 118606 91216 118662 91225
rect 118606 91151 118662 91160
rect 119986 91216 120042 91225
rect 119986 91151 120042 91160
rect 121366 91216 121422 91225
rect 121366 91151 121422 91160
rect 122746 91216 122802 91225
rect 122746 91151 122802 91160
rect 118516 77172 118568 77178
rect 118516 77114 118568 77120
rect 118620 53786 118648 91151
rect 120000 71738 120028 91151
rect 121380 75886 121408 91151
rect 122196 89004 122248 89010
rect 122196 88946 122248 88952
rect 122102 82240 122158 82249
rect 122102 82175 122158 82184
rect 121368 75880 121420 75886
rect 121368 75822 121420 75828
rect 119988 71732 120040 71738
rect 119988 71674 120040 71680
rect 119988 69692 120040 69698
rect 119988 69634 120040 69640
rect 118608 53780 118660 53786
rect 118608 53722 118660 53728
rect 117228 52420 117280 52426
rect 117228 52362 117280 52368
rect 119896 46300 119948 46306
rect 119896 46242 119948 46248
rect 118608 31068 118660 31074
rect 118608 31010 118660 31016
rect 117228 24200 117280 24206
rect 117228 24142 117280 24148
rect 116584 17332 116636 17338
rect 116584 17274 116636 17280
rect 117240 3534 117268 24142
rect 118620 3534 118648 31010
rect 119908 16574 119936 46242
rect 119816 16546 119936 16574
rect 119816 3534 119844 16546
rect 120000 6914 120028 69634
rect 119908 6886 120028 6914
rect 115204 3528 115256 3534
rect 115204 3470 115256 3476
rect 115848 3528 115900 3534
rect 115848 3470 115900 3476
rect 116400 3528 116452 3534
rect 116400 3470 116452 3476
rect 117228 3528 117280 3534
rect 117228 3470 117280 3476
rect 117596 3528 117648 3534
rect 117596 3470 117648 3476
rect 118608 3528 118660 3534
rect 118608 3470 118660 3476
rect 118792 3528 118844 3534
rect 118792 3470 118844 3476
rect 119804 3528 119856 3534
rect 119804 3470 119856 3476
rect 115216 480 115244 3470
rect 116412 480 116440 3470
rect 117608 480 117636 3470
rect 118804 480 118832 3470
rect 119908 480 119936 6886
rect 122116 3602 122144 82175
rect 122208 80034 122236 88946
rect 122760 84017 122788 91151
rect 122852 89690 122880 91287
rect 124126 91216 124182 91225
rect 124126 91151 124182 91160
rect 122840 89684 122892 89690
rect 122840 89626 122892 89632
rect 122746 84008 122802 84017
rect 122746 83943 122802 83952
rect 122196 80028 122248 80034
rect 122196 79970 122248 79976
rect 124140 73098 124168 91151
rect 125428 85542 125456 91287
rect 125506 91216 125562 91225
rect 125506 91151 125562 91160
rect 125416 85536 125468 85542
rect 125416 85478 125468 85484
rect 125520 78606 125548 91151
rect 126624 86601 126652 91831
rect 126900 91798 126928 92239
rect 130750 92032 130806 92041
rect 130750 91967 130806 91976
rect 126888 91792 126940 91798
rect 126888 91734 126940 91740
rect 126886 91624 126942 91633
rect 126886 91559 126942 91568
rect 126702 91352 126758 91361
rect 126702 91287 126758 91296
rect 126610 86592 126666 86601
rect 126610 86527 126666 86536
rect 125508 78600 125560 78606
rect 125508 78542 125560 78548
rect 124128 73092 124180 73098
rect 124128 73034 124180 73040
rect 126716 63510 126744 91287
rect 126794 91216 126850 91225
rect 126794 91151 126850 91160
rect 126704 63504 126756 63510
rect 126704 63446 126756 63452
rect 126808 59294 126836 91151
rect 126796 59288 126848 59294
rect 126796 59230 126848 59236
rect 126900 56574 126928 91559
rect 127990 91216 128046 91225
rect 127990 91151 128046 91160
rect 129646 91216 129702 91225
rect 129646 91151 129702 91160
rect 128004 91118 128032 91151
rect 127992 91112 128044 91118
rect 127992 91054 128044 91060
rect 129004 91112 129056 91118
rect 129004 91054 129056 91060
rect 129016 60654 129044 91054
rect 129660 70378 129688 91151
rect 130764 90409 130792 91967
rect 151634 91352 151690 91361
rect 151634 91287 151690 91296
rect 133786 91216 133842 91225
rect 133786 91151 133842 91160
rect 134430 91216 134486 91225
rect 134430 91151 134486 91160
rect 134708 91180 134760 91186
rect 130750 90400 130806 90409
rect 130750 90335 130806 90344
rect 129648 70372 129700 70378
rect 129648 70314 129700 70320
rect 133800 68950 133828 91151
rect 134444 87961 134472 91151
rect 134708 91122 134760 91128
rect 134720 88262 134748 91122
rect 151082 90400 151138 90409
rect 151082 90335 151138 90344
rect 134708 88256 134760 88262
rect 134708 88198 134760 88204
rect 134430 87952 134486 87961
rect 134430 87887 134486 87896
rect 151096 81326 151124 90335
rect 151648 85474 151676 91287
rect 151726 91216 151782 91225
rect 151726 91151 151782 91160
rect 153106 91216 153162 91225
rect 153106 91151 153162 91160
rect 151636 85468 151688 85474
rect 151636 85410 151688 85416
rect 151084 81320 151136 81326
rect 151084 81262 151136 81268
rect 151740 79966 151768 91151
rect 151728 79960 151780 79966
rect 151728 79902 151780 79908
rect 151082 76800 151138 76809
rect 151082 76735 151138 76744
rect 133788 68944 133840 68950
rect 133788 68886 133840 68892
rect 147034 67008 147090 67017
rect 147034 66943 147090 66952
rect 129004 60648 129056 60654
rect 129004 60590 129056 60596
rect 126888 56568 126940 56574
rect 126888 56510 126940 56516
rect 126244 46232 126296 46238
rect 126244 46174 126296 46180
rect 124128 32428 124180 32434
rect 124128 32370 124180 32376
rect 122748 29708 122800 29714
rect 122748 29650 122800 29656
rect 122104 3596 122156 3602
rect 122104 3538 122156 3544
rect 122760 3534 122788 29650
rect 124140 3534 124168 32370
rect 125508 21480 125560 21486
rect 125508 21422 125560 21428
rect 125520 3534 125548 21422
rect 126256 3641 126284 46174
rect 146944 39364 146996 39370
rect 146944 39306 146996 39312
rect 142804 33856 142856 33862
rect 142804 33798 142856 33804
rect 130384 28348 130436 28354
rect 130384 28290 130436 28296
rect 126242 3632 126298 3641
rect 126242 3567 126298 3576
rect 130396 3534 130424 28290
rect 142816 10402 142844 33798
rect 142804 10396 142856 10402
rect 142804 10338 142856 10344
rect 132958 10296 133014 10305
rect 132958 10231 133014 10240
rect 122288 3528 122340 3534
rect 121090 3496 121146 3505
rect 122288 3470 122340 3476
rect 122748 3528 122800 3534
rect 122748 3470 122800 3476
rect 123484 3528 123536 3534
rect 123484 3470 123536 3476
rect 124128 3528 124180 3534
rect 124128 3470 124180 3476
rect 124680 3528 124732 3534
rect 124680 3470 124732 3476
rect 125508 3528 125560 3534
rect 125508 3470 125560 3476
rect 129372 3528 129424 3534
rect 129372 3470 129424 3476
rect 130384 3528 130436 3534
rect 130384 3470 130436 3476
rect 121090 3431 121146 3440
rect 121104 480 121132 3431
rect 122300 480 122328 3470
rect 123496 480 123524 3470
rect 124692 480 124720 3470
rect 125874 3360 125930 3369
rect 125874 3295 125930 3304
rect 125888 480 125916 3295
rect 129384 480 129412 3470
rect 132972 480 133000 10231
rect 146956 4894 146984 39306
rect 147048 33794 147076 66943
rect 151096 56001 151124 76735
rect 153120 74458 153148 91151
rect 158732 89622 158760 93055
rect 162872 92410 162900 94386
rect 162860 92404 162912 92410
rect 162860 92346 162912 92352
rect 164148 91792 164200 91798
rect 164148 91734 164200 91740
rect 163502 90400 163558 90409
rect 163502 90335 163558 90344
rect 158720 89616 158772 89622
rect 158720 89558 158772 89564
rect 162214 89040 162270 89049
rect 160100 89004 160152 89010
rect 162214 88975 162270 88984
rect 160100 88946 160152 88952
rect 160112 85474 160140 88946
rect 160100 85468 160152 85474
rect 160100 85410 160152 85416
rect 160744 84856 160796 84862
rect 160744 84798 160796 84804
rect 153108 74452 153160 74458
rect 153108 74394 153160 74400
rect 151082 55992 151138 56001
rect 151082 55927 151138 55936
rect 151082 40624 151138 40633
rect 151082 40559 151138 40568
rect 147036 33788 147088 33794
rect 147036 33730 147088 33736
rect 151096 26926 151124 40559
rect 160756 39438 160784 84798
rect 162228 81326 162256 88975
rect 162216 81320 162268 81326
rect 162216 81262 162268 81268
rect 162124 80708 162176 80714
rect 162124 80650 162176 80656
rect 160744 39432 160796 39438
rect 160744 39374 160796 39380
rect 151084 26920 151136 26926
rect 151084 26862 151136 26868
rect 162136 9042 162164 80650
rect 163516 80034 163544 90335
rect 164160 88262 164188 91734
rect 164148 88256 164200 88262
rect 164148 88198 164200 88204
rect 164896 86737 164924 123422
rect 166264 121508 166316 121514
rect 166264 121450 166316 121456
rect 164976 100020 165028 100026
rect 164976 99962 165028 99968
rect 164988 92177 165016 99962
rect 165528 96688 165580 96694
rect 165528 96630 165580 96636
rect 165540 95169 165568 96630
rect 165620 96008 165672 96014
rect 165620 95950 165672 95956
rect 165526 95160 165582 95169
rect 165526 95095 165582 95104
rect 165632 94450 165660 95950
rect 165620 94444 165672 94450
rect 165620 94386 165672 94392
rect 166276 93226 166304 121450
rect 166356 106344 166408 106350
rect 166356 106286 166408 106292
rect 166264 93220 166316 93226
rect 166264 93162 166316 93168
rect 164974 92168 165030 92177
rect 164974 92103 165030 92112
rect 166368 88233 166396 106286
rect 166448 101448 166500 101454
rect 166448 101390 166500 101396
rect 166354 88224 166410 88233
rect 166354 88159 166410 88168
rect 164976 87644 165028 87650
rect 164976 87586 165028 87592
rect 164882 86728 164938 86737
rect 164882 86663 164938 86672
rect 163504 80028 163556 80034
rect 163504 79970 163556 79976
rect 164988 74361 165016 87586
rect 166460 85542 166488 101390
rect 166448 85536 166500 85542
rect 166448 85478 166500 85484
rect 167656 82754 167684 135254
rect 167748 109041 167776 137226
rect 167828 113212 167880 113218
rect 167828 113154 167880 113160
rect 167734 109032 167790 109041
rect 167734 108967 167790 108976
rect 167736 104916 167788 104922
rect 167736 104858 167788 104864
rect 167644 82748 167696 82754
rect 167644 82690 167696 82696
rect 167748 77246 167776 104858
rect 167840 85241 167868 113154
rect 168288 111784 168340 111790
rect 168286 111752 168288 111761
rect 168340 111752 168342 111761
rect 168286 111687 168342 111696
rect 168010 111072 168066 111081
rect 168010 111007 168066 111016
rect 167920 110424 167972 110430
rect 167918 110392 167920 110401
rect 167972 110392 167974 110401
rect 167918 110327 167974 110336
rect 168024 103514 168052 111007
rect 167932 103486 168052 103514
rect 167932 87961 167960 103486
rect 167918 87952 167974 87961
rect 167918 87887 167974 87896
rect 167826 85232 167882 85241
rect 167826 85167 167882 85176
rect 167736 77240 167788 77246
rect 167736 77182 167788 77188
rect 164974 74352 165030 74361
rect 164974 74287 165030 74296
rect 168392 28354 168420 251194
rect 168484 237425 168512 447335
rect 171140 432608 171192 432614
rect 171140 432550 171192 432556
rect 169760 400240 169812 400246
rect 169760 400182 169812 400188
rect 169024 353388 169076 353394
rect 169024 353330 169076 353336
rect 168470 237416 168526 237425
rect 168470 237351 168526 237360
rect 169036 222902 169064 353330
rect 169114 331528 169170 331537
rect 169114 331463 169170 331472
rect 169128 272542 169156 331463
rect 169772 295322 169800 400182
rect 170404 367804 170456 367810
rect 170404 367746 170456 367752
rect 170416 298353 170444 367746
rect 170496 332648 170548 332654
rect 170496 332590 170548 332596
rect 170508 309806 170536 332590
rect 170496 309800 170548 309806
rect 170496 309742 170548 309748
rect 170402 298344 170458 298353
rect 170402 298279 170458 298288
rect 170416 296714 170444 298279
rect 170416 296686 170536 296714
rect 169760 295316 169812 295322
rect 169760 295258 169812 295264
rect 169772 294642 169800 295258
rect 169760 294636 169812 294642
rect 169760 294578 169812 294584
rect 170404 293276 170456 293282
rect 170404 293218 170456 293224
rect 169208 274712 169260 274718
rect 169208 274654 169260 274660
rect 169116 272536 169168 272542
rect 169116 272478 169168 272484
rect 169220 247790 169248 274654
rect 169208 247784 169260 247790
rect 169208 247726 169260 247732
rect 170416 241505 170444 293218
rect 170508 253201 170536 296686
rect 171048 256760 171100 256766
rect 171048 256702 171100 256708
rect 170494 253192 170550 253201
rect 170494 253127 170550 253136
rect 170954 247072 171010 247081
rect 170954 247007 171010 247016
rect 170402 241496 170458 241505
rect 170402 241431 170458 241440
rect 170968 233889 170996 247007
rect 170954 233880 171010 233889
rect 170954 233815 171010 233824
rect 169024 222896 169076 222902
rect 169024 222838 169076 222844
rect 170402 213344 170458 213353
rect 170402 213279 170458 213288
rect 169116 180940 169168 180946
rect 169116 180882 169168 180888
rect 168470 174856 168526 174865
rect 168470 174791 168526 174800
rect 168484 172514 168512 174791
rect 168472 172508 168524 172514
rect 168472 172450 168524 172456
rect 169022 171320 169078 171329
rect 169022 171255 169078 171264
rect 169036 151094 169064 171255
rect 169128 171018 169156 180882
rect 169116 171012 169168 171018
rect 169116 170954 169168 170960
rect 170416 163538 170444 213279
rect 171060 202162 171088 256702
rect 171152 247081 171180 432550
rect 171232 396092 171284 396098
rect 171232 396034 171284 396040
rect 171244 268394 171272 396034
rect 176016 357536 176068 357542
rect 176016 357478 176068 357484
rect 175922 343904 175978 343913
rect 175922 343839 175978 343848
rect 173348 342372 173400 342378
rect 173348 342314 173400 342320
rect 171782 341048 171838 341057
rect 171782 340983 171838 340992
rect 171232 268388 171284 268394
rect 171232 268330 171284 268336
rect 171138 247072 171194 247081
rect 171138 247007 171194 247016
rect 171048 202156 171100 202162
rect 171048 202098 171100 202104
rect 170496 182300 170548 182306
rect 170496 182242 170548 182248
rect 170404 163532 170456 163538
rect 170404 163474 170456 163480
rect 170508 158710 170536 182242
rect 170496 158704 170548 158710
rect 170496 158646 170548 158652
rect 169024 151088 169076 151094
rect 169024 151030 169076 151036
rect 171796 145586 171824 340983
rect 173256 334076 173308 334082
rect 173256 334018 173308 334024
rect 173164 316804 173216 316810
rect 173164 316746 173216 316752
rect 172428 268388 172480 268394
rect 172428 268330 172480 268336
rect 172440 267889 172468 268330
rect 172426 267880 172482 267889
rect 172426 267815 172482 267824
rect 171876 264988 171928 264994
rect 171876 264930 171928 264936
rect 171888 213858 171916 264930
rect 173176 255513 173204 316746
rect 173268 278050 173296 334018
rect 173360 311166 173388 342314
rect 174634 339824 174690 339833
rect 174634 339759 174690 339768
rect 174542 336016 174598 336025
rect 174542 335951 174598 335960
rect 173348 311160 173400 311166
rect 173348 311102 173400 311108
rect 174556 300121 174584 335951
rect 174542 300112 174598 300121
rect 174542 300047 174598 300056
rect 174544 289944 174596 289950
rect 174544 289886 174596 289892
rect 174556 285666 174584 289886
rect 174544 285660 174596 285666
rect 174544 285602 174596 285608
rect 173348 282260 173400 282266
rect 173348 282202 173400 282208
rect 173256 278044 173308 278050
rect 173256 277986 173308 277992
rect 173256 260908 173308 260914
rect 173256 260850 173308 260856
rect 173162 255504 173218 255513
rect 173162 255439 173218 255448
rect 173164 248940 173216 248946
rect 173164 248882 173216 248888
rect 172518 241768 172574 241777
rect 172518 241703 172574 241712
rect 172532 236042 172560 241703
rect 172440 236014 172560 236042
rect 172440 230353 172468 236014
rect 172426 230344 172482 230353
rect 172426 230279 172482 230288
rect 172426 228440 172482 228449
rect 172426 228375 172482 228384
rect 172440 220794 172468 228375
rect 173176 226302 173204 248882
rect 173268 235793 173296 260850
rect 173254 235784 173310 235793
rect 173254 235719 173310 235728
rect 173360 229022 173388 282202
rect 173440 279472 173492 279478
rect 173440 279414 173492 279420
rect 173452 256766 173480 279414
rect 174544 270564 174596 270570
rect 174544 270506 174596 270512
rect 173440 256760 173492 256766
rect 173440 256702 173492 256708
rect 174176 248464 174228 248470
rect 174176 248406 174228 248412
rect 174188 243574 174216 248406
rect 174176 243568 174228 243574
rect 174176 243510 174228 243516
rect 173348 229016 173400 229022
rect 173348 228958 173400 228964
rect 173714 227760 173770 227769
rect 173714 227695 173770 227704
rect 173164 226296 173216 226302
rect 173164 226238 173216 226244
rect 173348 226296 173400 226302
rect 173348 226238 173400 226244
rect 172428 220788 172480 220794
rect 172428 220730 172480 220736
rect 171876 213852 171928 213858
rect 171876 213794 171928 213800
rect 171968 213240 172020 213246
rect 171968 213182 172020 213188
rect 171980 209545 172008 213182
rect 171966 209536 172022 209545
rect 171966 209471 172022 209480
rect 173256 202224 173308 202230
rect 173256 202166 173308 202172
rect 173162 187096 173218 187105
rect 173162 187031 173218 187040
rect 171874 178256 171930 178265
rect 171874 178191 171930 178200
rect 171888 162858 171916 178191
rect 171876 162852 171928 162858
rect 171876 162794 171928 162800
rect 171784 145580 171836 145586
rect 171784 145522 171836 145528
rect 171784 133952 171836 133958
rect 171784 133894 171836 133900
rect 170494 117328 170550 117337
rect 170494 117263 170550 117272
rect 170404 108316 170456 108322
rect 170404 108258 170456 108264
rect 169116 104168 169168 104174
rect 169116 104110 169168 104116
rect 169022 101416 169078 101425
rect 169022 101351 169078 101360
rect 168656 95940 168708 95946
rect 168656 95882 168708 95888
rect 168668 93129 168696 95882
rect 168654 93120 168710 93129
rect 168654 93055 168710 93064
rect 169036 81433 169064 101351
rect 169128 86873 169156 104110
rect 169114 86864 169170 86873
rect 169114 86799 169170 86808
rect 169022 81424 169078 81433
rect 169022 81359 169078 81368
rect 170416 78606 170444 108258
rect 170508 89593 170536 117263
rect 170680 116612 170732 116618
rect 170680 116554 170732 116560
rect 170588 93220 170640 93226
rect 170588 93162 170640 93168
rect 170494 89584 170550 89593
rect 170494 89519 170550 89528
rect 170404 78600 170456 78606
rect 170404 78542 170456 78548
rect 170600 67590 170628 93162
rect 170692 90982 170720 116554
rect 170680 90976 170732 90982
rect 170680 90918 170732 90924
rect 171796 88097 171824 133894
rect 172060 110492 172112 110498
rect 172060 110434 172112 110440
rect 171968 103556 172020 103562
rect 171968 103498 172020 103504
rect 171876 98048 171928 98054
rect 171876 97990 171928 97996
rect 171782 88088 171838 88097
rect 171782 88023 171838 88032
rect 170588 67584 170640 67590
rect 170588 67526 170640 67532
rect 171888 66162 171916 97990
rect 171980 74497 172008 103498
rect 172072 93673 172100 110434
rect 172058 93664 172114 93673
rect 172058 93599 172114 93608
rect 171966 74488 172022 74497
rect 171966 74423 172022 74432
rect 171876 66156 171928 66162
rect 171876 66098 171928 66104
rect 168380 28348 168432 28354
rect 168380 28290 168432 28296
rect 162124 9036 162176 9042
rect 162124 8978 162176 8984
rect 146944 4888 146996 4894
rect 136454 4856 136510 4865
rect 146944 4830 146996 4836
rect 136454 4791 136510 4800
rect 136468 480 136496 4791
rect 173176 4049 173204 187031
rect 173268 138718 173296 202166
rect 173360 173913 173388 226238
rect 173728 223553 173756 227695
rect 173714 223544 173770 223553
rect 173714 223479 173770 223488
rect 173440 178084 173492 178090
rect 173440 178026 173492 178032
rect 173346 173904 173402 173913
rect 173346 173839 173402 173848
rect 173452 165578 173480 178026
rect 173440 165572 173492 165578
rect 173440 165514 173492 165520
rect 173256 138712 173308 138718
rect 173256 138654 173308 138660
rect 173348 133204 173400 133210
rect 173348 133146 173400 133152
rect 173256 131164 173308 131170
rect 173256 131106 173308 131112
rect 173268 86601 173296 131106
rect 173360 92478 173388 133146
rect 173440 113280 173492 113286
rect 173440 113222 173492 113228
rect 173348 92472 173400 92478
rect 173348 92414 173400 92420
rect 173254 86592 173310 86601
rect 173254 86527 173310 86536
rect 173452 75886 173480 113222
rect 173440 75880 173492 75886
rect 173440 75822 173492 75828
rect 174556 50454 174584 270506
rect 174648 152522 174676 339759
rect 174728 305720 174780 305726
rect 174728 305662 174780 305668
rect 174740 281450 174768 305662
rect 174728 281444 174780 281450
rect 174728 281386 174780 281392
rect 175188 278792 175240 278798
rect 175188 278734 175240 278740
rect 175200 277370 175228 278734
rect 175188 277364 175240 277370
rect 175188 277306 175240 277312
rect 175832 256760 175884 256766
rect 175832 256702 175884 256708
rect 175844 253910 175872 256702
rect 175832 253904 175884 253910
rect 175832 253846 175884 253852
rect 174728 250504 174780 250510
rect 174728 250446 174780 250452
rect 174740 226234 174768 250446
rect 174728 226228 174780 226234
rect 174728 226170 174780 226176
rect 175936 160721 175964 343839
rect 176028 322318 176056 357478
rect 177396 350600 177448 350606
rect 177396 350542 177448 350548
rect 177302 330032 177358 330041
rect 177302 329967 177358 329976
rect 176016 322312 176068 322318
rect 176016 322254 176068 322260
rect 176014 319424 176070 319433
rect 176014 319359 176070 319368
rect 176028 297537 176056 319359
rect 176014 297528 176070 297537
rect 176014 297463 176070 297472
rect 176014 284608 176070 284617
rect 176014 284543 176070 284552
rect 176028 230450 176056 284543
rect 176108 249824 176160 249830
rect 176108 249766 176160 249772
rect 176120 235278 176148 249766
rect 176108 235272 176160 235278
rect 176108 235214 176160 235220
rect 176660 231736 176712 231742
rect 176660 231678 176712 231684
rect 176672 231130 176700 231678
rect 176660 231124 176712 231130
rect 176660 231066 176712 231072
rect 176016 230444 176068 230450
rect 176016 230386 176068 230392
rect 176014 182200 176070 182209
rect 176014 182135 176070 182144
rect 175922 160712 175978 160721
rect 175922 160647 175978 160656
rect 176028 157350 176056 182135
rect 176016 157344 176068 157350
rect 176016 157286 176068 157292
rect 174636 152516 174688 152522
rect 174636 152458 174688 152464
rect 175924 142860 175976 142866
rect 175924 142802 175976 142808
rect 174636 112464 174688 112470
rect 174636 112406 174688 112412
rect 174648 73098 174676 112406
rect 174728 102196 174780 102202
rect 174728 102138 174780 102144
rect 174740 85377 174768 102138
rect 175936 94081 175964 142802
rect 176016 131776 176068 131782
rect 176016 131718 176068 131724
rect 175922 94072 175978 94081
rect 175922 94007 175978 94016
rect 175924 90364 175976 90370
rect 175924 90306 175976 90312
rect 174726 85368 174782 85377
rect 174726 85303 174782 85312
rect 174636 73092 174688 73098
rect 174636 73034 174688 73040
rect 175936 70378 175964 90306
rect 176028 89010 176056 131718
rect 176016 89004 176068 89010
rect 176016 88946 176068 88952
rect 175924 70372 175976 70378
rect 175924 70314 175976 70320
rect 174544 50448 174596 50454
rect 174544 50390 174596 50396
rect 177316 6225 177344 329967
rect 177408 267034 177436 350542
rect 177488 328500 177540 328506
rect 177488 328442 177540 328448
rect 177500 285054 177528 328442
rect 178052 289105 178080 460906
rect 179420 451308 179472 451314
rect 179420 451250 179472 451256
rect 178682 353560 178738 353569
rect 178682 353495 178738 353504
rect 178696 320890 178724 353495
rect 178776 336864 178828 336870
rect 178776 336806 178828 336812
rect 178684 320884 178736 320890
rect 178684 320826 178736 320832
rect 178788 316810 178816 336806
rect 178776 316804 178828 316810
rect 178776 316746 178828 316752
rect 178682 293992 178738 294001
rect 178682 293927 178738 293936
rect 178038 289096 178094 289105
rect 178038 289031 178094 289040
rect 177488 285048 177540 285054
rect 177488 284990 177540 284996
rect 177396 267028 177448 267034
rect 177396 266970 177448 266976
rect 177856 265192 177908 265198
rect 177856 265134 177908 265140
rect 177396 253224 177448 253230
rect 177396 253166 177448 253172
rect 177408 236609 177436 253166
rect 177394 236600 177450 236609
rect 177394 236535 177450 236544
rect 177868 231130 177896 265134
rect 178696 264246 178724 293927
rect 178776 283892 178828 283898
rect 178776 283834 178828 283840
rect 178788 271182 178816 283834
rect 178776 271176 178828 271182
rect 178776 271118 178828 271124
rect 178868 269204 178920 269210
rect 178868 269146 178920 269152
rect 178684 264240 178736 264246
rect 178684 264182 178736 264188
rect 178684 262336 178736 262342
rect 178684 262278 178736 262284
rect 177948 233912 178000 233918
rect 177948 233854 178000 233860
rect 177856 231124 177908 231130
rect 177856 231066 177908 231072
rect 177394 207768 177450 207777
rect 177394 207703 177450 207712
rect 177408 155242 177436 207703
rect 177960 184210 177988 233854
rect 178696 229094 178724 262278
rect 178776 256080 178828 256086
rect 178776 256022 178828 256028
rect 178788 233918 178816 256022
rect 178880 248946 178908 269146
rect 178960 249824 179012 249830
rect 178960 249766 179012 249772
rect 178868 248940 178920 248946
rect 178868 248882 178920 248888
rect 178972 237017 179000 249766
rect 178958 237008 179014 237017
rect 178958 236943 179014 236952
rect 179432 235657 179460 451250
rect 202142 446040 202198 446049
rect 202142 445975 202198 445984
rect 188344 375420 188396 375426
rect 188344 375362 188396 375368
rect 185582 371376 185638 371385
rect 185582 371311 185638 371320
rect 181536 363044 181588 363050
rect 181536 362986 181588 362992
rect 181442 352064 181498 352073
rect 181442 351999 181498 352008
rect 180062 346624 180118 346633
rect 180062 346559 180118 346568
rect 180076 305697 180104 346559
rect 180156 310548 180208 310554
rect 180156 310490 180208 310496
rect 180062 305688 180118 305697
rect 180062 305623 180118 305632
rect 180064 245676 180116 245682
rect 180064 245618 180116 245624
rect 179418 235648 179474 235657
rect 179418 235583 179474 235592
rect 178776 233912 178828 233918
rect 178776 233854 178828 233860
rect 178696 229090 178908 229094
rect 178684 229084 178908 229090
rect 178736 229066 178908 229084
rect 178684 229026 178736 229032
rect 178684 225616 178736 225622
rect 178684 225558 178736 225564
rect 178696 216578 178724 225558
rect 178684 216572 178736 216578
rect 178684 216514 178736 216520
rect 178040 216504 178092 216510
rect 178040 216446 178092 216452
rect 178052 215393 178080 216446
rect 178038 215384 178094 215393
rect 178038 215319 178094 215328
rect 178682 214840 178738 214849
rect 178682 214775 178738 214784
rect 177948 184204 178000 184210
rect 177948 184146 178000 184152
rect 177486 183832 177542 183841
rect 177486 183767 177542 183776
rect 177500 160070 177528 183767
rect 177488 160064 177540 160070
rect 177488 160006 177540 160012
rect 177396 155236 177448 155242
rect 177396 155178 177448 155184
rect 177396 146328 177448 146334
rect 177396 146270 177448 146276
rect 177408 111081 177436 146270
rect 177394 111072 177450 111081
rect 177394 111007 177450 111016
rect 177578 111072 177634 111081
rect 177578 111007 177634 111016
rect 177394 108352 177450 108361
rect 177394 108287 177450 108296
rect 177408 71738 177436 108287
rect 177488 100768 177540 100774
rect 177488 100710 177540 100716
rect 177500 81297 177528 100710
rect 177592 93226 177620 111007
rect 177580 93220 177632 93226
rect 177580 93162 177632 93168
rect 177486 81288 177542 81297
rect 177486 81223 177542 81232
rect 177396 71732 177448 71738
rect 177396 71674 177448 71680
rect 178696 18698 178724 214775
rect 178776 192500 178828 192506
rect 178776 192442 178828 192448
rect 178788 141438 178816 192442
rect 178880 188358 178908 229066
rect 178868 188352 178920 188358
rect 178868 188294 178920 188300
rect 178868 176792 178920 176798
rect 178868 176734 178920 176740
rect 178880 158030 178908 176734
rect 178868 158024 178920 158030
rect 178868 157966 178920 157972
rect 178868 150476 178920 150482
rect 178868 150418 178920 150424
rect 178776 141432 178828 141438
rect 178776 141374 178828 141380
rect 178776 126268 178828 126274
rect 178776 126210 178828 126216
rect 178788 79966 178816 126210
rect 178880 111790 178908 150418
rect 178868 111784 178920 111790
rect 178868 111726 178920 111732
rect 178868 97300 178920 97306
rect 178868 97242 178920 97248
rect 178776 79960 178828 79966
rect 178776 79902 178828 79908
rect 178880 63442 178908 97242
rect 178868 63436 178920 63442
rect 178868 63378 178920 63384
rect 178684 18692 178736 18698
rect 178684 18634 178736 18640
rect 180076 13025 180104 245618
rect 180168 229090 180196 310490
rect 180248 273284 180300 273290
rect 180248 273226 180300 273232
rect 180260 235958 180288 273226
rect 180248 235952 180300 235958
rect 180248 235894 180300 235900
rect 180156 229084 180208 229090
rect 180156 229026 180208 229032
rect 180260 179382 180288 235894
rect 181456 207777 181484 351999
rect 181548 249121 181576 362986
rect 184296 353320 184348 353326
rect 184296 353262 184348 353268
rect 183008 345160 183060 345166
rect 183008 345102 183060 345108
rect 182822 338464 182878 338473
rect 182822 338399 182878 338408
rect 182836 330449 182864 338399
rect 182822 330440 182878 330449
rect 182822 330375 182878 330384
rect 183020 315353 183048 345102
rect 184204 329112 184256 329118
rect 184204 329054 184256 329060
rect 182822 315344 182878 315353
rect 182822 315279 182878 315288
rect 183006 315344 183062 315353
rect 183006 315279 183062 315288
rect 181626 291272 181682 291281
rect 181626 291207 181682 291216
rect 181640 256018 181668 291207
rect 182088 259480 182140 259486
rect 182088 259422 182140 259428
rect 181628 256012 181680 256018
rect 181628 255954 181680 255960
rect 181534 249112 181590 249121
rect 181534 249047 181590 249056
rect 181996 249076 182048 249082
rect 181996 249018 182048 249024
rect 181534 217288 181590 217297
rect 181534 217223 181590 217232
rect 181442 207768 181498 207777
rect 181442 207703 181498 207712
rect 180248 179376 180300 179382
rect 180248 179318 180300 179324
rect 181442 175400 181498 175409
rect 181442 175335 181498 175344
rect 181456 162790 181484 175335
rect 181444 162784 181496 162790
rect 181444 162726 181496 162732
rect 180156 149728 180208 149734
rect 180156 149670 180208 149676
rect 180168 110430 180196 149670
rect 181548 148374 181576 217223
rect 182008 216714 182036 249018
rect 181996 216708 182048 216714
rect 181996 216650 182048 216656
rect 182100 187105 182128 259422
rect 182836 231713 182864 315279
rect 183468 304292 183520 304298
rect 183468 304234 183520 304240
rect 183480 302326 183508 304234
rect 183468 302320 183520 302326
rect 183468 302262 183520 302268
rect 182914 280936 182970 280945
rect 182914 280871 182970 280880
rect 182822 231704 182878 231713
rect 182822 231639 182878 231648
rect 182928 219337 182956 280871
rect 183480 280158 183508 302262
rect 183468 280152 183520 280158
rect 183468 280094 183520 280100
rect 183100 274712 183152 274718
rect 183100 274654 183152 274660
rect 183008 270564 183060 270570
rect 183008 270506 183060 270512
rect 183020 256086 183048 270506
rect 183112 265198 183140 274654
rect 183100 265192 183152 265198
rect 183100 265134 183152 265140
rect 184216 264926 184244 329054
rect 184308 311234 184336 353262
rect 184296 311228 184348 311234
rect 184296 311170 184348 311176
rect 184388 305040 184440 305046
rect 184388 304982 184440 304988
rect 184296 285048 184348 285054
rect 184296 284990 184348 284996
rect 184204 264920 184256 264926
rect 184204 264862 184256 264868
rect 184204 262268 184256 262274
rect 184204 262210 184256 262216
rect 183468 256760 183520 256766
rect 183468 256702 183520 256708
rect 183008 256080 183060 256086
rect 183008 256022 183060 256028
rect 182914 219328 182970 219337
rect 182914 219263 182970 219272
rect 183480 198014 183508 256702
rect 183468 198008 183520 198014
rect 183468 197950 183520 197956
rect 182824 196648 182876 196654
rect 182824 196590 182876 196596
rect 182086 187096 182142 187105
rect 182086 187031 182142 187040
rect 181536 148368 181588 148374
rect 181536 148310 181588 148316
rect 181444 138032 181496 138038
rect 181444 137974 181496 137980
rect 180340 110560 180392 110566
rect 180340 110502 180392 110508
rect 180156 110424 180208 110430
rect 180156 110366 180208 110372
rect 180248 109064 180300 109070
rect 180248 109006 180300 109012
rect 180260 84114 180288 109006
rect 180352 90409 180380 110502
rect 180338 90400 180394 90409
rect 180338 90335 180394 90344
rect 180248 84108 180300 84114
rect 180248 84050 180300 84056
rect 181456 77178 181484 137974
rect 181536 94512 181588 94518
rect 181536 94454 181588 94460
rect 181548 82793 181576 94454
rect 181534 82784 181590 82793
rect 181534 82719 181590 82728
rect 181444 77172 181496 77178
rect 181444 77114 181496 77120
rect 182836 28354 182864 196590
rect 182914 179616 182970 179625
rect 182914 179551 182970 179560
rect 182928 164218 182956 179551
rect 182916 164212 182968 164218
rect 182916 164154 182968 164160
rect 182916 118720 182968 118726
rect 182916 118662 182968 118668
rect 182928 86902 182956 118662
rect 182916 86896 182968 86902
rect 182916 86838 182968 86844
rect 182824 28348 182876 28354
rect 182824 28290 182876 28296
rect 180062 13016 180118 13025
rect 180062 12951 180118 12960
rect 177302 6216 177358 6225
rect 177302 6151 177358 6160
rect 184216 4894 184244 262210
rect 184308 226302 184336 284990
rect 184400 281518 184428 304982
rect 185596 281625 185624 371311
rect 186964 358896 187016 358902
rect 186964 358838 187016 358844
rect 185768 282192 185820 282198
rect 185768 282134 185820 282140
rect 185582 281616 185638 281625
rect 185780 281586 185808 282134
rect 185582 281551 185638 281560
rect 185768 281580 185820 281586
rect 185768 281522 185820 281528
rect 186228 281580 186280 281586
rect 186228 281522 186280 281528
rect 184388 281512 184440 281518
rect 184388 281454 184440 281460
rect 185584 268388 185636 268394
rect 185584 268330 185636 268336
rect 184848 251864 184900 251870
rect 184848 251806 184900 251812
rect 184860 251258 184888 251806
rect 184848 251252 184900 251258
rect 184848 251194 184900 251200
rect 184388 242208 184440 242214
rect 184388 242150 184440 242156
rect 184400 229770 184428 242150
rect 184388 229764 184440 229770
rect 184388 229706 184440 229712
rect 184296 226296 184348 226302
rect 184296 226238 184348 226244
rect 184294 214024 184350 214033
rect 184294 213959 184350 213968
rect 184308 206922 184336 213959
rect 184296 206916 184348 206922
rect 184296 206858 184348 206864
rect 184294 198112 184350 198121
rect 184294 198047 184350 198056
rect 184308 126342 184336 198047
rect 184860 182850 184888 251194
rect 185596 224942 185624 268330
rect 185676 260976 185728 260982
rect 185676 260918 185728 260924
rect 185688 233306 185716 260918
rect 185676 233300 185728 233306
rect 185676 233242 185728 233248
rect 185584 224936 185636 224942
rect 185584 224878 185636 224884
rect 185596 219434 185624 224878
rect 185688 224233 185716 233242
rect 185674 224224 185730 224233
rect 185674 224159 185730 224168
rect 185596 219406 185716 219434
rect 185584 195288 185636 195294
rect 185584 195230 185636 195236
rect 184848 182844 184900 182850
rect 184848 182786 184900 182792
rect 184388 179512 184440 179518
rect 184388 179454 184440 179460
rect 184400 166938 184428 179454
rect 184388 166932 184440 166938
rect 184388 166874 184440 166880
rect 184296 126336 184348 126342
rect 184296 126278 184348 126284
rect 184388 124908 184440 124914
rect 184388 124850 184440 124856
rect 184296 118788 184348 118794
rect 184296 118730 184348 118736
rect 184308 89729 184336 118730
rect 184400 97209 184428 124850
rect 184386 97200 184442 97209
rect 184386 97135 184442 97144
rect 184388 93220 184440 93226
rect 184388 93162 184440 93168
rect 184294 89720 184350 89729
rect 184294 89655 184350 89664
rect 184400 69018 184428 93162
rect 184388 69012 184440 69018
rect 184388 68954 184440 68960
rect 185596 29646 185624 195230
rect 185688 175166 185716 219406
rect 186240 195294 186268 281522
rect 186976 266354 187004 358838
rect 187054 347984 187110 347993
rect 187054 347919 187110 347928
rect 187068 313342 187096 347919
rect 187056 313336 187108 313342
rect 187056 313278 187108 313284
rect 187608 313336 187660 313342
rect 187608 313278 187660 313284
rect 187054 295488 187110 295497
rect 187054 295423 187110 295432
rect 187068 286346 187096 295423
rect 187620 286346 187648 313278
rect 187056 286340 187108 286346
rect 187056 286282 187108 286288
rect 187608 286340 187660 286346
rect 187608 286282 187660 286288
rect 187056 277432 187108 277438
rect 187056 277374 187108 277380
rect 186964 266348 187016 266354
rect 186964 266290 187016 266296
rect 186962 247616 187018 247625
rect 186962 247551 187018 247560
rect 186976 198694 187004 247551
rect 187068 233238 187096 277374
rect 187146 276040 187202 276049
rect 187146 275975 187202 275984
rect 187160 234433 187188 275975
rect 188356 271969 188384 375362
rect 201500 372700 201552 372706
rect 201500 372642 201552 372648
rect 188436 369912 188488 369918
rect 188436 369854 188488 369860
rect 195334 369880 195390 369889
rect 188342 271960 188398 271969
rect 188342 271895 188398 271904
rect 188342 266384 188398 266393
rect 188342 266319 188398 266328
rect 187240 255332 187292 255338
rect 187240 255274 187292 255280
rect 187146 234424 187202 234433
rect 187146 234359 187202 234368
rect 187056 233232 187108 233238
rect 187056 233174 187108 233180
rect 187252 223514 187280 255274
rect 187240 223508 187292 223514
rect 187240 223450 187292 223456
rect 187252 214713 187280 223450
rect 187054 214704 187110 214713
rect 187054 214639 187110 214648
rect 187238 214704 187294 214713
rect 187238 214639 187294 214648
rect 186964 198688 187016 198694
rect 186964 198630 187016 198636
rect 186976 196654 187004 198630
rect 186964 196648 187016 196654
rect 186964 196590 187016 196596
rect 186228 195288 186280 195294
rect 186228 195230 186280 195236
rect 186962 188456 187018 188465
rect 186962 188391 187018 188400
rect 185766 175536 185822 175545
rect 185766 175471 185822 175480
rect 185676 175160 185728 175166
rect 185676 175102 185728 175108
rect 185780 168298 185808 175471
rect 185768 168292 185820 168298
rect 185768 168234 185820 168240
rect 186976 137358 187004 188391
rect 187068 176050 187096 214639
rect 187056 176044 187108 176050
rect 187056 175986 187108 175992
rect 186964 137352 187016 137358
rect 186964 137294 187016 137300
rect 185676 122868 185728 122874
rect 185676 122810 185728 122816
rect 185688 93158 185716 122810
rect 186964 117972 187016 117978
rect 186964 117914 187016 117920
rect 185676 93152 185728 93158
rect 185676 93094 185728 93100
rect 186976 66230 187004 117914
rect 186964 66224 187016 66230
rect 186964 66166 187016 66172
rect 185584 29640 185636 29646
rect 185584 29582 185636 29588
rect 188356 20058 188384 266319
rect 188448 244390 188476 369854
rect 195334 369815 195390 369824
rect 193864 356176 193916 356182
rect 193864 356118 193916 356124
rect 191104 354816 191156 354822
rect 191104 354758 191156 354764
rect 189724 331288 189776 331294
rect 189724 331230 189776 331236
rect 189736 258126 189764 331230
rect 189816 322312 189868 322318
rect 189816 322254 189868 322260
rect 189828 312594 189856 322254
rect 189816 312588 189868 312594
rect 189816 312530 189868 312536
rect 189814 305688 189870 305697
rect 189814 305623 189870 305632
rect 189724 258120 189776 258126
rect 189724 258062 189776 258068
rect 189724 254584 189776 254590
rect 189724 254526 189776 254532
rect 188528 253972 188580 253978
rect 188528 253914 188580 253920
rect 188436 244384 188488 244390
rect 188436 244326 188488 244332
rect 188436 231124 188488 231130
rect 188436 231066 188488 231072
rect 188448 196761 188476 231066
rect 188540 220697 188568 253914
rect 188988 245744 189040 245750
rect 188988 245686 189040 245692
rect 189000 228313 189028 245686
rect 189080 244316 189132 244322
rect 189080 244258 189132 244264
rect 189092 243001 189120 244258
rect 189078 242992 189134 243001
rect 189078 242927 189134 242936
rect 189736 237386 189764 254526
rect 189724 237380 189776 237386
rect 189724 237322 189776 237328
rect 188986 228304 189042 228313
rect 188986 228239 189042 228248
rect 188526 220688 188582 220697
rect 188526 220623 188582 220632
rect 188434 196752 188490 196761
rect 188434 196687 188490 196696
rect 189722 192536 189778 192545
rect 189722 192471 189778 192480
rect 188434 183696 188490 183705
rect 188434 183631 188490 183640
rect 188448 157282 188476 183631
rect 188436 157276 188488 157282
rect 188436 157218 188488 157224
rect 188434 142216 188490 142225
rect 188434 142151 188490 142160
rect 188448 59294 188476 142151
rect 188528 127016 188580 127022
rect 188528 126958 188580 126964
rect 188540 80073 188568 126958
rect 188526 80064 188582 80073
rect 188526 79999 188582 80008
rect 188436 59288 188488 59294
rect 188436 59230 188488 59236
rect 189736 32502 189764 192471
rect 189828 184385 189856 305623
rect 189908 260160 189960 260166
rect 189908 260102 189960 260108
rect 189920 244390 189948 260102
rect 191116 247042 191144 354758
rect 191196 309800 191248 309806
rect 191196 309742 191248 309748
rect 191104 247036 191156 247042
rect 191104 246978 191156 246984
rect 189908 244384 189960 244390
rect 189908 244326 189960 244332
rect 190368 244316 190420 244322
rect 190368 244258 190420 244264
rect 189908 242956 189960 242962
rect 189908 242898 189960 242904
rect 189920 231742 189948 242898
rect 189908 231736 189960 231742
rect 189908 231678 189960 231684
rect 190380 185706 190408 244258
rect 191208 234530 191236 309742
rect 191288 309188 191340 309194
rect 191288 309130 191340 309136
rect 191300 284306 191328 309130
rect 193128 307896 193180 307902
rect 193128 307838 193180 307844
rect 193034 299840 193090 299849
rect 193034 299775 193090 299784
rect 192574 287600 192630 287609
rect 192574 287535 192630 287544
rect 191288 284300 191340 284306
rect 191288 284242 191340 284248
rect 192484 271924 192536 271930
rect 192484 271866 192536 271872
rect 191748 258528 191800 258534
rect 191748 258470 191800 258476
rect 191760 258126 191788 258470
rect 191748 258120 191800 258126
rect 191748 258062 191800 258068
rect 191288 247784 191340 247790
rect 191288 247726 191340 247732
rect 191196 234524 191248 234530
rect 191196 234466 191248 234472
rect 191300 220794 191328 247726
rect 191656 244384 191708 244390
rect 191656 244326 191708 244332
rect 191288 220788 191340 220794
rect 191288 220730 191340 220736
rect 191196 216708 191248 216714
rect 191196 216650 191248 216656
rect 191104 210588 191156 210594
rect 191104 210530 191156 210536
rect 190368 185700 190420 185706
rect 190368 185642 190420 185648
rect 189814 184376 189870 184385
rect 189814 184311 189870 184320
rect 191116 141506 191144 210530
rect 191208 177313 191236 216650
rect 191668 211138 191696 244326
rect 191656 211132 191708 211138
rect 191656 211074 191708 211080
rect 191760 180033 191788 258062
rect 192496 249762 192524 271866
rect 192588 265674 192616 287535
rect 193048 277001 193076 299775
rect 193140 277370 193168 307838
rect 193876 301374 193904 356118
rect 195242 345264 195298 345273
rect 195242 345199 195298 345208
rect 195256 316713 195284 345199
rect 195242 316704 195298 316713
rect 195242 316639 195298 316648
rect 195242 313304 195298 313313
rect 195242 313239 195298 313248
rect 193864 301368 193916 301374
rect 193864 301310 193916 301316
rect 194508 301368 194560 301374
rect 194508 301310 194560 301316
rect 194520 300898 194548 301310
rect 194508 300892 194560 300898
rect 194508 300834 194560 300840
rect 193956 291304 194008 291310
rect 193956 291246 194008 291252
rect 193864 291236 193916 291242
rect 193864 291178 193916 291184
rect 193128 277364 193180 277370
rect 193128 277306 193180 277312
rect 193140 277166 193168 277306
rect 193128 277160 193180 277166
rect 193128 277102 193180 277108
rect 193034 276992 193090 277001
rect 193034 276927 193090 276936
rect 193036 270632 193088 270638
rect 193036 270574 193088 270580
rect 192576 265668 192628 265674
rect 192576 265610 192628 265616
rect 193048 258074 193076 270574
rect 193128 263628 193180 263634
rect 193128 263570 193180 263576
rect 192956 258046 193076 258074
rect 192576 251320 192628 251326
rect 192576 251262 192628 251268
rect 192484 249756 192536 249762
rect 192484 249698 192536 249704
rect 192588 248414 192616 251262
rect 192956 248441 192984 258046
rect 193036 249756 193088 249762
rect 193036 249698 193088 249704
rect 192496 248386 192616 248414
rect 192942 248432 192998 248441
rect 192496 243137 192524 248386
rect 192942 248367 192998 248376
rect 192576 247716 192628 247722
rect 192576 247658 192628 247664
rect 192482 243128 192538 243137
rect 192482 243063 192538 243072
rect 191840 220108 191892 220114
rect 191840 220050 191892 220056
rect 191852 219337 191880 220050
rect 191838 219328 191894 219337
rect 191838 219263 191894 219272
rect 192496 216753 192524 243063
rect 192588 227662 192616 247658
rect 192956 241534 192984 248367
rect 192944 241528 192996 241534
rect 192944 241470 192996 241476
rect 192576 227656 192628 227662
rect 192576 227598 192628 227604
rect 193048 222970 193076 249698
rect 193036 222964 193088 222970
rect 193036 222906 193088 222912
rect 192482 216744 192538 216753
rect 192482 216679 192538 216688
rect 192576 216708 192628 216714
rect 192576 216650 192628 216656
rect 192588 206990 192616 216650
rect 193034 213208 193090 213217
rect 193034 213143 193090 213152
rect 192576 206984 192628 206990
rect 192576 206926 192628 206932
rect 193048 183161 193076 213143
rect 193140 211818 193168 263570
rect 193876 222057 193904 291178
rect 193968 241505 193996 291246
rect 194048 262948 194100 262954
rect 194048 262890 194100 262896
rect 193954 241496 194010 241505
rect 193954 241431 194010 241440
rect 193862 222048 193918 222057
rect 193862 221983 193918 221992
rect 194060 213217 194088 262890
rect 194520 253910 194548 300834
rect 195060 267028 195112 267034
rect 195060 266970 195112 266976
rect 195072 259418 195100 266970
rect 195060 259412 195112 259418
rect 195060 259354 195112 259360
rect 194508 253904 194560 253910
rect 194508 253846 194560 253852
rect 194140 247104 194192 247110
rect 194140 247046 194192 247052
rect 194046 213208 194102 213217
rect 194046 213143 194102 213152
rect 193128 211812 193180 211818
rect 193128 211754 193180 211760
rect 194152 211070 194180 247046
rect 194506 241496 194562 241505
rect 194506 241431 194562 241440
rect 194520 240553 194548 241431
rect 194506 240544 194562 240553
rect 194506 240479 194562 240488
rect 194520 224330 194548 240479
rect 195058 225584 195114 225593
rect 195058 225519 195114 225528
rect 194508 224324 194560 224330
rect 194508 224266 194560 224272
rect 195072 222154 195100 225519
rect 195152 224256 195204 224262
rect 195152 224198 195204 224204
rect 195164 223582 195192 224198
rect 195152 223576 195204 223582
rect 195152 223518 195204 223524
rect 195152 222896 195204 222902
rect 195152 222838 195204 222844
rect 195164 222154 195192 222838
rect 195060 222148 195112 222154
rect 195060 222090 195112 222096
rect 195152 222148 195204 222154
rect 195152 222090 195204 222096
rect 194690 221776 194746 221785
rect 194690 221711 194746 221720
rect 194704 213897 194732 221711
rect 194690 213888 194746 213897
rect 194690 213823 194746 213832
rect 194784 211880 194836 211886
rect 194784 211822 194836 211828
rect 193128 211064 193180 211070
rect 193128 211006 193180 211012
rect 194140 211064 194192 211070
rect 194140 211006 194192 211012
rect 193140 210526 193168 211006
rect 193128 210520 193180 210526
rect 193128 210462 193180 210468
rect 193034 183152 193090 183161
rect 193034 183087 193090 183096
rect 191746 180024 191802 180033
rect 191746 179959 191802 179968
rect 191194 177304 191250 177313
rect 191194 177239 191250 177248
rect 193140 176633 193168 210462
rect 194796 206990 194824 211822
rect 194784 206984 194836 206990
rect 194784 206926 194836 206932
rect 193862 202192 193918 202201
rect 193862 202127 193918 202136
rect 193126 176624 193182 176633
rect 193126 176559 193182 176568
rect 191104 141500 191156 141506
rect 191104 141442 191156 141448
rect 191196 122120 191248 122126
rect 191196 122062 191248 122068
rect 191104 86284 191156 86290
rect 191104 86226 191156 86232
rect 189724 32496 189776 32502
rect 189724 32438 189776 32444
rect 188344 20052 188396 20058
rect 188344 19994 188396 20000
rect 184204 4888 184256 4894
rect 184204 4830 184256 4836
rect 173162 4040 173218 4049
rect 173162 3975 173218 3984
rect 191116 3505 191144 86226
rect 191208 60654 191236 122062
rect 191288 106412 191340 106418
rect 191288 106354 191340 106360
rect 191300 85513 191328 106354
rect 191286 85504 191342 85513
rect 191286 85439 191342 85448
rect 191196 60648 191248 60654
rect 191196 60590 191248 60596
rect 193876 43489 193904 202127
rect 193862 43480 193918 43489
rect 193862 43415 193918 43424
rect 195256 13161 195284 313239
rect 195348 283801 195376 369815
rect 198004 361684 198056 361690
rect 198004 361626 198056 361632
rect 195428 351960 195480 351966
rect 195428 351902 195480 351908
rect 195334 283792 195390 283801
rect 195334 283727 195390 283736
rect 195440 267510 195468 351902
rect 196716 346452 196768 346458
rect 196716 346394 196768 346400
rect 196624 320952 196676 320958
rect 196624 320894 196676 320900
rect 195520 285728 195572 285734
rect 195520 285670 195572 285676
rect 195428 267504 195480 267510
rect 195428 267446 195480 267452
rect 195532 262954 195560 285670
rect 195980 283960 196032 283966
rect 195980 283902 196032 283908
rect 195992 278089 196020 283902
rect 195978 278080 196034 278089
rect 195978 278015 196034 278024
rect 195888 272536 195940 272542
rect 195888 272478 195940 272484
rect 195900 271930 195928 272478
rect 195888 271924 195940 271930
rect 195888 271866 195940 271872
rect 195520 262948 195572 262954
rect 195520 262890 195572 262896
rect 195336 249960 195388 249966
rect 195336 249902 195388 249908
rect 195348 249082 195376 249902
rect 195336 249076 195388 249082
rect 195336 249018 195388 249024
rect 195334 241632 195390 241641
rect 195334 241567 195390 241576
rect 195348 230353 195376 241567
rect 195796 241528 195848 241534
rect 195796 241470 195848 241476
rect 195334 230344 195390 230353
rect 195334 230279 195390 230288
rect 195808 219502 195836 241470
rect 195900 229945 195928 271866
rect 196636 240446 196664 320894
rect 196728 314809 196756 346394
rect 196714 314800 196770 314809
rect 196714 314735 196770 314744
rect 197266 314800 197322 314809
rect 197266 314735 197322 314744
rect 197174 308408 197230 308417
rect 197174 308343 197230 308352
rect 197188 303686 197216 308343
rect 197176 303680 197228 303686
rect 197176 303622 197228 303628
rect 197280 301578 197308 314735
rect 197268 301572 197320 301578
rect 197268 301514 197320 301520
rect 198016 292505 198044 361626
rect 198096 346520 198148 346526
rect 198096 346462 198148 346468
rect 198108 330614 198136 346462
rect 198096 330608 198148 330614
rect 198096 330550 198148 330556
rect 199476 313948 199528 313954
rect 199476 313890 199528 313896
rect 199384 309256 199436 309262
rect 199384 309198 199436 309204
rect 198188 303680 198240 303686
rect 198188 303622 198240 303628
rect 198096 301572 198148 301578
rect 198096 301514 198148 301520
rect 198002 292496 198058 292505
rect 198002 292431 198058 292440
rect 198002 290184 198058 290193
rect 198002 290119 198058 290128
rect 196716 284980 196768 284986
rect 196716 284922 196768 284928
rect 196728 247353 196756 284922
rect 197358 282432 197414 282441
rect 197358 282367 197414 282376
rect 197372 281586 197400 282367
rect 197360 281580 197412 281586
rect 197360 281522 197412 281528
rect 197360 281444 197412 281450
rect 197360 281386 197412 281392
rect 197372 280809 197400 281386
rect 197358 280800 197414 280809
rect 197358 280735 197414 280744
rect 197450 280256 197506 280265
rect 197450 280191 197506 280200
rect 197360 280152 197412 280158
rect 197360 280094 197412 280100
rect 197372 279449 197400 280094
rect 197464 279478 197492 280191
rect 197452 279472 197504 279478
rect 197358 279440 197414 279449
rect 197452 279414 197504 279420
rect 197358 279375 197414 279384
rect 197358 278624 197414 278633
rect 197280 278582 197358 278610
rect 197280 278050 197308 278582
rect 197358 278559 197414 278568
rect 197268 278044 197320 278050
rect 197268 277986 197320 277992
rect 197174 249112 197230 249121
rect 197174 249047 197230 249056
rect 196714 247344 196770 247353
rect 196714 247279 196770 247288
rect 196714 243808 196770 243817
rect 196714 243743 196770 243752
rect 196624 240440 196676 240446
rect 196624 240382 196676 240388
rect 195886 229936 195942 229945
rect 195886 229871 195942 229880
rect 196728 223417 196756 243743
rect 197082 231568 197138 231577
rect 197082 231503 197138 231512
rect 197096 230625 197124 231503
rect 197082 230616 197138 230625
rect 197082 230551 197138 230560
rect 197096 228449 197124 230551
rect 197082 228440 197138 228449
rect 197082 228375 197138 228384
rect 196714 223408 196770 223417
rect 196714 223343 196770 223352
rect 195796 219496 195848 219502
rect 195796 219438 195848 219444
rect 195808 219337 195836 219438
rect 195794 219328 195850 219337
rect 195794 219263 195850 219272
rect 195334 215384 195390 215393
rect 195334 215319 195390 215328
rect 195348 203561 195376 215319
rect 195334 203552 195390 203561
rect 195334 203487 195390 203496
rect 195334 202328 195390 202337
rect 195334 202263 195390 202272
rect 195348 135930 195376 202263
rect 197188 188465 197216 249047
rect 197280 197985 197308 277986
rect 197360 277160 197412 277166
rect 197360 277102 197412 277108
rect 197372 276729 197400 277102
rect 197358 276720 197414 276729
rect 198016 276690 198044 290119
rect 198108 278089 198136 301514
rect 198200 282985 198228 303622
rect 198278 288552 198334 288561
rect 198278 288487 198334 288496
rect 198186 282976 198242 282985
rect 198186 282911 198242 282920
rect 198094 278080 198150 278089
rect 198094 278015 198150 278024
rect 197358 276655 197414 276664
rect 198004 276684 198056 276690
rect 198004 276626 198056 276632
rect 198292 276010 198320 288487
rect 198738 285832 198794 285841
rect 198738 285767 198794 285776
rect 198752 282266 198780 285767
rect 198740 282260 198792 282266
rect 198740 282202 198792 282208
rect 198280 276004 198332 276010
rect 198280 275946 198332 275952
rect 197450 275088 197506 275097
rect 197450 275023 197506 275032
rect 197464 274718 197492 275023
rect 197452 274712 197504 274718
rect 197452 274654 197504 274660
rect 197360 274644 197412 274650
rect 197360 274586 197412 274592
rect 197372 274553 197400 274586
rect 197358 274544 197414 274553
rect 197358 274479 197414 274488
rect 197358 273728 197414 273737
rect 197358 273663 197414 273672
rect 197372 273290 197400 273663
rect 197360 273284 197412 273290
rect 197360 273226 197412 273232
rect 197358 272912 197414 272921
rect 197358 272847 197414 272856
rect 197372 271930 197400 272847
rect 197360 271924 197412 271930
rect 197360 271866 197412 271872
rect 197358 271552 197414 271561
rect 197358 271487 197414 271496
rect 197372 270570 197400 271487
rect 197450 271008 197506 271017
rect 197450 270943 197506 270952
rect 197464 270638 197492 270943
rect 197452 270632 197504 270638
rect 197452 270574 197504 270580
rect 197360 270564 197412 270570
rect 197360 270506 197412 270512
rect 197358 270192 197414 270201
rect 197358 270127 197414 270136
rect 197372 269210 197400 270127
rect 197360 269204 197412 269210
rect 197360 269146 197412 269152
rect 197360 269068 197412 269074
rect 197360 269010 197412 269016
rect 197372 268841 197400 269010
rect 197358 268832 197414 268841
rect 197358 268767 197414 268776
rect 197360 267504 197412 267510
rect 197360 267446 197412 267452
rect 197372 266665 197400 267446
rect 197358 266656 197414 266665
rect 197358 266591 197414 266600
rect 197360 266348 197412 266354
rect 197360 266290 197412 266296
rect 197372 265849 197400 266290
rect 197358 265840 197414 265849
rect 197358 265775 197414 265784
rect 197360 264920 197412 264926
rect 197360 264862 197412 264868
rect 197372 264489 197400 264862
rect 197358 264480 197414 264489
rect 197358 264415 197414 264424
rect 197358 263664 197414 263673
rect 197358 263599 197360 263608
rect 197412 263599 197414 263608
rect 197360 263570 197412 263576
rect 197360 262336 197412 262342
rect 197358 262304 197360 262313
rect 197412 262304 197414 262313
rect 197358 262239 197414 262248
rect 197450 261488 197506 261497
rect 197450 261423 197506 261432
rect 197360 260976 197412 260982
rect 197358 260944 197360 260953
rect 197412 260944 197414 260953
rect 197464 260914 197492 261423
rect 197358 260879 197414 260888
rect 197452 260908 197504 260914
rect 197452 260850 197504 260856
rect 197358 260128 197414 260137
rect 197358 260063 197414 260072
rect 197372 259486 197400 260063
rect 197360 259480 197412 259486
rect 197360 259422 197412 259428
rect 197452 259412 197504 259418
rect 197452 259354 197504 259360
rect 197358 259312 197414 259321
rect 197358 259247 197414 259256
rect 197372 258534 197400 259247
rect 197464 258777 197492 259354
rect 197450 258768 197506 258777
rect 197450 258703 197506 258712
rect 197360 258528 197412 258534
rect 197360 258470 197412 258476
rect 197358 257952 197414 257961
rect 197358 257887 197414 257896
rect 197372 256766 197400 257887
rect 197360 256760 197412 256766
rect 197360 256702 197412 256708
rect 197358 256592 197414 256601
rect 197358 256527 197414 256536
rect 197372 255338 197400 256527
rect 197360 255332 197412 255338
rect 197360 255274 197412 255280
rect 198002 255232 198058 255241
rect 198002 255167 198058 255176
rect 197358 254416 197414 254425
rect 197358 254351 197414 254360
rect 197372 253978 197400 254351
rect 197360 253972 197412 253978
rect 197360 253914 197412 253920
rect 197452 253904 197504 253910
rect 197452 253846 197504 253852
rect 197464 253609 197492 253846
rect 197450 253600 197506 253609
rect 197450 253535 197506 253544
rect 197450 252240 197506 252249
rect 197450 252175 197506 252184
rect 197358 251696 197414 251705
rect 197358 251631 197414 251640
rect 197372 251258 197400 251631
rect 197464 251326 197492 252175
rect 197452 251320 197504 251326
rect 197452 251262 197504 251268
rect 197360 251252 197412 251258
rect 197360 251194 197412 251200
rect 197450 250880 197506 250889
rect 197450 250815 197506 250824
rect 197358 250064 197414 250073
rect 197358 249999 197414 250008
rect 197372 249830 197400 249999
rect 197464 249966 197492 250815
rect 197452 249960 197504 249966
rect 197452 249902 197504 249908
rect 197360 249824 197412 249830
rect 197360 249766 197412 249772
rect 197452 249756 197504 249762
rect 197452 249698 197504 249704
rect 197464 249529 197492 249698
rect 197450 249520 197506 249529
rect 197450 249455 197506 249464
rect 197358 247888 197414 247897
rect 197358 247823 197414 247832
rect 197372 247110 197400 247823
rect 197360 247104 197412 247110
rect 197360 247046 197412 247052
rect 197452 247036 197504 247042
rect 197452 246978 197504 246984
rect 197358 246528 197414 246537
rect 197358 246463 197414 246472
rect 197372 245750 197400 246463
rect 197464 245993 197492 246978
rect 197450 245984 197506 245993
rect 197450 245919 197506 245928
rect 197360 245744 197412 245750
rect 197360 245686 197412 245692
rect 197450 245168 197506 245177
rect 197450 245103 197506 245112
rect 197464 244390 197492 245103
rect 197452 244384 197504 244390
rect 197358 244352 197414 244361
rect 197452 244326 197504 244332
rect 197358 244287 197360 244296
rect 197412 244287 197414 244296
rect 197360 244258 197412 244264
rect 197910 242176 197966 242185
rect 197910 242111 197966 242120
rect 197924 241534 197952 242111
rect 197912 241528 197964 241534
rect 198016 241505 198044 255167
rect 197912 241470 197964 241476
rect 198002 241496 198058 241505
rect 198002 241431 198058 241440
rect 198740 235272 198792 235278
rect 198740 235214 198792 235220
rect 198752 234598 198780 235214
rect 198740 234592 198792 234598
rect 198740 234534 198792 234540
rect 199396 233170 199424 309198
rect 199488 302161 199516 313890
rect 199474 302152 199530 302161
rect 199474 302087 199530 302096
rect 200946 302152 201002 302161
rect 200946 302087 201002 302096
rect 200960 301073 200988 302087
rect 200946 301064 201002 301073
rect 200946 300999 201002 301008
rect 201314 301064 201370 301073
rect 201314 300999 201370 301008
rect 200580 295384 200632 295390
rect 200580 295326 200632 295332
rect 199476 294024 199528 294030
rect 199476 293966 199528 293972
rect 199488 267714 199516 293966
rect 200394 292496 200450 292505
rect 200394 292431 200450 292440
rect 200120 284436 200172 284442
rect 200120 284378 200172 284384
rect 199568 284368 199620 284374
rect 199568 284310 199620 284316
rect 199580 268394 199608 284310
rect 200132 283898 200160 284378
rect 200408 284172 200436 292431
rect 200592 290465 200620 295326
rect 201130 292496 201186 292505
rect 201130 292431 201186 292440
rect 201144 291825 201172 292431
rect 201130 291816 201186 291825
rect 201130 291751 201186 291760
rect 200578 290456 200634 290465
rect 200578 290391 200634 290400
rect 200764 286340 200816 286346
rect 200764 286282 200816 286288
rect 200776 284172 200804 286282
rect 201328 284172 201356 300999
rect 201512 285326 201540 372642
rect 202156 352782 202184 445975
rect 582392 432614 582420 484599
rect 582654 471472 582710 471481
rect 582654 471407 582710 471416
rect 582470 458144 582526 458153
rect 582470 458079 582526 458088
rect 582484 451246 582512 458079
rect 582472 451240 582524 451246
rect 582472 451182 582524 451188
rect 582380 432608 582432 432614
rect 582380 432550 582432 432556
rect 582378 431624 582434 431633
rect 582378 431559 582434 431568
rect 582392 403646 582420 431559
rect 582380 403640 582432 403646
rect 582380 403582 582432 403588
rect 228364 376780 228416 376786
rect 228364 376722 228416 376728
rect 221462 367160 221518 367169
rect 221462 367095 221518 367104
rect 212908 365016 212960 365022
rect 212908 364958 212960 364964
rect 207664 357468 207716 357474
rect 207664 357410 207716 357416
rect 206282 353696 206338 353705
rect 206282 353631 206338 353640
rect 202144 352776 202196 352782
rect 202144 352718 202196 352724
rect 202788 352776 202840 352782
rect 202788 352718 202840 352724
rect 202800 352578 202828 352718
rect 204902 352608 204958 352617
rect 202788 352572 202840 352578
rect 204902 352543 204958 352552
rect 202788 352514 202840 352520
rect 202142 327176 202198 327185
rect 202142 327111 202198 327120
rect 202156 306374 202184 327111
rect 201696 306346 202184 306374
rect 201696 303657 201724 306346
rect 201682 303648 201738 303657
rect 201682 303583 201738 303592
rect 201500 285320 201552 285326
rect 201500 285262 201552 285268
rect 201696 284172 201724 303583
rect 202800 293282 202828 352514
rect 204258 342408 204314 342417
rect 204258 342343 204314 342352
rect 203524 335436 203576 335442
rect 203524 335378 203576 335384
rect 202788 293276 202840 293282
rect 202788 293218 202840 293224
rect 203536 292777 203564 335378
rect 203616 324964 203668 324970
rect 203616 324906 203668 324912
rect 203628 306374 203656 324906
rect 203628 306346 203748 306374
rect 203720 295458 203748 306346
rect 203708 295452 203760 295458
rect 203708 295394 203760 295400
rect 203522 292768 203578 292777
rect 203522 292703 203578 292712
rect 202142 289912 202198 289921
rect 202142 289847 202198 289856
rect 202156 284186 202184 289847
rect 203156 285728 203208 285734
rect 203156 285670 203208 285676
rect 202420 285320 202472 285326
rect 202420 285262 202472 285268
rect 202432 284186 202460 285262
rect 202156 284158 202262 284186
rect 202432 284158 202814 284186
rect 203168 284172 203196 285670
rect 203720 284172 203748 295394
rect 204166 292768 204222 292777
rect 204166 292703 204222 292712
rect 204180 285734 204208 292703
rect 204168 285728 204220 285734
rect 204272 285705 204300 342343
rect 204352 294636 204404 294642
rect 204352 294578 204404 294584
rect 204364 291650 204392 294578
rect 204352 291644 204404 291650
rect 204352 291586 204404 291592
rect 204916 285734 204944 352543
rect 204996 322992 205048 322998
rect 204996 322934 205048 322940
rect 205008 310486 205036 322934
rect 204996 310480 205048 310486
rect 204996 310422 205048 310428
rect 206296 302297 206324 353631
rect 207676 331906 207704 357410
rect 210422 348392 210478 348401
rect 210422 348327 210478 348336
rect 209042 334248 209098 334257
rect 209042 334183 209098 334192
rect 207664 331900 207716 331906
rect 207664 331842 207716 331848
rect 207754 331256 207810 331265
rect 207754 331191 207810 331200
rect 206376 319524 206428 319530
rect 206376 319466 206428 319472
rect 206388 309097 206416 319466
rect 206374 309088 206430 309097
rect 206374 309023 206430 309032
rect 206926 309088 206982 309097
rect 206926 309023 206982 309032
rect 206940 307873 206968 309023
rect 206926 307864 206982 307873
rect 206926 307799 206982 307808
rect 206282 302288 206338 302297
rect 206282 302223 206338 302232
rect 206650 302288 206706 302297
rect 206650 302223 206706 302232
rect 205548 285796 205600 285802
rect 205548 285738 205600 285744
rect 204904 285728 204956 285734
rect 204168 285670 204220 285676
rect 204258 285696 204314 285705
rect 204904 285670 204956 285676
rect 205178 285696 205234 285705
rect 204258 285631 204314 285640
rect 205178 285631 205234 285640
rect 204258 284608 204314 284617
rect 204258 284543 204314 284552
rect 204272 284172 204300 284543
rect 201958 284064 202014 284073
rect 202156 284050 202184 284158
rect 202014 284022 202184 284050
rect 201958 283999 202014 284008
rect 204352 283960 204404 283966
rect 205192 283914 205220 285631
rect 205560 284172 205588 285738
rect 206098 284336 206154 284345
rect 206098 284271 206154 284280
rect 206112 284172 206140 284271
rect 206664 284172 206692 302223
rect 206940 287054 206968 307799
rect 207768 306474 207796 331191
rect 208492 318844 208544 318850
rect 208492 318786 208544 318792
rect 207756 306468 207808 306474
rect 207756 306410 207808 306416
rect 207768 296714 207796 306410
rect 207584 296686 207796 296714
rect 206940 287026 207060 287054
rect 207032 284172 207060 287026
rect 207584 284172 207612 296686
rect 208400 288516 208452 288522
rect 208400 288458 208452 288464
rect 208412 287706 208440 288458
rect 208400 287700 208452 287706
rect 208400 287642 208452 287648
rect 208400 287564 208452 287570
rect 208400 287506 208452 287512
rect 208124 285728 208176 285734
rect 208124 285670 208176 285676
rect 208136 284172 208164 285670
rect 208412 285326 208440 287506
rect 208400 285320 208452 285326
rect 208400 285262 208452 285268
rect 208504 284172 208532 318786
rect 209056 309233 209084 334183
rect 209134 332616 209190 332625
rect 209134 332551 209190 332560
rect 209148 318850 209176 332551
rect 209136 318844 209188 318850
rect 209136 318786 209188 318792
rect 209964 310480 210016 310486
rect 209964 310422 210016 310428
rect 209976 309369 210004 310422
rect 209962 309360 210018 309369
rect 209962 309295 210018 309304
rect 209042 309224 209098 309233
rect 209042 309159 209098 309168
rect 209410 309224 209466 309233
rect 209410 309159 209466 309168
rect 208584 291644 208636 291650
rect 208584 291586 208636 291592
rect 208596 287570 208624 291586
rect 208584 287564 208636 287570
rect 208584 287506 208636 287512
rect 208676 285320 208728 285326
rect 208676 285262 208728 285268
rect 208688 284186 208716 285262
rect 208688 284158 209070 284186
rect 209424 284172 209452 309159
rect 210436 305017 210464 348327
rect 211158 331392 211214 331401
rect 211158 331327 211214 331336
rect 210514 309360 210570 309369
rect 210514 309295 210570 309304
rect 210422 305008 210478 305017
rect 210422 304943 210478 304952
rect 209964 293276 210016 293282
rect 209964 293218 210016 293224
rect 209976 284172 210004 293218
rect 210528 284172 210556 309295
rect 210882 290048 210938 290057
rect 210882 289983 210938 289992
rect 210896 287094 210924 289983
rect 210884 287088 210936 287094
rect 210884 287030 210936 287036
rect 210896 284172 210924 287030
rect 205362 283928 205418 283937
rect 204404 283908 204654 283914
rect 204352 283902 204654 283908
rect 200120 283892 200172 283898
rect 204364 283886 204654 283902
rect 205192 283900 205362 283914
rect 205206 283886 205362 283900
rect 211172 283914 211200 331327
rect 211802 329216 211858 329225
rect 211802 329151 211858 329160
rect 211816 284889 211844 329151
rect 211986 293992 212042 294001
rect 211986 293927 212042 293936
rect 212000 292913 212028 293927
rect 211986 292904 212042 292913
rect 211986 292839 212042 292848
rect 211802 284880 211858 284889
rect 211802 284815 211858 284824
rect 212000 284172 212028 292839
rect 212354 284880 212410 284889
rect 212354 284815 212410 284824
rect 212368 284172 212396 284815
rect 212920 284172 212948 364958
rect 215942 363080 215998 363089
rect 215942 363015 215998 363024
rect 214564 360256 214616 360262
rect 214564 360198 214616 360204
rect 213828 330540 213880 330546
rect 213828 330482 213880 330488
rect 213458 289096 213514 289105
rect 213458 289031 213514 289040
rect 213472 284172 213500 289031
rect 213840 284172 213868 330482
rect 214576 298858 214604 360198
rect 215390 336832 215446 336841
rect 215390 336767 215446 336776
rect 214746 305008 214802 305017
rect 214746 304943 214802 304952
rect 214564 298852 214616 298858
rect 214564 298794 214616 298800
rect 214760 284172 214788 304943
rect 215300 300960 215352 300966
rect 215300 300902 215352 300908
rect 215312 284172 215340 300902
rect 215404 284050 215432 336767
rect 215956 313993 215984 363015
rect 220082 338328 220138 338337
rect 220082 338263 220138 338272
rect 216036 338156 216088 338162
rect 216036 338098 216088 338104
rect 215942 313984 215998 313993
rect 215942 313919 215998 313928
rect 215944 303748 215996 303754
rect 215944 303690 215996 303696
rect 215956 293350 215984 303690
rect 216048 300966 216076 338098
rect 218702 336968 218758 336977
rect 218702 336903 218758 336912
rect 218716 320210 218744 336903
rect 218704 320204 218756 320210
rect 218704 320146 218756 320152
rect 219348 320204 219400 320210
rect 219348 320146 219400 320152
rect 218704 311908 218756 311914
rect 218704 311850 218756 311856
rect 216036 300960 216088 300966
rect 216036 300902 216088 300908
rect 216588 298784 216640 298790
rect 216588 298726 216640 298732
rect 216600 294710 216628 298726
rect 216680 295384 216732 295390
rect 216680 295326 216732 295332
rect 216588 294704 216640 294710
rect 216588 294646 216640 294652
rect 216692 294001 216720 295326
rect 218716 294642 218744 311850
rect 218704 294636 218756 294642
rect 218704 294578 218756 294584
rect 218060 294024 218112 294030
rect 216678 293992 216734 294001
rect 216678 293927 216734 293936
rect 217690 293992 217746 294001
rect 218060 293966 218112 293972
rect 217690 293927 217746 293936
rect 215944 293344 215996 293350
rect 215944 293286 215996 293292
rect 215484 292596 215536 292602
rect 215484 292538 215536 292544
rect 215496 288386 215524 292538
rect 215484 288380 215536 288386
rect 215484 288322 215536 288328
rect 216680 284980 216732 284986
rect 216680 284922 216732 284928
rect 216692 284889 216720 284922
rect 216678 284880 216734 284889
rect 216678 284815 216734 284824
rect 216772 284776 216824 284782
rect 216772 284718 216824 284724
rect 216784 284442 216812 284718
rect 216772 284436 216824 284442
rect 216772 284378 216824 284384
rect 216784 284172 216812 284378
rect 217324 284368 217376 284374
rect 217324 284310 217376 284316
rect 217336 284172 217364 284310
rect 217704 284172 217732 293927
rect 218072 291854 218100 293966
rect 218610 292632 218666 292641
rect 218610 292567 218666 292576
rect 218060 291848 218112 291854
rect 218060 291790 218112 291796
rect 218060 288516 218112 288522
rect 218060 288458 218112 288464
rect 218072 288386 218100 288458
rect 218060 288380 218112 288386
rect 218060 288322 218112 288328
rect 218242 286376 218298 286385
rect 218242 286311 218298 286320
rect 218256 284172 218284 286311
rect 218624 284172 218652 292567
rect 218704 286340 218756 286346
rect 218704 286282 218756 286288
rect 218716 285841 218744 286282
rect 219360 285938 219388 320146
rect 219716 318436 219768 318442
rect 219716 318378 219768 318384
rect 219728 317490 219756 318378
rect 219716 317484 219768 317490
rect 219716 317426 219768 317432
rect 219440 287088 219492 287094
rect 219440 287030 219492 287036
rect 219348 285932 219400 285938
rect 219348 285874 219400 285880
rect 218702 285832 218758 285841
rect 218702 285767 218758 285776
rect 218716 284186 218744 285767
rect 219452 284782 219480 287030
rect 219440 284776 219492 284782
rect 219440 284718 219492 284724
rect 218716 284158 219190 284186
rect 219728 284172 219756 317426
rect 220096 311914 220124 338263
rect 220176 334008 220228 334014
rect 220176 333950 220228 333956
rect 220188 318442 220216 333950
rect 220176 318436 220228 318442
rect 220176 318378 220228 318384
rect 220084 311908 220136 311914
rect 220084 311850 220136 311856
rect 220728 311908 220780 311914
rect 220728 311850 220780 311856
rect 220636 288516 220688 288522
rect 220636 288458 220688 288464
rect 220082 284336 220138 284345
rect 220082 284271 220138 284280
rect 220096 284172 220124 284271
rect 220648 284172 220676 288458
rect 220740 285705 220768 311850
rect 221188 285932 221240 285938
rect 221188 285874 221240 285880
rect 220726 285696 220782 285705
rect 220726 285631 220782 285640
rect 221200 284172 221228 285874
rect 221476 285841 221504 367095
rect 224224 358828 224276 358834
rect 224224 358770 224276 358776
rect 222844 349852 222896 349858
rect 222844 349794 222896 349800
rect 221554 334384 221610 334393
rect 221554 334319 221610 334328
rect 221568 310593 221596 334319
rect 221554 310584 221610 310593
rect 221554 310519 221610 310528
rect 221462 285832 221518 285841
rect 221462 285767 221518 285776
rect 221568 284172 221596 310519
rect 222856 291961 222884 349794
rect 222936 347812 222988 347818
rect 222936 347754 222988 347760
rect 222948 296857 222976 347754
rect 222934 296848 222990 296857
rect 222934 296783 222990 296792
rect 222842 291952 222898 291961
rect 222842 291887 222898 291896
rect 222948 287054 222976 296783
rect 223028 291236 223080 291242
rect 223028 291178 223080 291184
rect 223580 291236 223632 291242
rect 223580 291178 223632 291184
rect 222856 287026 222976 287054
rect 222106 285696 222162 285705
rect 222106 285631 222162 285640
rect 222120 284172 222148 285631
rect 222856 284186 222884 287026
rect 222502 284158 222884 284186
rect 223040 284172 223068 291178
rect 223592 288454 223620 291178
rect 223580 288448 223632 288454
rect 223580 288390 223632 288396
rect 223592 284172 223620 288390
rect 223946 285696 224002 285705
rect 223946 285631 224002 285640
rect 223960 284172 223988 285631
rect 224236 284345 224264 358770
rect 224316 345092 224368 345098
rect 224316 345034 224368 345040
rect 224328 304298 224356 345034
rect 226430 342544 226486 342553
rect 226430 342479 226486 342488
rect 225604 341012 225656 341018
rect 225604 340954 225656 340960
rect 225418 327448 225474 327457
rect 225418 327383 225474 327392
rect 224868 318096 224920 318102
rect 224868 318038 224920 318044
rect 224880 314702 224908 318038
rect 224868 314696 224920 314702
rect 224868 314638 224920 314644
rect 224316 304292 224368 304298
rect 224316 304234 224368 304240
rect 224684 287700 224736 287706
rect 224684 287642 224736 287648
rect 224696 287162 224724 287642
rect 224684 287156 224736 287162
rect 224684 287098 224736 287104
rect 224222 284336 224278 284345
rect 224222 284271 224278 284280
rect 224696 284186 224724 287098
rect 224880 287054 224908 314638
rect 224880 287026 225000 287054
rect 224526 284158 224724 284186
rect 224972 284186 225000 287026
rect 224972 284158 225078 284186
rect 225432 284172 225460 327383
rect 225616 299713 225644 340954
rect 226340 313404 226392 313410
rect 226340 313346 226392 313352
rect 226352 309126 226380 313346
rect 226340 309120 226392 309126
rect 226340 309062 226392 309068
rect 225602 299704 225658 299713
rect 225602 299639 225658 299648
rect 225970 297528 226026 297537
rect 225970 297463 226026 297472
rect 225984 284172 226012 297463
rect 216034 284064 216090 284073
rect 215404 284022 216034 284050
rect 216034 283999 216090 284008
rect 211618 283928 211674 283937
rect 211172 283886 211618 283914
rect 205362 283863 205418 283872
rect 214470 283928 214526 283937
rect 214406 283886 214470 283914
rect 211618 283863 211674 283872
rect 214470 283863 214526 283872
rect 215942 283928 215998 283937
rect 226444 283914 226472 342479
rect 226982 332752 227038 332761
rect 226982 332687 227038 332696
rect 226996 284345 227024 332687
rect 227810 299704 227866 299713
rect 227810 299639 227866 299648
rect 227444 298852 227496 298858
rect 227444 298794 227496 298800
rect 226982 284336 227038 284345
rect 226982 284271 227038 284280
rect 226996 284186 227024 284271
rect 226918 284158 227024 284186
rect 227456 284172 227484 298794
rect 227824 284172 227852 299639
rect 228376 298489 228404 376722
rect 331220 372632 331272 372638
rect 331220 372574 331272 372580
rect 232504 371340 232556 371346
rect 232504 371282 232556 371288
rect 231124 368552 231176 368558
rect 231124 368494 231176 368500
rect 230480 354748 230532 354754
rect 230480 354690 230532 354696
rect 228454 335472 228510 335481
rect 228454 335407 228510 335416
rect 228468 307834 228496 335407
rect 230386 330440 230442 330449
rect 230386 330375 230442 330384
rect 230020 311228 230072 311234
rect 230020 311170 230072 311176
rect 230032 310729 230060 311170
rect 230018 310720 230074 310729
rect 230018 310655 230074 310664
rect 228456 307828 228508 307834
rect 228456 307770 228508 307776
rect 228916 307828 228968 307834
rect 228916 307770 228968 307776
rect 228362 298480 228418 298489
rect 228362 298415 228418 298424
rect 228364 294704 228416 294710
rect 228364 294646 228416 294652
rect 228376 284172 228404 294646
rect 228928 284172 228956 307770
rect 229006 298480 229062 298489
rect 229006 298415 229062 298424
rect 229020 285682 229048 298415
rect 230032 296714 230060 310655
rect 229848 296686 230060 296714
rect 229020 285654 229140 285682
rect 229112 284186 229140 285654
rect 229112 284158 229310 284186
rect 229848 284172 229876 296686
rect 230400 284172 230428 330375
rect 230492 284481 230520 354690
rect 231136 299470 231164 368494
rect 231124 299464 231176 299470
rect 231124 299406 231176 299412
rect 231122 290184 231178 290193
rect 231122 290119 231178 290128
rect 230478 284472 230534 284481
rect 231136 284442 231164 290119
rect 231306 287192 231362 287201
rect 231306 287127 231362 287136
rect 230478 284407 230534 284416
rect 230756 284436 230808 284442
rect 230756 284378 230808 284384
rect 231124 284436 231176 284442
rect 231124 284378 231176 284384
rect 230768 284172 230796 284378
rect 231320 284172 231348 287127
rect 232516 285841 232544 371282
rect 240508 371272 240560 371278
rect 240508 371214 240560 371220
rect 233882 357504 233938 357513
rect 233882 357439 233938 357448
rect 232594 323640 232650 323649
rect 232594 323575 232650 323584
rect 232502 285832 232558 285841
rect 232502 285767 232558 285776
rect 231674 284472 231730 284481
rect 231674 284407 231730 284416
rect 231688 284172 231716 284407
rect 232516 284186 232544 285767
rect 232608 285734 232636 323575
rect 233148 299464 233200 299470
rect 233148 299406 233200 299412
rect 233160 298178 233188 299406
rect 233148 298172 233200 298178
rect 233148 298114 233200 298120
rect 232596 285728 232648 285734
rect 232596 285670 232648 285676
rect 232778 284744 232834 284753
rect 232778 284679 232834 284688
rect 232254 284158 232544 284186
rect 232792 284172 232820 284679
rect 233160 284172 233188 298114
rect 233896 289814 233924 357439
rect 238024 356108 238076 356114
rect 238024 356050 238076 356056
rect 234618 353424 234674 353433
rect 234618 353359 234674 353368
rect 233974 328672 234030 328681
rect 233974 328607 234030 328616
rect 233988 295390 234016 328607
rect 233976 295384 234028 295390
rect 233976 295326 234028 295332
rect 233884 289808 233936 289814
rect 233884 289750 233936 289756
rect 233988 284186 234016 295326
rect 234252 285728 234304 285734
rect 234252 285670 234304 285676
rect 233726 284158 234016 284186
rect 234264 284172 234292 285670
rect 234632 284172 234660 353359
rect 236644 320884 236696 320890
rect 236644 320826 236696 320832
rect 236000 311160 236052 311166
rect 236000 311102 236052 311108
rect 235172 293276 235224 293282
rect 235172 293218 235224 293224
rect 235184 284172 235212 293218
rect 235540 289808 235592 289814
rect 235540 289750 235592 289756
rect 235552 284172 235580 289750
rect 226798 283928 226854 283937
rect 215998 283886 216246 283914
rect 226444 283886 226798 283914
rect 215942 283863 215998 283872
rect 236012 283914 236040 311102
rect 236656 299577 236684 320826
rect 238036 312497 238064 356050
rect 239404 331900 239456 331906
rect 239404 331842 239456 331848
rect 238206 327312 238262 327321
rect 238206 327247 238262 327256
rect 238116 319456 238168 319462
rect 238116 319398 238168 319404
rect 238022 312488 238078 312497
rect 238022 312423 238078 312432
rect 236826 299840 236882 299849
rect 236826 299775 236882 299784
rect 236642 299568 236698 299577
rect 236642 299503 236698 299512
rect 236458 287328 236514 287337
rect 236458 287263 236514 287272
rect 236472 286346 236500 287263
rect 236460 286340 236512 286346
rect 236460 286282 236512 286288
rect 236656 284172 236684 299503
rect 236736 293344 236788 293350
rect 236736 293286 236788 293292
rect 236748 288454 236776 293286
rect 236840 293185 236868 299775
rect 238128 296714 238156 319398
rect 238220 298110 238248 327247
rect 239220 312588 239272 312594
rect 239220 312530 239272 312536
rect 239232 307766 239260 312530
rect 239220 307760 239272 307766
rect 239220 307702 239272 307708
rect 239416 302433 239444 331842
rect 239496 306400 239548 306406
rect 239496 306342 239548 306348
rect 239402 302424 239458 302433
rect 239402 302359 239458 302368
rect 238208 298104 238260 298110
rect 238208 298046 238260 298052
rect 238668 298104 238720 298110
rect 238668 298046 238720 298052
rect 238680 296750 238708 298046
rect 237944 296686 238156 296714
rect 238668 296744 238720 296750
rect 238668 296686 238720 296692
rect 236826 293176 236882 293185
rect 236826 293111 236882 293120
rect 236736 288448 236788 288454
rect 236736 288390 236788 288396
rect 236748 284186 236776 288390
rect 237944 285734 237972 296686
rect 238574 290184 238630 290193
rect 238574 290119 238630 290128
rect 238114 287600 238170 287609
rect 238114 287535 238170 287544
rect 237564 285728 237616 285734
rect 237564 285670 237616 285676
rect 237932 285728 237984 285734
rect 237932 285670 237984 285676
rect 236748 284158 237038 284186
rect 237576 284172 237604 285670
rect 238128 284617 238156 287535
rect 238114 284608 238170 284617
rect 238114 284543 238170 284552
rect 238128 284172 238156 284543
rect 238588 284186 238616 290119
rect 238680 285682 238708 296686
rect 239508 288425 239536 306342
rect 239586 302424 239642 302433
rect 239586 302359 239642 302368
rect 239494 288416 239550 288425
rect 239494 288351 239550 288360
rect 238680 285654 238800 285682
rect 238510 284158 238616 284186
rect 238772 284186 238800 285654
rect 238772 284158 239062 284186
rect 239600 284172 239628 302359
rect 239954 291272 240010 291281
rect 239954 291207 240010 291216
rect 239968 284172 239996 291207
rect 240048 284980 240100 284986
rect 240048 284922 240100 284928
rect 240060 284345 240088 284922
rect 240046 284336 240102 284345
rect 240046 284271 240102 284280
rect 240520 284172 240548 371214
rect 327078 368520 327134 368529
rect 327078 368455 327134 368464
rect 251272 367124 251324 367130
rect 251272 367066 251324 367072
rect 243176 365764 243228 365770
rect 243176 365706 243228 365712
rect 241520 361616 241572 361622
rect 241520 361558 241572 361564
rect 240782 313984 240838 313993
rect 240782 313919 240838 313928
rect 240796 306374 240824 313919
rect 240796 306346 240916 306374
rect 240888 294030 240916 306346
rect 241426 295488 241482 295497
rect 241426 295423 241482 295432
rect 240876 294024 240928 294030
rect 240876 293966 240928 293972
rect 240888 284172 240916 293966
rect 241440 284172 241468 295423
rect 241532 293282 241560 361558
rect 242164 326392 242216 326398
rect 242164 326334 242216 326340
rect 243082 326360 243138 326369
rect 241520 293276 241572 293282
rect 241520 293218 241572 293224
rect 241980 284368 242032 284374
rect 241980 284310 242032 284316
rect 241992 284186 242020 284310
rect 242176 284186 242204 326334
rect 243082 326295 243138 326304
rect 242256 316736 242308 316742
rect 242256 316678 242308 316684
rect 242268 306374 242296 316678
rect 242532 307760 242584 307766
rect 242532 307702 242584 307708
rect 242544 306374 242572 307702
rect 242268 306346 242388 306374
rect 242544 306346 242848 306374
rect 242360 285977 242388 306346
rect 242820 287054 242848 306346
rect 242820 287026 242940 287054
rect 242346 285968 242402 285977
rect 242346 285903 242402 285912
rect 241992 284172 242204 284186
rect 242360 284172 242388 285903
rect 242912 284172 242940 287026
rect 242006 284158 242204 284172
rect 243096 284050 243124 326295
rect 243188 284209 243216 365706
rect 251180 362976 251232 362982
rect 251180 362918 251232 362924
rect 249800 349172 249852 349178
rect 249800 349114 249852 349120
rect 246304 343664 246356 343670
rect 246304 343606 246356 343612
rect 244280 339516 244332 339522
rect 244280 339458 244332 339464
rect 243912 302252 243964 302258
rect 243912 302194 243964 302200
rect 243818 288416 243874 288425
rect 243818 288351 243874 288360
rect 243174 284200 243230 284209
rect 243832 284172 243860 288351
rect 243924 287054 243952 302194
rect 243924 287026 244044 287054
rect 243912 284436 243964 284442
rect 243912 284378 243964 284384
rect 243174 284135 243230 284144
rect 243634 284064 243690 284073
rect 243096 284022 243634 284050
rect 243634 283999 243690 284008
rect 236274 283928 236330 283937
rect 236012 283886 236274 283914
rect 226798 283863 226854 283872
rect 243924 283898 243952 284378
rect 236274 283863 236330 283872
rect 243912 283892 243964 283898
rect 200120 283834 200172 283840
rect 243912 283834 243964 283840
rect 244016 276162 244044 287026
rect 244292 283257 244320 339458
rect 246028 315308 246080 315314
rect 246028 315250 246080 315256
rect 245752 305652 245804 305658
rect 245752 305594 245804 305600
rect 244464 299600 244516 299606
rect 244464 299542 244516 299548
rect 244372 291848 244424 291854
rect 244372 291790 244424 291796
rect 244278 283248 244334 283257
rect 244278 283183 244334 283192
rect 244016 276146 244320 276162
rect 244016 276140 244332 276146
rect 244016 276134 244280 276140
rect 244280 276082 244332 276088
rect 199660 269136 199712 269142
rect 199660 269078 199712 269084
rect 199568 268388 199620 268394
rect 199568 268330 199620 268336
rect 199476 267708 199528 267714
rect 199476 267650 199528 267656
rect 199474 263120 199530 263129
rect 199474 263055 199530 263064
rect 199488 245857 199516 263055
rect 199672 257417 199700 269078
rect 199658 257408 199714 257417
rect 199658 257343 199714 257352
rect 199934 257408 199990 257417
rect 199934 257343 199990 257352
rect 199948 248414 199976 257343
rect 200026 253056 200082 253065
rect 200026 252991 200082 253000
rect 200040 248577 200068 252991
rect 244384 250345 244412 291790
rect 244476 268841 244504 299542
rect 244556 289876 244608 289882
rect 244556 289818 244608 289824
rect 244462 268832 244518 268841
rect 244462 268767 244518 268776
rect 244476 267782 244504 268767
rect 244464 267776 244516 267782
rect 244464 267718 244516 267724
rect 244568 260953 244596 289818
rect 245382 283248 245438 283257
rect 245382 283183 245438 283192
rect 245396 282946 245424 283183
rect 245384 282940 245436 282946
rect 245384 282882 245436 282888
rect 245658 282432 245714 282441
rect 245658 282367 245714 282376
rect 245672 281586 245700 282367
rect 245660 281580 245712 281586
rect 245660 281522 245712 281528
rect 245658 281072 245714 281081
rect 245658 281007 245714 281016
rect 245672 280226 245700 281007
rect 245660 280220 245712 280226
rect 245660 280162 245712 280168
rect 244646 278896 244702 278905
rect 244646 278831 244702 278840
rect 244554 260944 244610 260953
rect 244554 260879 244610 260888
rect 244462 256048 244518 256057
rect 244462 255983 244518 255992
rect 244370 250336 244426 250345
rect 244200 250294 244370 250322
rect 200026 248568 200082 248577
rect 200026 248503 200082 248512
rect 199948 248386 200068 248414
rect 199474 245848 199530 245857
rect 199474 245783 199530 245792
rect 199384 233164 199436 233170
rect 199384 233106 199436 233112
rect 198096 219496 198148 219502
rect 198096 219438 198148 219444
rect 198002 216744 198058 216753
rect 198002 216679 198058 216688
rect 197266 197976 197322 197985
rect 197266 197911 197322 197920
rect 197174 188456 197230 188465
rect 197174 188391 197230 188400
rect 198016 145654 198044 216679
rect 198108 172417 198136 219438
rect 199488 202201 199516 245783
rect 199842 244624 199898 244633
rect 199842 244559 199898 244568
rect 199568 243568 199620 243574
rect 199568 243510 199620 243516
rect 199580 235958 199608 243510
rect 199856 240145 199884 244559
rect 199936 240508 199988 240514
rect 199936 240450 199988 240456
rect 199948 240417 199976 240450
rect 199934 240408 199990 240417
rect 199934 240343 199990 240352
rect 199842 240136 199898 240145
rect 199842 240071 199898 240080
rect 199568 235952 199620 235958
rect 199568 235894 199620 235900
rect 200040 220114 200068 248386
rect 244200 242298 244228 250294
rect 244370 250271 244426 250280
rect 244370 247344 244426 247353
rect 244370 247279 244426 247288
rect 244200 242270 244320 242298
rect 244292 242214 244320 242270
rect 244280 242208 244332 242214
rect 244280 242150 244332 242156
rect 244002 241360 244058 241369
rect 244002 241295 244058 241304
rect 200120 240780 200172 240786
rect 200120 240722 200172 240728
rect 200132 240378 200160 240722
rect 200120 240372 200172 240378
rect 200120 240314 200172 240320
rect 200118 240272 200174 240281
rect 200118 240207 200174 240216
rect 200132 233866 200160 240207
rect 200224 238649 200252 240244
rect 200304 240168 200356 240174
rect 200592 240145 200620 240244
rect 201040 240168 201092 240174
rect 200304 240110 200356 240116
rect 200578 240136 200634 240145
rect 200210 238640 200266 238649
rect 200210 238575 200266 238584
rect 200224 235498 200252 238575
rect 200316 237969 200344 240110
rect 201144 240122 201172 240244
rect 201092 240116 201172 240122
rect 201040 240110 201172 240116
rect 201408 240168 201460 240174
rect 201512 240122 201540 240244
rect 201460 240116 201540 240122
rect 201408 240110 201540 240116
rect 201052 240094 201172 240110
rect 201420 240094 201540 240110
rect 200578 240071 200634 240080
rect 200302 237960 200358 237969
rect 200302 237895 200358 237904
rect 200592 237425 200620 240071
rect 201144 238754 201172 240094
rect 201144 238726 201356 238754
rect 200578 237416 200634 237425
rect 200578 237351 200634 237360
rect 200224 235470 200344 235498
rect 200132 233838 200252 233866
rect 200120 229764 200172 229770
rect 200120 229706 200172 229712
rect 200132 228993 200160 229706
rect 200118 228984 200174 228993
rect 200118 228919 200174 228928
rect 200224 227769 200252 233838
rect 200316 230450 200344 235470
rect 200304 230444 200356 230450
rect 200304 230386 200356 230392
rect 200210 227760 200266 227769
rect 200210 227695 200266 227704
rect 200854 227760 200910 227769
rect 200854 227695 200910 227704
rect 200028 220108 200080 220114
rect 200028 220050 200080 220056
rect 200762 215928 200818 215937
rect 200762 215863 200818 215872
rect 199474 202192 199530 202201
rect 199474 202127 199530 202136
rect 200776 197334 200804 215863
rect 200868 210361 200896 227695
rect 200854 210352 200910 210361
rect 200854 210287 200910 210296
rect 201328 202230 201356 238726
rect 201406 237416 201462 237425
rect 201406 237351 201462 237360
rect 201316 202224 201368 202230
rect 201316 202166 201368 202172
rect 200764 197328 200816 197334
rect 200764 197270 200816 197276
rect 201420 196722 201448 237351
rect 201408 196716 201460 196722
rect 201408 196658 201460 196664
rect 201512 192506 201540 240094
rect 202064 238649 202092 240244
rect 202616 238754 202644 240244
rect 202248 238726 202644 238754
rect 202050 238640 202106 238649
rect 202050 238575 202106 238584
rect 202248 238513 202276 238726
rect 202234 238504 202290 238513
rect 202234 238439 202290 238448
rect 202144 230444 202196 230450
rect 202144 230386 202196 230392
rect 201500 192500 201552 192506
rect 201500 192442 201552 192448
rect 202156 187066 202184 230386
rect 202248 213353 202276 238439
rect 202234 213344 202290 213353
rect 202234 213279 202290 213288
rect 202984 205601 203012 240244
rect 203536 238754 203564 240244
rect 203168 238726 203564 238754
rect 204088 238754 204116 240244
rect 204088 238726 204208 238754
rect 203168 212401 203196 238726
rect 204180 234530 204208 238726
rect 204456 237289 204484 240244
rect 204442 237280 204498 237289
rect 204442 237215 204498 237224
rect 204168 234524 204220 234530
rect 204168 234466 204220 234472
rect 204180 233918 204208 234466
rect 204168 233912 204220 233918
rect 203522 233880 203578 233889
rect 204168 233854 204220 233860
rect 203522 233815 203578 233824
rect 203536 219337 203564 233815
rect 205008 226137 205036 240244
rect 204994 226128 205050 226137
rect 204994 226063 205050 226072
rect 205008 224262 205036 226063
rect 204996 224256 205048 224262
rect 204996 224198 205048 224204
rect 205086 224224 205142 224233
rect 205086 224159 205142 224168
rect 203522 219328 203578 219337
rect 203522 219263 203578 219272
rect 204996 215960 205048 215966
rect 204996 215902 205048 215908
rect 204902 215384 204958 215393
rect 204902 215319 204958 215328
rect 203154 212392 203210 212401
rect 203154 212327 203210 212336
rect 203168 209774 203196 212327
rect 203168 209746 203564 209774
rect 202970 205592 203026 205601
rect 202970 205527 203026 205536
rect 203536 199510 203564 209746
rect 203614 205592 203670 205601
rect 203614 205527 203670 205536
rect 203524 199504 203576 199510
rect 203524 199446 203576 199452
rect 202328 192568 202380 192574
rect 202328 192510 202380 192516
rect 202144 187060 202196 187066
rect 202144 187002 202196 187008
rect 202234 186960 202290 186969
rect 202234 186895 202290 186904
rect 198094 172408 198150 172417
rect 198094 172343 198150 172352
rect 198004 145648 198056 145654
rect 198004 145590 198056 145596
rect 196716 143608 196768 143614
rect 196716 143550 196768 143556
rect 195336 135924 195388 135930
rect 195336 135866 195388 135872
rect 195336 128376 195388 128382
rect 195336 128318 195388 128324
rect 195348 57934 195376 128318
rect 196624 126336 196676 126342
rect 196624 126278 196676 126284
rect 195336 57928 195388 57934
rect 195336 57870 195388 57876
rect 196636 31142 196664 126278
rect 196728 90370 196756 143550
rect 199384 141432 199436 141438
rect 199384 141374 199436 141380
rect 198096 138712 198148 138718
rect 198096 138654 198148 138660
rect 198004 134564 198056 134570
rect 198004 134506 198056 134512
rect 196716 90364 196768 90370
rect 196716 90306 196768 90312
rect 196716 89004 196768 89010
rect 196716 88946 196768 88952
rect 196624 31136 196676 31142
rect 196624 31078 196676 31084
rect 195242 13152 195298 13161
rect 195242 13087 195298 13096
rect 191102 3496 191158 3505
rect 191102 3431 191158 3440
rect 196728 2174 196756 88946
rect 196806 84824 196862 84833
rect 196806 84759 196862 84768
rect 196820 6186 196848 84759
rect 198016 68950 198044 134506
rect 198108 91769 198136 138654
rect 198094 91760 198150 91769
rect 198094 91695 198150 91704
rect 198096 90364 198148 90370
rect 198096 90306 198148 90312
rect 198004 68944 198056 68950
rect 198004 68886 198056 68892
rect 198108 29714 198136 90306
rect 199396 33794 199424 141374
rect 202144 137352 202196 137358
rect 202144 137294 202196 137300
rect 200856 125656 200908 125662
rect 200856 125598 200908 125604
rect 200764 104984 200816 104990
rect 200764 104926 200816 104932
rect 199474 95840 199530 95849
rect 199474 95775 199530 95784
rect 199488 64870 199516 95775
rect 200776 78674 200804 104926
rect 200868 101454 200896 125598
rect 200856 101448 200908 101454
rect 200856 101390 200908 101396
rect 200764 78668 200816 78674
rect 200764 78610 200816 78616
rect 199476 64864 199528 64870
rect 199476 64806 199528 64812
rect 199384 33788 199436 33794
rect 199384 33730 199436 33736
rect 198096 29708 198148 29714
rect 198096 29650 198148 29656
rect 202156 10402 202184 137294
rect 202248 73817 202276 186895
rect 202340 124982 202368 192510
rect 203628 181490 203656 205527
rect 203524 181484 203576 181490
rect 203524 181426 203576 181432
rect 203616 181484 203668 181490
rect 203616 181426 203668 181432
rect 202328 124976 202380 124982
rect 202328 124918 202380 124924
rect 202326 112432 202382 112441
rect 202326 112367 202382 112376
rect 202234 73808 202290 73817
rect 202234 73743 202290 73752
rect 202340 59362 202368 112367
rect 203536 104281 203564 181426
rect 204916 178673 204944 215319
rect 205008 201414 205036 215902
rect 205100 213217 205128 224159
rect 205376 216617 205404 240244
rect 205928 229094 205956 240244
rect 205928 229066 206416 229094
rect 206284 227792 206336 227798
rect 206284 227734 206336 227740
rect 205638 222184 205694 222193
rect 205638 222119 205694 222128
rect 205652 221649 205680 222119
rect 205638 221640 205694 221649
rect 205638 221575 205694 221584
rect 205362 216608 205418 216617
rect 205362 216543 205418 216552
rect 205376 215393 205404 216543
rect 205362 215384 205418 215393
rect 205362 215319 205418 215328
rect 205086 213208 205142 213217
rect 205086 213143 205142 213152
rect 204996 201408 205048 201414
rect 204996 201350 205048 201356
rect 206296 183025 206324 227734
rect 206388 220833 206416 229066
rect 206480 221649 206508 240244
rect 206848 229090 206876 240244
rect 206836 229084 206888 229090
rect 206836 229026 206888 229032
rect 206848 227798 206876 229026
rect 206928 227928 206980 227934
rect 206928 227870 206980 227876
rect 206836 227792 206888 227798
rect 206836 227734 206888 227740
rect 206466 221640 206522 221649
rect 206466 221575 206522 221584
rect 206374 220824 206430 220833
rect 206374 220759 206430 220768
rect 206388 200802 206416 220759
rect 206376 200796 206428 200802
rect 206376 200738 206428 200744
rect 206940 184249 206968 227870
rect 207400 216753 207428 240244
rect 207952 238754 207980 240244
rect 207676 238746 207980 238754
rect 207664 238740 207980 238746
rect 207716 238726 207980 238740
rect 207664 238682 207716 238688
rect 207386 216744 207442 216753
rect 207386 216679 207442 216688
rect 207676 198082 207704 238682
rect 208320 227934 208348 240244
rect 208400 239420 208452 239426
rect 208400 239362 208452 239368
rect 208412 238746 208440 239362
rect 208400 238740 208452 238746
rect 208400 238682 208452 238688
rect 208872 234433 208900 240244
rect 209042 237416 209098 237425
rect 209042 237351 209098 237360
rect 208858 234424 208914 234433
rect 208858 234359 208914 234368
rect 208308 227928 208360 227934
rect 208308 227870 208360 227876
rect 207754 216744 207810 216753
rect 207754 216679 207810 216688
rect 207664 198076 207716 198082
rect 207664 198018 207716 198024
rect 207768 195974 207796 216679
rect 209056 209710 209084 237351
rect 209240 232937 209268 240244
rect 209792 238754 209820 240244
rect 209792 238726 209912 238754
rect 209686 233880 209742 233889
rect 209686 233815 209742 233824
rect 209226 232928 209282 232937
rect 209226 232863 209282 232872
rect 209044 209704 209096 209710
rect 209044 209646 209096 209652
rect 208400 208412 208452 208418
rect 208400 208354 208452 208360
rect 208412 206825 208440 208354
rect 208398 206816 208454 206825
rect 208398 206751 208454 206760
rect 207756 195968 207808 195974
rect 207756 195910 207808 195916
rect 209056 186969 209084 209646
rect 209700 208418 209728 233815
rect 209884 225010 209912 238726
rect 210344 235657 210372 240244
rect 210330 235648 210386 235657
rect 210330 235583 210386 235592
rect 209872 225004 209924 225010
rect 209872 224946 209924 224952
rect 209884 221785 209912 224946
rect 209870 221776 209926 221785
rect 209870 221711 209926 221720
rect 210712 209774 210740 240244
rect 211264 237425 211292 240244
rect 211250 237416 211306 237425
rect 211250 237351 211306 237360
rect 211816 232937 211844 240244
rect 211802 232928 211858 232937
rect 211802 232863 211858 232872
rect 212184 229094 212212 240244
rect 212630 232928 212686 232937
rect 212630 232863 212686 232872
rect 211816 229066 212212 229094
rect 211068 228472 211120 228478
rect 211068 228414 211120 228420
rect 211080 226234 211108 228414
rect 211816 226370 211844 229066
rect 211804 226364 211856 226370
rect 211804 226306 211856 226312
rect 211068 226228 211120 226234
rect 211068 226170 211120 226176
rect 210436 209746 210740 209774
rect 210436 209545 210464 209746
rect 210422 209536 210478 209545
rect 210422 209471 210478 209480
rect 209688 208412 209740 208418
rect 209688 208354 209740 208360
rect 209042 186960 209098 186969
rect 209042 186895 209098 186904
rect 206926 184240 206982 184249
rect 206926 184175 206982 184184
rect 206282 183016 206338 183025
rect 206282 182951 206338 182960
rect 204902 178664 204958 178673
rect 204902 178599 204958 178608
rect 204904 176044 204956 176050
rect 204904 175986 204956 175992
rect 203616 136672 203668 136678
rect 203616 136614 203668 136620
rect 203522 104272 203578 104281
rect 203522 104207 203578 104216
rect 203524 98116 203576 98122
rect 203524 98058 203576 98064
rect 203536 60722 203564 98058
rect 203628 84153 203656 136614
rect 203614 84144 203670 84153
rect 203614 84079 203670 84088
rect 203524 60716 203576 60722
rect 203524 60658 203576 60664
rect 202328 59356 202380 59362
rect 202328 59298 202380 59304
rect 204916 35290 204944 175986
rect 204996 145580 205048 145586
rect 204996 145522 205048 145528
rect 204904 35284 204956 35290
rect 204904 35226 204956 35232
rect 205008 26926 205036 145522
rect 209044 141500 209096 141506
rect 209044 141442 209096 141448
rect 206282 132560 206338 132569
rect 206282 132495 206338 132504
rect 206296 92313 206324 132495
rect 206374 115968 206430 115977
rect 206374 115903 206430 115912
rect 206388 93226 206416 115903
rect 206376 93220 206428 93226
rect 206376 93162 206428 93168
rect 206282 92304 206338 92313
rect 206282 92239 206338 92248
rect 206284 84924 206336 84930
rect 206284 84866 206336 84872
rect 205088 40792 205140 40798
rect 205088 40734 205140 40740
rect 205100 26994 205128 40734
rect 206296 33862 206324 84866
rect 206284 33856 206336 33862
rect 206284 33798 206336 33804
rect 205088 26988 205140 26994
rect 205088 26930 205140 26936
rect 204996 26920 205048 26926
rect 204996 26862 205048 26868
rect 209056 25634 209084 141442
rect 209226 120728 209282 120737
rect 209226 120663 209282 120672
rect 209134 104136 209190 104145
rect 209134 104071 209190 104080
rect 209148 73166 209176 104071
rect 209240 97306 209268 120663
rect 210436 97986 210464 209471
rect 211816 200025 211844 226306
rect 212644 219434 212672 232863
rect 212632 219428 212684 219434
rect 212632 219370 212684 219376
rect 212644 210458 212672 219370
rect 212632 210452 212684 210458
rect 212632 210394 212684 210400
rect 211802 200016 211858 200025
rect 211802 199951 211858 199960
rect 212736 194546 212764 240244
rect 213104 237425 213132 240244
rect 213656 238754 213684 240244
rect 213656 238726 213868 238754
rect 213656 238649 213684 238726
rect 213642 238640 213698 238649
rect 213642 238575 213698 238584
rect 213090 237416 213146 237425
rect 213090 237351 213146 237360
rect 213736 204264 213788 204270
rect 213736 204206 213788 204212
rect 213748 203017 213776 204206
rect 213734 203008 213790 203017
rect 213734 202943 213790 202952
rect 212724 194540 212776 194546
rect 212724 194482 212776 194488
rect 213840 194041 213868 238726
rect 214208 238678 214236 240244
rect 214196 238672 214248 238678
rect 214196 238614 214248 238620
rect 214208 232558 214236 238614
rect 214576 237289 214604 240244
rect 214562 237280 214618 237289
rect 214562 237215 214618 237224
rect 214656 233912 214708 233918
rect 214656 233854 214708 233860
rect 214564 233164 214616 233170
rect 214564 233106 214616 233112
rect 214196 232552 214248 232558
rect 214196 232494 214248 232500
rect 214576 203590 214604 233106
rect 214668 221542 214696 233854
rect 215128 233170 215156 240244
rect 215116 233164 215168 233170
rect 215116 233106 215168 233112
rect 214656 221536 214708 221542
rect 214656 221478 214708 221484
rect 215208 221468 215260 221474
rect 215208 221410 215260 221416
rect 215220 218890 215248 221410
rect 215208 218884 215260 218890
rect 215208 218826 215260 218832
rect 214656 207664 214708 207670
rect 214656 207606 214708 207612
rect 214668 207097 214696 207606
rect 214654 207088 214710 207097
rect 214654 207023 214710 207032
rect 214564 203584 214616 203590
rect 214564 203526 214616 203532
rect 214668 195401 214696 207023
rect 215680 204202 215708 240244
rect 216048 234569 216076 240244
rect 216600 238406 216628 240244
rect 216588 238400 216640 238406
rect 216588 238342 216640 238348
rect 216034 234560 216090 234569
rect 216034 234495 216090 234504
rect 216678 234016 216734 234025
rect 216678 233951 216734 233960
rect 215944 233844 215996 233850
rect 215944 233786 215996 233792
rect 215668 204196 215720 204202
rect 215668 204138 215720 204144
rect 215680 200114 215708 204138
rect 215956 204105 215984 233786
rect 216692 231810 216720 233951
rect 216680 231804 216732 231810
rect 216680 231746 216732 231752
rect 217152 229094 217180 240244
rect 217152 229066 217272 229094
rect 217244 217977 217272 229066
rect 217322 222320 217378 222329
rect 217322 222255 217378 222264
rect 217230 217968 217286 217977
rect 217336 217938 217364 222255
rect 217230 217903 217286 217912
rect 217324 217932 217376 217938
rect 217244 217297 217272 217903
rect 217324 217874 217376 217880
rect 217230 217288 217286 217297
rect 217230 217223 217286 217232
rect 217520 211041 217548 240244
rect 218072 238754 218100 240244
rect 218072 238726 218192 238754
rect 218060 238400 218112 238406
rect 218060 238342 218112 238348
rect 218072 238105 218100 238342
rect 218058 238096 218114 238105
rect 218058 238031 218114 238040
rect 218164 237522 218192 238726
rect 218152 237516 218204 237522
rect 218152 237458 218204 237464
rect 217506 211032 217562 211041
rect 217506 210967 217562 210976
rect 215942 204096 215998 204105
rect 215942 204031 215998 204040
rect 217520 200114 217548 210967
rect 215680 200086 216076 200114
rect 214654 195392 214710 195401
rect 214654 195327 214710 195336
rect 213826 194032 213882 194041
rect 213826 193967 213882 193976
rect 216048 177993 216076 200086
rect 217428 200086 217548 200114
rect 217324 190528 217376 190534
rect 217324 190470 217376 190476
rect 216034 177984 216090 177993
rect 216034 177919 216090 177928
rect 217336 169046 217364 190470
rect 217428 189786 217456 200086
rect 218440 190505 218468 240244
rect 218704 237516 218756 237522
rect 218704 237458 218756 237464
rect 218716 227633 218744 237458
rect 218702 227624 218758 227633
rect 218702 227559 218758 227568
rect 218704 222964 218756 222970
rect 218704 222906 218756 222912
rect 218716 192545 218744 222906
rect 218992 214033 219020 240244
rect 219544 238754 219572 240244
rect 219912 238754 219940 240244
rect 219544 238726 219664 238754
rect 219912 238746 220216 238754
rect 219636 222154 219664 238726
rect 219900 238740 220216 238746
rect 219952 238726 220216 238740
rect 219900 238682 219952 238688
rect 220084 237516 220136 237522
rect 220084 237458 220136 237464
rect 219624 222148 219676 222154
rect 219624 222090 219676 222096
rect 218978 214024 219034 214033
rect 218978 213959 219034 213968
rect 218992 207670 219020 213959
rect 218980 207664 219032 207670
rect 218980 207606 219032 207612
rect 220096 198665 220124 237458
rect 220188 228410 220216 238726
rect 220464 233238 220492 240244
rect 220818 239456 220874 239465
rect 220818 239391 220874 239400
rect 220832 238746 220860 239391
rect 220820 238740 220872 238746
rect 220820 238682 220872 238688
rect 221016 233850 221044 240244
rect 221004 233844 221056 233850
rect 221004 233786 221056 233792
rect 220452 233232 220504 233238
rect 220452 233174 220504 233180
rect 220728 233232 220780 233238
rect 220728 233174 220780 233180
rect 220740 231198 220768 233174
rect 220728 231192 220780 231198
rect 220728 231134 220780 231140
rect 220176 228404 220228 228410
rect 220176 228346 220228 228352
rect 221384 201482 221412 240244
rect 221936 237522 221964 240244
rect 222304 238746 222332 240244
rect 222856 238754 222884 240244
rect 222292 238740 222344 238746
rect 222292 238682 222344 238688
rect 222396 238726 222884 238754
rect 222304 237522 222332 238682
rect 221924 237516 221976 237522
rect 221924 237458 221976 237464
rect 222292 237516 222344 237522
rect 222292 237458 222344 237464
rect 222106 233880 222162 233889
rect 222106 233815 222108 233824
rect 222160 233815 222162 233824
rect 222108 233786 222160 233792
rect 221464 229764 221516 229770
rect 221464 229706 221516 229712
rect 221476 217841 221504 229706
rect 222396 226302 222424 238726
rect 223408 238649 223436 240244
rect 223394 238640 223450 238649
rect 223394 238575 223450 238584
rect 222844 237516 222896 237522
rect 222844 237458 222896 237464
rect 222936 237516 222988 237522
rect 222936 237458 222988 237464
rect 222384 226296 222436 226302
rect 222384 226238 222436 226244
rect 222396 225078 222424 226238
rect 222384 225072 222436 225078
rect 222384 225014 222436 225020
rect 221462 217832 221518 217841
rect 221462 217767 221518 217776
rect 222856 206310 222884 237458
rect 222948 227662 222976 237458
rect 223408 232529 223436 238575
rect 223776 237522 223804 240244
rect 224328 239873 224356 240244
rect 224314 239864 224370 239873
rect 224314 239799 224370 239808
rect 224328 239465 224356 239799
rect 224314 239456 224370 239465
rect 224314 239391 224370 239400
rect 224776 238128 224828 238134
rect 224776 238070 224828 238076
rect 224788 237969 224816 238070
rect 224774 237960 224830 237969
rect 224774 237895 224830 237904
rect 223764 237516 223816 237522
rect 223764 237458 223816 237464
rect 223394 232520 223450 232529
rect 223394 232455 223450 232464
rect 224222 231704 224278 231713
rect 224222 231639 224278 231648
rect 222936 227656 222988 227662
rect 222936 227598 222988 227604
rect 222844 206304 222896 206310
rect 222844 206246 222896 206252
rect 221372 201476 221424 201482
rect 221372 201418 221424 201424
rect 222948 199481 222976 227598
rect 223028 225072 223080 225078
rect 223028 225014 223080 225020
rect 223040 210497 223068 225014
rect 224236 218822 224264 231639
rect 224224 218816 224276 218822
rect 224224 218758 224276 218764
rect 223026 210488 223082 210497
rect 223026 210423 223082 210432
rect 222934 199472 222990 199481
rect 222934 199407 222990 199416
rect 220082 198656 220138 198665
rect 220082 198591 220138 198600
rect 218702 192536 218758 192545
rect 218702 192471 218758 192480
rect 218426 190496 218482 190505
rect 218426 190431 218482 190440
rect 217416 189780 217468 189786
rect 217416 189722 217468 189728
rect 218440 189038 218468 190431
rect 218428 189032 218480 189038
rect 218428 188974 218480 188980
rect 220082 178120 220138 178129
rect 220082 178055 220138 178064
rect 217324 169040 217376 169046
rect 217324 168982 217376 168988
rect 220096 155854 220124 178055
rect 221464 163532 221516 163538
rect 221464 163474 221516 163480
rect 220084 155848 220136 155854
rect 220084 155790 220136 155796
rect 213184 155236 213236 155242
rect 213184 155178 213236 155184
rect 211896 129804 211948 129810
rect 211896 129746 211948 129752
rect 211804 109132 211856 109138
rect 211804 109074 211856 109080
rect 210424 97980 210476 97986
rect 210424 97922 210476 97928
rect 209228 97300 209280 97306
rect 209228 97242 209280 97248
rect 211816 82822 211844 109074
rect 211908 104174 211936 129746
rect 211896 104168 211948 104174
rect 211896 104110 211948 104116
rect 211804 82816 211856 82822
rect 211804 82758 211856 82764
rect 209136 73160 209188 73166
rect 209136 73102 209188 73108
rect 213196 39438 213224 155178
rect 214564 153264 214616 153270
rect 214564 153206 214616 153212
rect 213276 129872 213328 129878
rect 213276 129814 213328 129820
rect 213288 64802 213316 129814
rect 214576 96014 214604 153206
rect 217324 152516 217376 152522
rect 217324 152458 217376 152464
rect 214656 151836 214708 151842
rect 214656 151778 214708 151784
rect 214668 126274 214696 151778
rect 214656 126268 214708 126274
rect 214656 126210 214708 126216
rect 214656 99408 214708 99414
rect 214656 99350 214708 99356
rect 214564 96008 214616 96014
rect 214564 95950 214616 95956
rect 214668 74526 214696 99350
rect 214656 74520 214708 74526
rect 214656 74462 214708 74468
rect 214562 73944 214618 73953
rect 214562 73879 214618 73888
rect 213276 64796 213328 64802
rect 213276 64738 213328 64744
rect 213184 39432 213236 39438
rect 213184 39374 213236 39380
rect 209044 25628 209096 25634
rect 209044 25570 209096 25576
rect 214576 13122 214604 73879
rect 214656 58676 214708 58682
rect 214656 58618 214708 58624
rect 214668 40798 214696 58618
rect 217336 40798 217364 152458
rect 218796 145648 218848 145654
rect 218796 145590 218848 145596
rect 218702 104272 218758 104281
rect 218702 104207 218758 104216
rect 214656 40792 214708 40798
rect 214656 40734 214708 40740
rect 217324 40792 217376 40798
rect 217324 40734 217376 40740
rect 214564 13116 214616 13122
rect 214564 13058 214616 13064
rect 202144 10396 202196 10402
rect 202144 10338 202196 10344
rect 196808 6180 196860 6186
rect 196808 6122 196860 6128
rect 218716 4865 218744 104207
rect 218808 101454 218836 145590
rect 220084 135924 220136 135930
rect 220084 135866 220136 135872
rect 218796 101448 218848 101454
rect 218796 101390 218848 101396
rect 220096 11665 220124 135866
rect 220176 125724 220228 125730
rect 220176 125666 220228 125672
rect 220188 63510 220216 125666
rect 221476 83502 221504 163474
rect 222936 151904 222988 151910
rect 222936 151846 222988 151852
rect 222842 141400 222898 141409
rect 222842 141335 222898 141344
rect 222856 120766 222884 141335
rect 222948 137290 222976 151846
rect 224224 140820 224276 140826
rect 224224 140762 224276 140768
rect 222936 137284 222988 137290
rect 222936 137226 222988 137232
rect 222844 120760 222896 120766
rect 222844 120702 222896 120708
rect 224236 112470 224264 140762
rect 224788 119377 224816 237895
rect 224880 231713 224908 240244
rect 225248 240145 225276 240244
rect 225234 240136 225290 240145
rect 225234 240071 225290 240080
rect 224866 231704 224922 231713
rect 224866 231639 224922 231648
rect 224868 218748 224920 218754
rect 224868 218690 224920 218696
rect 224880 218113 224908 218690
rect 225800 218113 225828 240244
rect 224866 218104 224922 218113
rect 224866 218039 224922 218048
rect 225786 218104 225842 218113
rect 225786 218039 225842 218048
rect 224774 119368 224830 119377
rect 224774 119303 224830 119312
rect 224316 116000 224368 116006
rect 224316 115942 224368 115948
rect 224224 112464 224276 112470
rect 224224 112406 224276 112412
rect 224328 91050 224356 115942
rect 224880 96014 224908 218039
rect 226168 205465 226196 240244
rect 226720 238134 226748 240244
rect 226708 238128 226760 238134
rect 226708 238070 226760 238076
rect 226984 238060 227036 238066
rect 226984 238002 227036 238008
rect 226996 215937 227024 238002
rect 226982 215928 227038 215937
rect 226982 215863 227038 215872
rect 227272 210905 227300 240244
rect 227640 238649 227668 240244
rect 228192 240145 228220 240244
rect 228178 240136 228234 240145
rect 228178 240071 228234 240080
rect 228744 240009 228772 240244
rect 228730 240000 228786 240009
rect 228730 239935 228786 239944
rect 227626 238640 227682 238649
rect 227626 238575 227682 238584
rect 229112 225078 229140 240244
rect 229664 229770 229692 240244
rect 230216 234025 230244 240244
rect 230584 238241 230612 240244
rect 230570 238232 230626 238241
rect 230570 238167 230626 238176
rect 230202 234016 230258 234025
rect 230202 233951 230258 233960
rect 229652 229764 229704 229770
rect 229652 229706 229704 229712
rect 229100 225072 229152 225078
rect 229100 225014 229152 225020
rect 229744 225072 229796 225078
rect 229744 225014 229796 225020
rect 227258 210896 227314 210905
rect 227258 210831 227314 210840
rect 226154 205456 226210 205465
rect 226154 205391 226210 205400
rect 226168 200870 226196 205391
rect 226156 200864 226208 200870
rect 226156 200806 226208 200812
rect 227272 200114 227300 210831
rect 229756 206961 229784 225014
rect 231136 209778 231164 240244
rect 231504 233209 231532 240244
rect 231952 240168 232004 240174
rect 231950 240136 231952 240145
rect 232004 240136 232006 240145
rect 231950 240071 232006 240080
rect 231490 233200 231546 233209
rect 231490 233135 231546 233144
rect 232056 231946 232084 240244
rect 232502 239592 232558 239601
rect 232502 239527 232558 239536
rect 232044 231940 232096 231946
rect 232044 231882 232096 231888
rect 231124 209772 231176 209778
rect 231124 209714 231176 209720
rect 231136 209098 231164 209714
rect 231124 209092 231176 209098
rect 231124 209034 231176 209040
rect 229742 206952 229798 206961
rect 229742 206887 229798 206896
rect 226996 200086 227300 200114
rect 226996 182889 227024 200086
rect 228362 189952 228418 189961
rect 228362 189887 228418 189896
rect 227718 183152 227774 183161
rect 227718 183087 227774 183096
rect 226982 182880 227038 182889
rect 226982 182815 227038 182824
rect 227732 178022 227760 183087
rect 227720 178016 227772 178022
rect 227720 177958 227772 177964
rect 226984 148368 227036 148374
rect 226984 148310 227036 148316
rect 225604 120148 225656 120154
rect 225604 120090 225656 120096
rect 224868 96008 224920 96014
rect 224868 95950 224920 95956
rect 224316 91044 224368 91050
rect 224316 90986 224368 90992
rect 221464 83496 221516 83502
rect 221464 83438 221516 83444
rect 224222 74080 224278 74089
rect 224222 74015 224278 74024
rect 220176 63504 220228 63510
rect 220176 63446 220228 63452
rect 224236 14550 224264 74015
rect 225616 52426 225644 120090
rect 226996 90409 227024 148310
rect 226982 90400 227038 90409
rect 226982 90335 227038 90344
rect 225604 52420 225656 52426
rect 225604 52362 225656 52368
rect 224224 14544 224276 14550
rect 224224 14486 224276 14492
rect 220082 11656 220138 11665
rect 220082 11591 220138 11600
rect 218702 4856 218758 4865
rect 218702 4791 218758 4800
rect 228376 3602 228404 189887
rect 231124 185632 231176 185638
rect 231124 185574 231176 185580
rect 229836 140888 229888 140894
rect 229836 140830 229888 140836
rect 229744 127084 229796 127090
rect 229744 127026 229796 127032
rect 228456 124976 228508 124982
rect 228456 124918 228508 124924
rect 228468 24177 228496 124918
rect 229756 93945 229784 127026
rect 229848 108322 229876 140830
rect 230480 113280 230532 113286
rect 230480 113222 230532 113228
rect 230492 113150 230520 113222
rect 230480 113144 230532 113150
rect 230480 113086 230532 113092
rect 229836 108316 229888 108322
rect 229836 108258 229888 108264
rect 229742 93936 229798 93945
rect 229742 93871 229798 93880
rect 229834 93120 229890 93129
rect 229834 93055 229890 93064
rect 229744 77988 229796 77994
rect 229744 77930 229796 77936
rect 228454 24168 228510 24177
rect 228454 24103 228510 24112
rect 228364 3596 228416 3602
rect 228364 3538 228416 3544
rect 229756 3466 229784 77930
rect 229848 35222 229876 93055
rect 229836 35216 229888 35222
rect 229836 35158 229888 35164
rect 231136 3534 231164 185574
rect 231216 182232 231268 182238
rect 231216 182174 231268 182180
rect 231228 164150 231256 182174
rect 231584 179444 231636 179450
rect 231584 179386 231636 179392
rect 231596 173806 231624 179386
rect 231584 173800 231636 173806
rect 231584 173742 231636 173748
rect 231216 164144 231268 164150
rect 231216 164086 231268 164092
rect 231216 144968 231268 144974
rect 231216 144910 231268 144916
rect 231228 89049 231256 144910
rect 231306 135552 231362 135561
rect 231306 135487 231362 135496
rect 231320 123486 231348 135487
rect 231308 123480 231360 123486
rect 231308 123422 231360 123428
rect 231308 107704 231360 107710
rect 231308 107646 231360 107652
rect 231214 89040 231270 89049
rect 231214 88975 231270 88984
rect 231320 84182 231348 107646
rect 231308 84176 231360 84182
rect 231308 84118 231360 84124
rect 231124 3528 231176 3534
rect 231124 3470 231176 3476
rect 229744 3460 229796 3466
rect 229744 3402 229796 3408
rect 232516 3369 232544 239527
rect 232608 238513 232636 240244
rect 232686 240000 232742 240009
rect 232686 239935 232742 239944
rect 232594 238504 232650 238513
rect 232594 238439 232650 238448
rect 232594 229936 232650 229945
rect 232594 229871 232650 229880
rect 232608 205057 232636 229871
rect 232700 221474 232728 239935
rect 232976 231849 233004 240244
rect 233148 231940 233200 231946
rect 233148 231882 233200 231888
rect 232962 231840 233018 231849
rect 232962 231775 233018 231784
rect 233160 230382 233188 231882
rect 233148 230376 233200 230382
rect 233148 230318 233200 230324
rect 232688 221468 232740 221474
rect 232688 221410 232740 221416
rect 232594 205048 232650 205057
rect 232594 204983 232650 204992
rect 233148 204944 233200 204950
rect 233148 204886 233200 204892
rect 233160 188358 233188 204886
rect 233528 202881 233556 240244
rect 233884 237448 233936 237454
rect 233884 237390 233936 237396
rect 233896 229945 233924 237390
rect 234080 234666 234108 240244
rect 234068 234660 234120 234666
rect 234068 234602 234120 234608
rect 234080 233073 234108 234602
rect 234066 233064 234122 233073
rect 234066 232999 234122 233008
rect 233882 229936 233938 229945
rect 233882 229871 233938 229880
rect 233976 221536 234028 221542
rect 233976 221478 234028 221484
rect 233514 202872 233570 202881
rect 233514 202807 233570 202816
rect 233884 199436 233936 199442
rect 233884 199378 233936 199384
rect 232596 188352 232648 188358
rect 232596 188294 232648 188300
rect 233148 188352 233200 188358
rect 233148 188294 233200 188300
rect 232608 180169 232636 188294
rect 232594 180160 232650 180169
rect 232594 180095 232650 180104
rect 232688 139460 232740 139466
rect 232688 139402 232740 139408
rect 232700 124914 232728 139402
rect 232688 124908 232740 124914
rect 232688 124850 232740 124856
rect 232596 124228 232648 124234
rect 232596 124170 232648 124176
rect 232608 89690 232636 124170
rect 232596 89684 232648 89690
rect 232596 89626 232648 89632
rect 232594 87544 232650 87553
rect 232594 87479 232650 87488
rect 232608 31074 232636 87479
rect 232596 31068 232648 31074
rect 232596 31010 232648 31016
rect 233896 6186 233924 199378
rect 233988 193934 234016 221478
rect 234448 204950 234476 240244
rect 235000 224913 235028 240244
rect 235368 238513 235396 240244
rect 235816 240168 235868 240174
rect 235920 240122 235948 240244
rect 235868 240116 235948 240122
rect 235816 240110 235948 240116
rect 235828 240094 235948 240110
rect 236472 238649 236500 240244
rect 236458 238640 236514 238649
rect 236458 238575 236514 238584
rect 235354 238504 235410 238513
rect 235354 238439 235410 238448
rect 234986 224904 235042 224913
rect 234986 224839 235042 224848
rect 236840 219434 236868 240244
rect 237392 237454 237420 240244
rect 237944 240145 237972 240244
rect 237930 240136 237986 240145
rect 237930 240071 237986 240080
rect 237380 237448 237432 237454
rect 237944 237425 237972 240071
rect 237380 237390 237432 237396
rect 237930 237416 237986 237425
rect 237930 237351 237986 237360
rect 238022 221640 238078 221649
rect 238022 221575 238078 221584
rect 236748 219406 236868 219434
rect 236748 215393 236776 219406
rect 235998 215384 236054 215393
rect 235998 215319 236054 215328
rect 236734 215384 236790 215393
rect 236734 215319 236790 215328
rect 236012 215218 236040 215319
rect 236000 215212 236052 215218
rect 236000 215154 236052 215160
rect 234436 204944 234488 204950
rect 234436 204886 234488 204892
rect 233976 193928 234028 193934
rect 233976 193870 234028 193876
rect 236644 193860 236696 193866
rect 236644 193802 236696 193808
rect 233976 183592 234028 183598
rect 233976 183534 234028 183540
rect 233988 172446 234016 183534
rect 233976 172440 234028 172446
rect 233976 172382 234028 172388
rect 233976 138712 234028 138718
rect 233976 138654 234028 138660
rect 233988 74458 234016 138654
rect 235264 135380 235316 135386
rect 235264 135322 235316 135328
rect 234066 133104 234122 133113
rect 234066 133039 234122 133048
rect 234080 98705 234108 133039
rect 234160 107772 234212 107778
rect 234160 107714 234212 107720
rect 234066 98696 234122 98705
rect 234066 98631 234122 98640
rect 234172 81394 234200 107714
rect 235276 91798 235304 135322
rect 236000 117360 236052 117366
rect 236000 117302 236052 117308
rect 236012 116618 236040 117302
rect 236000 116612 236052 116618
rect 236000 116554 236052 116560
rect 235356 113280 235408 113286
rect 235356 113222 235408 113228
rect 235264 91792 235316 91798
rect 235264 91734 235316 91740
rect 235368 88330 235396 113222
rect 235908 91792 235960 91798
rect 235908 91734 235960 91740
rect 235356 88324 235408 88330
rect 235356 88266 235408 88272
rect 234160 81388 234212 81394
rect 234160 81330 234212 81336
rect 233976 74452 234028 74458
rect 233976 74394 234028 74400
rect 235920 6914 235948 91734
rect 236656 89049 236684 193802
rect 238036 181558 238064 221575
rect 238312 216345 238340 240244
rect 238864 238066 238892 240244
rect 239232 240009 239260 240244
rect 239218 240000 239274 240009
rect 239218 239935 239274 239944
rect 238852 238060 238904 238066
rect 238852 238002 238904 238008
rect 238666 237416 238722 237425
rect 238666 237351 238722 237360
rect 238680 221542 238708 237351
rect 239784 226273 239812 240244
rect 240336 239494 240364 240244
rect 240324 239488 240376 239494
rect 240324 239430 240376 239436
rect 240336 238066 240364 239430
rect 240324 238060 240376 238066
rect 240324 238002 240376 238008
rect 240704 237153 240732 240244
rect 240784 237448 240836 237454
rect 240784 237390 240836 237396
rect 240690 237144 240746 237153
rect 240690 237079 240746 237088
rect 240796 233306 240824 237390
rect 240784 233300 240836 233306
rect 240784 233242 240836 233248
rect 239770 226264 239826 226273
rect 239770 226199 239826 226208
rect 238668 221536 238720 221542
rect 238668 221478 238720 221484
rect 238298 216336 238354 216345
rect 238298 216271 238354 216280
rect 240796 215966 240824 233242
rect 241256 231742 241284 240244
rect 241808 238649 241836 240244
rect 241794 238640 241850 238649
rect 241794 238575 241850 238584
rect 242176 238377 242204 240244
rect 242254 239456 242310 239465
rect 242254 239391 242310 239400
rect 242162 238368 242218 238377
rect 242162 238303 242218 238312
rect 241244 231736 241296 231742
rect 241244 231678 241296 231684
rect 241428 231736 241480 231742
rect 241428 231678 241480 231684
rect 241440 231130 241468 231678
rect 241428 231124 241480 231130
rect 241428 231066 241480 231072
rect 240784 215960 240836 215966
rect 240784 215902 240836 215908
rect 242164 211812 242216 211818
rect 242164 211754 242216 211760
rect 240782 192672 240838 192681
rect 240782 192607 240838 192616
rect 238024 181552 238076 181558
rect 238024 181494 238076 181500
rect 238114 180840 238170 180849
rect 238114 180775 238170 180784
rect 237380 178016 237432 178022
rect 237380 177958 237432 177964
rect 237392 176769 237420 177958
rect 238022 177032 238078 177041
rect 238022 176967 238078 176976
rect 237378 176760 237434 176769
rect 237378 176695 237434 176704
rect 238036 161362 238064 176967
rect 238128 166025 238156 180775
rect 238114 166016 238170 166025
rect 238114 165951 238170 165960
rect 238024 161356 238076 161362
rect 238024 161298 238076 161304
rect 240138 160712 240194 160721
rect 240138 160647 240194 160656
rect 238024 143676 238076 143682
rect 238024 143618 238076 143624
rect 238036 122126 238064 143618
rect 238116 124296 238168 124302
rect 238116 124238 238168 124244
rect 238024 122120 238076 122126
rect 238024 122062 238076 122068
rect 236736 120760 236788 120766
rect 236736 120702 236788 120708
rect 236748 91050 236776 120702
rect 238024 120216 238076 120222
rect 238024 120158 238076 120164
rect 236736 91044 236788 91050
rect 236736 90986 236788 90992
rect 236642 89040 236698 89049
rect 236642 88975 236698 88984
rect 236642 87680 236698 87689
rect 236642 87615 236698 87624
rect 235998 61568 236054 61577
rect 235998 61503 236054 61512
rect 236012 58682 236040 61503
rect 236000 58676 236052 58682
rect 236000 58618 236052 58624
rect 236656 47598 236684 87615
rect 238036 62082 238064 120158
rect 238128 93906 238156 124238
rect 239404 121576 239456 121582
rect 239404 121518 239456 121524
rect 238208 114572 238260 114578
rect 238208 114514 238260 114520
rect 238116 93900 238168 93906
rect 238116 93842 238168 93848
rect 238220 91089 238248 114514
rect 238206 91080 238262 91089
rect 238206 91015 238262 91024
rect 238114 86184 238170 86193
rect 238114 86119 238170 86128
rect 238024 62076 238076 62082
rect 238024 62018 238076 62024
rect 236644 47592 236696 47598
rect 236644 47534 236696 47540
rect 238024 47592 238076 47598
rect 238024 47534 238076 47540
rect 236642 32464 236698 32473
rect 236642 32399 236698 32408
rect 236656 17338 236684 32399
rect 238036 18630 238064 47534
rect 238128 28257 238156 86119
rect 239416 53786 239444 121518
rect 239404 53780 239456 53786
rect 239404 53722 239456 53728
rect 238114 28248 238170 28257
rect 238114 28183 238170 28192
rect 238024 18624 238076 18630
rect 238024 18566 238076 18572
rect 236644 17332 236696 17338
rect 236644 17274 236696 17280
rect 238024 17264 238076 17270
rect 238024 17206 238076 17212
rect 235828 6886 235948 6914
rect 233884 6180 233936 6186
rect 233884 6122 233936 6128
rect 232502 3360 232558 3369
rect 232502 3295 232558 3304
rect 196716 2168 196768 2174
rect 196716 2110 196768 2116
rect 235828 480 235856 6886
rect 238036 2174 238064 17206
rect 239312 3596 239364 3602
rect 239312 3538 239364 3544
rect 238024 2168 238076 2174
rect 238024 2110 238076 2116
rect 239324 480 239352 3538
rect 240152 490 240180 160647
rect 240796 15978 240824 192607
rect 242176 189854 242204 211754
rect 242268 192574 242296 239391
rect 242728 237386 242756 240244
rect 243280 237454 243308 240244
rect 243268 237448 243320 237454
rect 243268 237390 243320 237396
rect 242716 237380 242768 237386
rect 242716 237322 242768 237328
rect 243648 235958 243676 240244
rect 243636 235952 243688 235958
rect 243636 235894 243688 235900
rect 243648 235278 243676 235894
rect 243636 235272 243688 235278
rect 242346 235240 242402 235249
rect 243636 235214 243688 235220
rect 242346 235175 242402 235184
rect 242360 225593 242388 235175
rect 242346 225584 242402 225593
rect 242346 225519 242402 225528
rect 244016 209681 244044 241295
rect 244096 240780 244148 240786
rect 244096 240722 244148 240728
rect 244108 234569 244136 240722
rect 244280 237448 244332 237454
rect 244280 237390 244332 237396
rect 244094 234560 244150 234569
rect 244094 234495 244150 234504
rect 244002 209672 244058 209681
rect 244002 209607 244058 209616
rect 244292 208350 244320 237390
rect 244384 227361 244412 247279
rect 244370 227352 244426 227361
rect 244370 227287 244426 227296
rect 244476 219337 244504 255983
rect 244660 235793 244688 278831
rect 245660 276140 245712 276146
rect 245660 276082 245712 276088
rect 245672 271017 245700 276082
rect 245764 273170 245792 305594
rect 245844 294636 245896 294642
rect 245844 294578 245896 294584
rect 245856 276282 245884 294578
rect 245934 294536 245990 294545
rect 245934 294471 245990 294480
rect 245844 276276 245896 276282
rect 245844 276218 245896 276224
rect 245948 276162 245976 294471
rect 246040 276729 246068 315250
rect 246316 312594 246344 343606
rect 247132 330608 247184 330614
rect 247132 330550 247184 330556
rect 246304 312588 246356 312594
rect 246304 312530 246356 312536
rect 247040 304292 247092 304298
rect 247040 304234 247092 304240
rect 246304 300892 246356 300898
rect 246304 300834 246356 300840
rect 246316 294642 246344 300834
rect 246304 294636 246356 294642
rect 246304 294578 246356 294584
rect 246120 282872 246172 282878
rect 246120 282814 246172 282820
rect 246132 281625 246160 282814
rect 246118 281616 246174 281625
rect 246118 281551 246174 281560
rect 246120 281512 246172 281518
rect 246120 281454 246172 281460
rect 246132 280265 246160 281454
rect 246118 280256 246174 280265
rect 246118 280191 246174 280200
rect 246118 279440 246174 279449
rect 246118 279375 246174 279384
rect 246132 278798 246160 279375
rect 246120 278792 246172 278798
rect 246120 278734 246172 278740
rect 246120 278044 246172 278050
rect 246120 277986 246172 277992
rect 246132 277545 246160 277986
rect 246118 277536 246174 277545
rect 246118 277471 246174 277480
rect 246026 276720 246082 276729
rect 246026 276655 246028 276664
rect 246080 276655 246082 276664
rect 246028 276626 246080 276632
rect 246040 276595 246068 276626
rect 246028 276276 246080 276282
rect 246028 276218 246080 276224
rect 245856 276134 245976 276162
rect 245856 274530 245884 276134
rect 245936 276004 245988 276010
rect 245936 275946 245988 275952
rect 245948 275913 245976 275946
rect 245934 275904 245990 275913
rect 245934 275839 245990 275848
rect 245934 274544 245990 274553
rect 245856 274502 245934 274530
rect 245934 274479 245990 274488
rect 245948 273970 245976 274479
rect 245936 273964 245988 273970
rect 245936 273906 245988 273912
rect 245842 273728 245898 273737
rect 245842 273663 245898 273672
rect 245856 273290 245884 273663
rect 245844 273284 245896 273290
rect 245844 273226 245896 273232
rect 245934 273184 245990 273193
rect 245764 273142 245884 273170
rect 245856 272542 245884 273142
rect 245934 273119 245990 273128
rect 245948 272610 245976 273119
rect 245936 272604 245988 272610
rect 245936 272546 245988 272552
rect 245844 272536 245896 272542
rect 246040 272490 246068 276218
rect 245844 272478 245896 272484
rect 245856 272377 245884 272478
rect 245948 272462 246068 272490
rect 245842 272368 245898 272377
rect 245842 272303 245898 272312
rect 245750 271552 245806 271561
rect 245750 271487 245806 271496
rect 245764 271182 245792 271487
rect 245752 271176 245804 271182
rect 245752 271118 245804 271124
rect 245658 271008 245714 271017
rect 245658 270943 245714 270952
rect 245660 270496 245712 270502
rect 245660 270438 245712 270444
rect 245672 270201 245700 270438
rect 245658 270192 245714 270201
rect 245658 270127 245714 270136
rect 245948 269822 245976 272462
rect 246302 271008 246358 271017
rect 246302 270943 246358 270952
rect 245936 269816 245988 269822
rect 245936 269758 245988 269764
rect 245948 269657 245976 269758
rect 245934 269648 245990 269657
rect 245934 269583 245990 269592
rect 245936 268388 245988 268394
rect 245936 268330 245988 268336
rect 245948 268025 245976 268330
rect 245934 268016 245990 268025
rect 245934 267951 245990 267960
rect 246026 267472 246082 267481
rect 246026 267407 246082 267416
rect 245936 267028 245988 267034
rect 245936 266970 245988 266976
rect 245948 266665 245976 266970
rect 245934 266656 245990 266665
rect 245934 266591 245990 266600
rect 246040 266422 246068 267407
rect 246028 266416 246080 266422
rect 246028 266358 246080 266364
rect 245752 266348 245804 266354
rect 245752 266290 245804 266296
rect 245764 265305 245792 266290
rect 245844 266280 245896 266286
rect 245844 266222 245896 266228
rect 245856 265849 245884 266222
rect 245842 265840 245898 265849
rect 245842 265775 245898 265784
rect 245750 265296 245806 265305
rect 245750 265231 245806 265240
rect 245936 264920 245988 264926
rect 245936 264862 245988 264868
rect 245842 264480 245898 264489
rect 245842 264415 245898 264424
rect 245856 263634 245884 264415
rect 245948 263945 245976 264862
rect 245934 263936 245990 263945
rect 245934 263871 245990 263880
rect 245844 263628 245896 263634
rect 245844 263570 245896 263576
rect 245750 263120 245806 263129
rect 245750 263055 245806 263064
rect 244922 260944 244978 260953
rect 244922 260879 244924 260888
rect 244976 260879 244978 260888
rect 244924 260850 244976 260856
rect 245764 258074 245792 263055
rect 245934 262304 245990 262313
rect 245934 262239 245936 262248
rect 245988 262239 245990 262248
rect 245936 262210 245988 262216
rect 245842 261760 245898 261769
rect 245842 261695 245898 261704
rect 245856 260234 245884 261695
rect 245936 260840 245988 260846
rect 245936 260782 245988 260788
rect 245844 260228 245896 260234
rect 245844 260170 245896 260176
rect 245948 259593 245976 260782
rect 245934 259584 245990 259593
rect 245934 259519 245990 259528
rect 245844 259412 245896 259418
rect 245844 259354 245896 259360
rect 245856 258233 245884 259354
rect 245934 258768 245990 258777
rect 245934 258703 245936 258712
rect 245988 258703 245990 258712
rect 245936 258674 245988 258680
rect 245842 258224 245898 258233
rect 245842 258159 245898 258168
rect 245764 258046 245884 258074
rect 245658 256592 245714 256601
rect 245658 256527 245714 256536
rect 244922 248704 244978 248713
rect 244922 248639 244978 248648
rect 244936 246362 244964 248639
rect 244924 246356 244976 246362
rect 244924 246298 244976 246304
rect 244646 235784 244702 235793
rect 244646 235719 244702 235728
rect 245672 228993 245700 256527
rect 245752 252476 245804 252482
rect 245752 252418 245804 252424
rect 245764 251705 245792 252418
rect 245750 251696 245806 251705
rect 245750 251631 245806 251640
rect 245750 250880 245806 250889
rect 245750 250815 245806 250824
rect 245764 249830 245792 250815
rect 245752 249824 245804 249830
rect 245752 249766 245804 249772
rect 245856 248414 245884 258046
rect 246026 255232 246082 255241
rect 246026 255167 246082 255176
rect 246040 253978 246068 255167
rect 246028 253972 246080 253978
rect 246028 253914 246080 253920
rect 245936 253904 245988 253910
rect 245934 253872 245936 253881
rect 245988 253872 245990 253881
rect 245934 253807 245990 253816
rect 245934 253056 245990 253065
rect 245934 252991 245990 253000
rect 245948 252890 245976 252991
rect 245936 252884 245988 252890
rect 245936 252826 245988 252832
rect 245936 249552 245988 249558
rect 245934 249520 245936 249529
rect 245988 249520 245990 249529
rect 245934 249455 245990 249464
rect 245856 248386 246068 248414
rect 245934 248160 245990 248169
rect 245934 248095 245990 248104
rect 245948 247722 245976 248095
rect 245936 247716 245988 247722
rect 245936 247658 245988 247664
rect 245842 245168 245898 245177
rect 245842 245103 245898 245112
rect 245750 240816 245806 240825
rect 245750 240751 245806 240760
rect 245764 240174 245792 240751
rect 245752 240168 245804 240174
rect 245752 240110 245804 240116
rect 245856 238754 245884 245103
rect 245934 244624 245990 244633
rect 245934 244559 245990 244568
rect 245948 244322 245976 244559
rect 245936 244316 245988 244322
rect 245936 244258 245988 244264
rect 246040 239601 246068 248386
rect 246120 247716 246172 247722
rect 246120 247658 246172 247664
rect 246026 239592 246082 239601
rect 246026 239527 246082 239536
rect 246132 238754 246160 247658
rect 246316 244905 246344 270943
rect 246946 252240 247002 252249
rect 247052 252226 247080 304234
rect 247144 278089 247172 330550
rect 248420 322244 248472 322250
rect 248420 322186 248472 322192
rect 247224 289944 247276 289950
rect 247224 289886 247276 289892
rect 247130 278080 247186 278089
rect 247130 278015 247186 278024
rect 247236 257417 247264 289886
rect 247222 257408 247278 257417
rect 247222 257343 247224 257352
rect 247276 257343 247278 257352
rect 247224 257314 247276 257320
rect 247236 257283 247264 257314
rect 248432 254425 248460 322186
rect 249064 316804 249116 316810
rect 249064 316746 249116 316752
rect 248510 288552 248566 288561
rect 248510 288487 248566 288496
rect 248418 254416 248474 254425
rect 248418 254351 248474 254360
rect 248524 252890 248552 288487
rect 248604 271176 248656 271182
rect 248604 271118 248656 271124
rect 248512 252884 248564 252890
rect 248512 252826 248564 252832
rect 247002 252198 247080 252226
rect 246946 252175 247002 252184
rect 246394 245984 246450 245993
rect 246394 245919 246450 245928
rect 246408 245682 246436 245919
rect 246396 245676 246448 245682
rect 246396 245618 246448 245624
rect 247040 245676 247092 245682
rect 247040 245618 247092 245624
rect 246302 244896 246358 244905
rect 246302 244831 246358 244840
rect 246394 243808 246450 243817
rect 246394 243743 246450 243752
rect 246408 242962 246436 243743
rect 246396 242956 246448 242962
rect 246396 242898 246448 242904
rect 246302 242448 246358 242457
rect 246302 242383 246358 242392
rect 246316 241534 246344 242383
rect 246304 241528 246356 241534
rect 246304 241470 246356 241476
rect 245764 238726 245884 238754
rect 245948 238726 246160 238754
rect 245658 228984 245714 228993
rect 245658 228919 245714 228928
rect 245672 227769 245700 228919
rect 245658 227760 245714 227769
rect 245658 227695 245714 227704
rect 245764 219434 245792 238726
rect 245948 235929 245976 238726
rect 245934 235920 245990 235929
rect 245934 235855 245990 235864
rect 246302 227760 246358 227769
rect 246302 227695 246358 227704
rect 245580 219406 245792 219434
rect 244462 219328 244518 219337
rect 244462 219263 244518 219272
rect 245580 218890 245608 219406
rect 245568 218884 245620 218890
rect 245568 218826 245620 218832
rect 244280 208344 244332 208350
rect 244280 208286 244332 208292
rect 244292 207058 244320 208286
rect 244280 207052 244332 207058
rect 244280 206994 244332 207000
rect 244924 207052 244976 207058
rect 244924 206994 244976 207000
rect 242256 192568 242308 192574
rect 242256 192510 242308 192516
rect 242164 189848 242216 189854
rect 241518 189816 241574 189825
rect 242164 189790 242216 189796
rect 241518 189751 241574 189760
rect 240874 133920 240930 133929
rect 240874 133855 240930 133864
rect 240888 111081 240916 133855
rect 240874 111072 240930 111081
rect 240874 111007 240930 111016
rect 241532 16574 241560 189751
rect 242164 186992 242216 186998
rect 242164 186934 242216 186940
rect 241532 16546 241744 16574
rect 240784 15972 240836 15978
rect 240784 15914 240836 15920
rect 240230 7032 240286 7041
rect 240230 6967 240286 6976
rect 240244 4049 240272 6967
rect 240230 4040 240286 4049
rect 240230 3975 240286 3984
rect 240336 598 240548 626
rect 240336 490 240364 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 462 240364 490
rect 240520 480 240548 598
rect 241716 480 241744 16546
rect 242176 3466 242204 186934
rect 244278 184376 244334 184385
rect 244278 184311 244334 184320
rect 243542 142760 243598 142769
rect 243542 142695 243598 142704
rect 242256 142180 242308 142186
rect 242256 142122 242308 142128
rect 242268 56574 242296 142122
rect 242256 56568 242308 56574
rect 242256 56510 242308 56516
rect 242900 20052 242952 20058
rect 242900 19994 242952 20000
rect 242912 16574 242940 19994
rect 242912 16546 243492 16574
rect 242898 6216 242954 6225
rect 242898 6151 242954 6160
rect 242164 3460 242216 3466
rect 242164 3402 242216 3408
rect 242912 480 242940 6151
rect 243464 3210 243492 16546
rect 243556 3369 243584 142695
rect 243728 122936 243780 122942
rect 243728 122878 243780 122884
rect 243740 113150 243768 122878
rect 243728 113144 243780 113150
rect 243728 113086 243780 113092
rect 243636 111920 243688 111926
rect 243636 111862 243688 111868
rect 243648 87650 243676 111862
rect 243636 87644 243688 87650
rect 243636 87586 243688 87592
rect 243634 82376 243690 82385
rect 243634 82311 243690 82320
rect 243648 40633 243676 82311
rect 243634 40624 243690 40633
rect 243634 40559 243690 40568
rect 244292 16574 244320 184311
rect 244936 176497 244964 206994
rect 245580 184278 245608 218826
rect 245658 200832 245714 200841
rect 245658 200767 245714 200776
rect 245568 184272 245620 184278
rect 245568 184214 245620 184220
rect 244922 176488 244978 176497
rect 244922 176423 244978 176432
rect 245016 136740 245068 136746
rect 245016 136682 245068 136688
rect 244924 111852 244976 111858
rect 244924 111794 244976 111800
rect 244936 55214 244964 111794
rect 245028 91497 245056 136682
rect 245014 91488 245070 91497
rect 245014 91423 245070 91432
rect 245014 80880 245070 80889
rect 245014 80815 245070 80824
rect 245028 66910 245056 80815
rect 245016 66904 245068 66910
rect 245016 66846 245068 66852
rect 244924 55208 244976 55214
rect 244924 55150 244976 55156
rect 245672 16574 245700 200767
rect 246316 95033 246344 227695
rect 247052 213858 247080 245618
rect 247224 242956 247276 242962
rect 247224 242898 247276 242904
rect 247132 241528 247184 241534
rect 247132 241470 247184 241476
rect 247144 228478 247172 241470
rect 247236 234598 247264 242898
rect 248616 238754 248644 271118
rect 249076 270570 249104 316746
rect 249708 281580 249760 281586
rect 249708 281522 249760 281528
rect 249720 279478 249748 281522
rect 249708 279472 249760 279478
rect 249708 279414 249760 279420
rect 249064 270564 249116 270570
rect 249064 270506 249116 270512
rect 249064 252884 249116 252890
rect 249064 252826 249116 252832
rect 248432 238726 248644 238754
rect 248432 236722 248460 238726
rect 248340 236706 248460 236722
rect 248328 236700 248460 236706
rect 248380 236694 248460 236700
rect 248328 236642 248380 236648
rect 247224 234592 247276 234598
rect 247224 234534 247276 234540
rect 247132 228472 247184 228478
rect 247132 228414 247184 228420
rect 247040 213852 247092 213858
rect 247040 213794 247092 213800
rect 248340 210633 248368 236642
rect 249076 229770 249104 252826
rect 249812 249558 249840 349114
rect 249890 317520 249946 317529
rect 249890 317455 249946 317464
rect 249904 276010 249932 317455
rect 249982 298208 250038 298217
rect 249982 298143 250038 298152
rect 249996 278050 250024 298143
rect 250444 285796 250496 285802
rect 250444 285738 250496 285744
rect 249984 278044 250036 278050
rect 249984 277986 250036 277992
rect 249892 276004 249944 276010
rect 249892 275946 249944 275952
rect 249892 273284 249944 273290
rect 249892 273226 249944 273232
rect 249800 249552 249852 249558
rect 249800 249494 249852 249500
rect 249708 240100 249760 240106
rect 249708 240042 249760 240048
rect 249720 235249 249748 240042
rect 249706 235240 249762 235249
rect 249706 235175 249762 235184
rect 249064 229764 249116 229770
rect 249064 229706 249116 229712
rect 249904 216714 249932 273226
rect 250076 266416 250128 266422
rect 250076 266358 250128 266364
rect 249984 253972 250036 253978
rect 249984 253914 250036 253920
rect 249996 220794 250024 253914
rect 250088 240106 250116 266358
rect 250456 261526 250484 285738
rect 251192 264926 251220 362918
rect 251284 272610 251312 367066
rect 262218 364440 262274 364449
rect 262218 364375 262274 364384
rect 252558 356144 252614 356153
rect 252558 356079 252614 356088
rect 251362 347848 251418 347857
rect 251362 347783 251418 347792
rect 251376 282878 251404 347783
rect 251454 295624 251510 295633
rect 251454 295559 251510 295568
rect 251364 282872 251416 282878
rect 251364 282814 251416 282820
rect 251364 278792 251416 278798
rect 251364 278734 251416 278740
rect 251272 272604 251324 272610
rect 251272 272546 251324 272552
rect 251180 264920 251232 264926
rect 251180 264862 251232 264868
rect 251180 262268 251232 262274
rect 251180 262210 251232 262216
rect 250444 261520 250496 261526
rect 250444 261462 250496 261468
rect 250076 240100 250128 240106
rect 250076 240042 250128 240048
rect 249984 220788 250036 220794
rect 249984 220730 250036 220736
rect 251088 220788 251140 220794
rect 251088 220730 251140 220736
rect 251100 220182 251128 220730
rect 251088 220176 251140 220182
rect 251088 220118 251140 220124
rect 249892 216708 249944 216714
rect 249892 216650 249944 216656
rect 250628 216708 250680 216714
rect 250628 216650 250680 216656
rect 248326 210624 248382 210633
rect 248326 210559 248382 210568
rect 247682 207768 247738 207777
rect 247682 207703 247738 207712
rect 246396 153332 246448 153338
rect 246396 153274 246448 153280
rect 246408 131782 246436 153274
rect 246488 146396 246540 146402
rect 246488 146338 246540 146344
rect 246500 134570 246528 146338
rect 246488 134564 246540 134570
rect 246488 134506 246540 134512
rect 246396 131776 246448 131782
rect 246396 131718 246448 131724
rect 246394 119368 246450 119377
rect 246394 119303 246450 119312
rect 246408 95198 246436 119303
rect 246396 95192 246448 95198
rect 246396 95134 246448 95140
rect 246302 95024 246358 95033
rect 246302 94959 246358 94968
rect 246304 93220 246356 93226
rect 246304 93162 246356 93168
rect 244292 16546 245240 16574
rect 245672 16546 245976 16574
rect 243542 3360 243598 3369
rect 243542 3295 243598 3304
rect 243464 3182 244136 3210
rect 244108 480 244136 3182
rect 245212 480 245240 16546
rect 245948 490 245976 16546
rect 246316 15910 246344 93162
rect 246304 15904 246356 15910
rect 246304 15846 246356 15852
rect 247696 6225 247724 207703
rect 250442 204912 250498 204921
rect 250442 204847 250498 204856
rect 247776 194608 247828 194614
rect 247776 194550 247828 194556
rect 247788 169697 247816 194550
rect 249062 179480 249118 179489
rect 249062 179415 249118 179424
rect 248604 173868 248656 173874
rect 248604 173810 248656 173816
rect 248616 172961 248644 173810
rect 248602 172952 248658 172961
rect 248602 172887 248658 172896
rect 248604 172508 248656 172514
rect 248604 172450 248656 172456
rect 248616 171601 248644 172450
rect 248602 171592 248658 171601
rect 248602 171527 248658 171536
rect 247774 169688 247830 169697
rect 247774 169623 247830 169632
rect 248420 167000 248472 167006
rect 248418 166968 248420 166977
rect 248472 166968 248474 166977
rect 248418 166903 248474 166912
rect 248512 166932 248564 166938
rect 248512 166874 248564 166880
rect 248524 166433 248552 166874
rect 248510 166424 248566 166433
rect 248510 166359 248566 166368
rect 248420 165572 248472 165578
rect 248420 165514 248472 165520
rect 248432 165073 248460 165514
rect 248418 165064 248474 165073
rect 248418 164999 248474 165008
rect 248512 164212 248564 164218
rect 248512 164154 248564 164160
rect 248420 164144 248472 164150
rect 248420 164086 248472 164092
rect 248432 163713 248460 164086
rect 248418 163704 248474 163713
rect 248418 163639 248474 163648
rect 248524 163033 248552 164154
rect 248510 163024 248566 163033
rect 248510 162959 248566 162968
rect 248420 162852 248472 162858
rect 248420 162794 248472 162800
rect 248432 162353 248460 162794
rect 248512 162784 248564 162790
rect 248512 162726 248564 162732
rect 248418 162344 248474 162353
rect 248418 162279 248474 162288
rect 248524 161809 248552 162726
rect 248510 161800 248566 161809
rect 248510 161735 248566 161744
rect 248512 161424 248564 161430
rect 248512 161366 248564 161372
rect 248420 161356 248472 161362
rect 248420 161298 248472 161304
rect 248432 161129 248460 161298
rect 248418 161120 248474 161129
rect 248418 161055 248474 161064
rect 248524 160449 248552 161366
rect 248510 160440 248566 160449
rect 248510 160375 248566 160384
rect 248420 160064 248472 160070
rect 248420 160006 248472 160012
rect 248432 159089 248460 160006
rect 248418 159080 248474 159089
rect 248418 159015 248474 159024
rect 248420 158704 248472 158710
rect 248420 158646 248472 158652
rect 248432 158409 248460 158646
rect 248418 158400 248474 158409
rect 248418 158335 248474 158344
rect 249076 157729 249104 179415
rect 249524 176656 249576 176662
rect 249524 176598 249576 176604
rect 249248 175976 249300 175982
rect 249248 175918 249300 175924
rect 249156 169040 249208 169046
rect 249260 169017 249288 175918
rect 249536 175681 249564 176598
rect 249706 176488 249762 176497
rect 249706 176423 249762 176432
rect 249522 175672 249578 175681
rect 249522 175607 249578 175616
rect 249720 175370 249748 176423
rect 249708 175364 249760 175370
rect 249708 175306 249760 175312
rect 249708 175228 249760 175234
rect 249708 175170 249760 175176
rect 249720 175001 249748 175170
rect 249706 174992 249762 175001
rect 249706 174927 249762 174936
rect 249708 173800 249760 173806
rect 249708 173742 249760 173748
rect 249720 173641 249748 173742
rect 249706 173632 249762 173641
rect 249706 173567 249762 173576
rect 249340 172440 249392 172446
rect 249340 172382 249392 172388
rect 249352 172281 249380 172382
rect 249338 172272 249394 172281
rect 249338 172207 249394 172216
rect 249616 171080 249668 171086
rect 249616 171022 249668 171028
rect 249706 171048 249762 171057
rect 249628 170377 249656 171022
rect 249706 170983 249708 170992
rect 249760 170983 249762 170992
rect 249708 170954 249760 170960
rect 249614 170368 249670 170377
rect 249614 170303 249670 170312
rect 249708 169720 249760 169726
rect 249706 169688 249708 169697
rect 249760 169688 249762 169697
rect 249706 169623 249762 169632
rect 249156 168982 249208 168988
rect 249246 169008 249302 169017
rect 249168 159769 249196 168982
rect 249246 168943 249302 168952
rect 249616 168360 249668 168366
rect 249616 168302 249668 168308
rect 249706 168328 249762 168337
rect 249628 167657 249656 168302
rect 249706 168263 249708 168272
rect 249760 168263 249762 168272
rect 249708 168234 249760 168240
rect 249614 167648 249670 167657
rect 249614 167583 249670 167592
rect 249154 159760 249210 159769
rect 249154 159695 249210 159704
rect 249432 158024 249484 158030
rect 249432 157966 249484 157972
rect 249062 157720 249118 157729
rect 249062 157655 249118 157664
rect 249154 154456 249210 154465
rect 249154 154391 249210 154400
rect 249168 153270 249196 154391
rect 249156 153264 249208 153270
rect 249156 153206 249208 153212
rect 248970 153096 249026 153105
rect 248970 153031 249026 153040
rect 248984 151842 249012 153031
rect 249338 152552 249394 152561
rect 249338 152487 249394 152496
rect 248972 151836 249024 151842
rect 248972 151778 249024 151784
rect 249246 151192 249302 151201
rect 249246 151127 249302 151136
rect 248972 151088 249024 151094
rect 248972 151030 249024 151036
rect 248984 149161 249012 151030
rect 249260 149734 249288 151127
rect 249248 149728 249300 149734
rect 249248 149670 249300 149676
rect 248970 149152 249026 149161
rect 248970 149087 249026 149096
rect 249246 147928 249302 147937
rect 249246 147863 249302 147872
rect 249154 147248 249210 147257
rect 249154 147183 249210 147192
rect 249168 146334 249196 147183
rect 249156 146328 249208 146334
rect 249156 146270 249208 146276
rect 249154 144528 249210 144537
rect 249154 144463 249210 144472
rect 249168 143614 249196 144463
rect 249156 143608 249208 143614
rect 249156 143550 249208 143556
rect 249154 140584 249210 140593
rect 249154 140519 249210 140528
rect 248970 139904 249026 139913
rect 248970 139839 249026 139848
rect 247774 132832 247830 132841
rect 247774 132767 247830 132776
rect 247788 112441 247816 132767
rect 248984 132494 249012 139839
rect 249168 139466 249196 140519
rect 249156 139460 249208 139466
rect 249156 139402 249208 139408
rect 249062 139224 249118 139233
rect 249062 139159 249118 139168
rect 249076 135130 249104 139159
rect 249154 138000 249210 138009
rect 249154 137935 249210 137944
rect 249168 136746 249196 137935
rect 249156 136740 249208 136746
rect 249156 136682 249208 136688
rect 249154 136640 249210 136649
rect 249154 136575 249210 136584
rect 249168 135318 249196 136575
rect 249156 135312 249208 135318
rect 249156 135254 249208 135260
rect 249076 135102 249196 135130
rect 248984 132466 249104 132494
rect 248970 124128 249026 124137
rect 248970 124063 249026 124072
rect 248984 122874 249012 124063
rect 248972 122868 249024 122874
rect 248972 122810 249024 122816
rect 248786 122088 248842 122097
rect 248786 122023 248842 122032
rect 248800 121582 248828 122023
rect 248788 121576 248840 121582
rect 248788 121518 248840 121524
rect 248786 119504 248842 119513
rect 248786 119439 248842 119448
rect 248800 118726 248828 119439
rect 248788 118720 248840 118726
rect 248788 118662 248840 118668
rect 248786 118144 248842 118153
rect 248786 118079 248842 118088
rect 248800 117366 248828 118079
rect 248788 117360 248840 117366
rect 248788 117302 248840 117308
rect 248786 116784 248842 116793
rect 248786 116719 248842 116728
rect 248800 116006 248828 116719
rect 248788 116000 248840 116006
rect 248788 115942 248840 115948
rect 247866 115016 247922 115025
rect 247866 114951 247922 114960
rect 247774 112432 247830 112441
rect 247774 112367 247830 112376
rect 247880 95946 247908 114951
rect 248970 112160 249026 112169
rect 248970 112095 249026 112104
rect 248984 111926 249012 112095
rect 248972 111920 249024 111926
rect 248972 111862 249024 111868
rect 248970 110800 249026 110809
rect 248970 110735 249026 110744
rect 248984 110566 249012 110735
rect 248972 110560 249024 110566
rect 248972 110502 249024 110508
rect 248786 106176 248842 106185
rect 248786 106111 248842 106120
rect 248800 104922 248828 106111
rect 248788 104916 248840 104922
rect 248788 104858 248840 104864
rect 248510 103592 248566 103601
rect 248510 103527 248566 103536
rect 248524 101425 248552 103527
rect 248786 101552 248842 101561
rect 248786 101487 248842 101496
rect 248510 101416 248566 101425
rect 248510 101351 248566 101360
rect 247868 95940 247920 95946
rect 247868 95882 247920 95888
rect 248800 94518 248828 101487
rect 249076 100026 249104 132466
rect 249168 108361 249196 135102
rect 249260 133210 249288 147863
rect 249352 138718 249380 152487
rect 249444 148481 249472 157966
rect 249616 157344 249668 157350
rect 249616 157286 249668 157292
rect 249628 156505 249656 157286
rect 249708 157276 249760 157282
rect 249708 157218 249760 157224
rect 249720 157185 249748 157218
rect 249706 157176 249762 157185
rect 249706 157111 249762 157120
rect 249614 156496 249670 156505
rect 249614 156431 249670 156440
rect 249708 155916 249760 155922
rect 249708 155858 249760 155864
rect 249616 155848 249668 155854
rect 249720 155825 249748 155858
rect 249616 155790 249668 155796
rect 249706 155816 249762 155825
rect 249628 155145 249656 155790
rect 249706 155751 249762 155760
rect 249614 155136 249670 155145
rect 249614 155071 249670 155080
rect 249706 153776 249762 153785
rect 249706 153711 249762 153720
rect 249720 153338 249748 153711
rect 249708 153332 249760 153338
rect 249708 153274 249760 153280
rect 249708 151904 249760 151910
rect 249706 151872 249708 151881
rect 249760 151872 249762 151881
rect 249706 151807 249762 151816
rect 249706 150512 249762 150521
rect 249706 150447 249708 150456
rect 249760 150447 249762 150456
rect 249708 150418 249760 150424
rect 249616 150408 249668 150414
rect 249616 150350 249668 150356
rect 249628 149841 249656 150350
rect 249614 149832 249670 149841
rect 249614 149767 249670 149776
rect 249430 148472 249486 148481
rect 249430 148407 249486 148416
rect 249706 146568 249762 146577
rect 249706 146503 249762 146512
rect 249720 146402 249748 146503
rect 249708 146396 249760 146402
rect 249708 146338 249760 146344
rect 249614 145888 249670 145897
rect 249614 145823 249670 145832
rect 249628 142866 249656 145823
rect 249706 145208 249762 145217
rect 249706 145143 249762 145152
rect 249720 144974 249748 145143
rect 249708 144968 249760 144974
rect 249708 144910 249760 144916
rect 249706 143848 249762 143857
rect 249706 143783 249762 143792
rect 249720 143682 249748 143783
rect 249708 143676 249760 143682
rect 249708 143618 249760 143624
rect 249616 142860 249668 142866
rect 249616 142802 249668 142808
rect 249706 142624 249762 142633
rect 249706 142559 249762 142568
rect 249720 142186 249748 142559
rect 249708 142180 249760 142186
rect 249708 142122 249760 142128
rect 249614 141944 249670 141953
rect 249614 141879 249670 141888
rect 249628 140894 249656 141879
rect 249706 141264 249762 141273
rect 249706 141199 249762 141208
rect 249616 140888 249668 140894
rect 249616 140830 249668 140836
rect 249720 140826 249748 141199
rect 249708 140820 249760 140826
rect 249708 140762 249760 140768
rect 249340 138712 249392 138718
rect 249340 138654 249392 138660
rect 249706 138680 249762 138689
rect 249706 138615 249762 138624
rect 249720 138038 249748 138615
rect 249708 138032 249760 138038
rect 249708 137974 249760 137980
rect 249706 137320 249762 137329
rect 249706 137255 249762 137264
rect 249720 136678 249748 137255
rect 249708 136672 249760 136678
rect 249708 136614 249760 136620
rect 249706 135960 249762 135969
rect 249706 135895 249762 135904
rect 249720 135386 249748 135895
rect 249708 135380 249760 135386
rect 249708 135322 249760 135328
rect 249706 134600 249762 134609
rect 249706 134535 249762 134544
rect 249720 133958 249748 134535
rect 249708 133952 249760 133958
rect 249708 133894 249760 133900
rect 249248 133204 249300 133210
rect 249248 133146 249300 133152
rect 249706 132016 249762 132025
rect 249706 131951 249762 131960
rect 249246 131336 249302 131345
rect 249246 131271 249302 131280
rect 249260 120737 249288 131271
rect 249720 131170 249748 131951
rect 249708 131164 249760 131170
rect 249708 131106 249760 131112
rect 249614 130656 249670 130665
rect 249614 130591 249670 130600
rect 249628 129878 249656 130591
rect 249706 129976 249762 129985
rect 249706 129911 249762 129920
rect 249616 129872 249668 129878
rect 249616 129814 249668 129820
rect 249720 129810 249748 129911
rect 249708 129804 249760 129810
rect 249708 129746 249760 129752
rect 249706 129296 249762 129305
rect 249706 129231 249762 129240
rect 249720 128382 249748 129231
rect 249708 128376 249760 128382
rect 249708 128318 249760 128324
rect 249614 128072 249670 128081
rect 249614 128007 249670 128016
rect 249628 127022 249656 128007
rect 249706 127392 249762 127401
rect 249706 127327 249762 127336
rect 249720 127090 249748 127327
rect 249708 127084 249760 127090
rect 249708 127026 249760 127032
rect 249616 127016 249668 127022
rect 249616 126958 249668 126964
rect 249614 126712 249670 126721
rect 249614 126647 249670 126656
rect 249628 125730 249656 126647
rect 249706 126032 249762 126041
rect 249706 125967 249762 125976
rect 249616 125724 249668 125730
rect 249616 125666 249668 125672
rect 249720 125662 249748 125967
rect 249708 125656 249760 125662
rect 249708 125598 249760 125604
rect 249614 125352 249670 125361
rect 249614 125287 249670 125296
rect 249628 124302 249656 125287
rect 249706 124672 249762 124681
rect 249706 124607 249762 124616
rect 249616 124296 249668 124302
rect 249616 124238 249668 124244
rect 249720 124234 249748 124607
rect 249708 124228 249760 124234
rect 249708 124170 249760 124176
rect 249522 123448 249578 123457
rect 249522 123383 249578 123392
rect 249536 122942 249564 123383
rect 249524 122936 249576 122942
rect 249524 122878 249576 122884
rect 249706 122768 249762 122777
rect 249706 122703 249762 122712
rect 249720 121514 249748 122703
rect 249708 121508 249760 121514
rect 249708 121450 249760 121456
rect 249614 121408 249670 121417
rect 249614 121343 249670 121352
rect 249246 120728 249302 120737
rect 249246 120663 249302 120672
rect 249628 120154 249656 121343
rect 249706 120728 249762 120737
rect 249706 120663 249762 120672
rect 249720 120222 249748 120663
rect 249708 120216 249760 120222
rect 249708 120158 249760 120164
rect 249616 120148 249668 120154
rect 249616 120090 249668 120096
rect 249706 120048 249762 120057
rect 249706 119983 249762 119992
rect 249614 118824 249670 118833
rect 249720 118794 249748 119983
rect 249614 118759 249670 118768
rect 249708 118788 249760 118794
rect 249628 117978 249656 118759
rect 249708 118730 249760 118736
rect 249616 117972 249668 117978
rect 249616 117914 249668 117920
rect 249706 114880 249762 114889
rect 249706 114815 249762 114824
rect 249720 114578 249748 114815
rect 249708 114572 249760 114578
rect 249708 114514 249760 114520
rect 249614 114200 249670 114209
rect 249614 114135 249670 114144
rect 249628 113218 249656 114135
rect 249706 113520 249762 113529
rect 249706 113455 249762 113464
rect 249720 113286 249748 113455
rect 249708 113280 249760 113286
rect 249708 113222 249760 113228
rect 249616 113212 249668 113218
rect 249616 113154 249668 113160
rect 249246 112840 249302 112849
rect 249246 112775 249302 112784
rect 249260 111858 249288 112775
rect 249248 111852 249300 111858
rect 249248 111794 249300 111800
rect 249246 111480 249302 111489
rect 249246 111415 249302 111424
rect 249260 110498 249288 111415
rect 249248 110492 249300 110498
rect 249248 110434 249300 110440
rect 249614 110256 249670 110265
rect 249614 110191 249670 110200
rect 249628 109070 249656 110191
rect 249706 109576 249762 109585
rect 249706 109511 249762 109520
rect 249720 109138 249748 109511
rect 249708 109132 249760 109138
rect 249708 109074 249760 109080
rect 249616 109064 249668 109070
rect 249616 109006 249668 109012
rect 249706 108896 249762 108905
rect 249706 108831 249762 108840
rect 249154 108352 249210 108361
rect 249154 108287 249210 108296
rect 249522 108216 249578 108225
rect 249522 108151 249578 108160
rect 249536 107710 249564 108151
rect 249720 107778 249748 108831
rect 249708 107772 249760 107778
rect 249708 107714 249760 107720
rect 249524 107704 249576 107710
rect 249524 107646 249576 107652
rect 249706 107536 249762 107545
rect 249706 107471 249762 107480
rect 249522 106856 249578 106865
rect 249522 106791 249578 106800
rect 249536 106350 249564 106791
rect 249720 106418 249748 107471
rect 249708 106412 249760 106418
rect 249708 106354 249760 106360
rect 249524 106344 249576 106350
rect 249524 106286 249576 106292
rect 249706 105632 249762 105641
rect 249706 105567 249762 105576
rect 249720 104990 249748 105567
rect 249708 104984 249760 104990
rect 249614 104952 249670 104961
rect 249708 104926 249760 104932
rect 249614 104887 249670 104896
rect 249628 104145 249656 104887
rect 249706 104272 249762 104281
rect 249706 104207 249762 104216
rect 249614 104136 249670 104145
rect 249614 104071 249670 104080
rect 249720 103562 249748 104207
rect 249708 103556 249760 103562
rect 249708 103498 249760 103504
rect 249706 102912 249762 102921
rect 249706 102847 249762 102856
rect 249246 102232 249302 102241
rect 249720 102202 249748 102847
rect 249246 102167 249302 102176
rect 249708 102196 249760 102202
rect 249154 101008 249210 101017
rect 249154 100943 249210 100952
rect 249168 100774 249196 100943
rect 249156 100768 249208 100774
rect 249156 100710 249208 100716
rect 249064 100020 249116 100026
rect 249064 99962 249116 99968
rect 249260 98002 249288 102167
rect 249708 102138 249760 102144
rect 249706 100328 249762 100337
rect 249706 100263 249762 100272
rect 249522 99648 249578 99657
rect 249522 99583 249578 99592
rect 249168 97974 249288 98002
rect 248788 94512 248840 94518
rect 248788 94454 248840 94460
rect 249062 89176 249118 89185
rect 249062 89111 249118 89120
rect 248418 71224 248474 71233
rect 248418 71159 248474 71168
rect 247682 6216 247738 6225
rect 247682 6151 247738 6160
rect 247592 3528 247644 3534
rect 247592 3470 247644 3476
rect 246224 598 246436 626
rect 246224 490 246252 598
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 462 246252 490
rect 246408 480 246436 598
rect 247604 480 247632 3470
rect 248432 490 248460 71159
rect 249076 47598 249104 89111
rect 249168 66201 249196 97974
rect 249246 96928 249302 96937
rect 249246 96863 249302 96872
rect 249154 66192 249210 66201
rect 249154 66127 249210 66136
rect 249260 63481 249288 96863
rect 249338 96384 249394 96393
rect 249338 96319 249394 96328
rect 249352 86970 249380 96319
rect 249536 95849 249564 99583
rect 249720 99414 249748 100263
rect 249708 99408 249760 99414
rect 249708 99350 249760 99356
rect 249614 98968 249670 98977
rect 249614 98903 249670 98912
rect 249628 98054 249656 98903
rect 249706 98288 249762 98297
rect 249706 98223 249762 98232
rect 249720 98122 249748 98223
rect 249708 98116 249760 98122
rect 249708 98058 249760 98064
rect 249616 98048 249668 98054
rect 249616 97990 249668 97996
rect 249706 97608 249762 97617
rect 249706 97543 249762 97552
rect 249720 96694 249748 97543
rect 249708 96688 249760 96694
rect 249708 96630 249760 96636
rect 249522 95840 249578 95849
rect 249522 95775 249578 95784
rect 249340 86964 249392 86970
rect 249340 86906 249392 86912
rect 249798 75304 249854 75313
rect 249798 75239 249854 75248
rect 249246 63472 249302 63481
rect 249246 63407 249302 63416
rect 249064 47592 249116 47598
rect 249064 47534 249116 47540
rect 249812 16574 249840 75239
rect 249812 16546 250024 16574
rect 248616 598 248828 626
rect 248616 490 248644 598
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 462 248644 490
rect 248800 480 248828 598
rect 249996 480 250024 16546
rect 250456 3534 250484 204847
rect 250534 178120 250590 178129
rect 250534 178055 250590 178064
rect 250548 49094 250576 178055
rect 250640 177342 250668 216650
rect 251192 205630 251220 262210
rect 251376 224777 251404 278734
rect 251468 259865 251496 295559
rect 251824 272604 251876 272610
rect 251824 272546 251876 272552
rect 251454 259856 251510 259865
rect 251454 259791 251510 259800
rect 251836 232665 251864 272546
rect 252572 240145 252600 356079
rect 255318 355328 255374 355337
rect 255318 355263 255374 355272
rect 252652 336796 252704 336802
rect 252652 336738 252704 336744
rect 252558 240136 252614 240145
rect 252558 240071 252614 240080
rect 252664 238377 252692 336738
rect 254032 309188 254084 309194
rect 254032 309130 254084 309136
rect 252744 296812 252796 296818
rect 252744 296754 252796 296760
rect 252756 260846 252784 296754
rect 253938 290184 253994 290193
rect 253938 290119 253994 290128
rect 253204 287156 253256 287162
rect 253204 287098 253256 287104
rect 253216 271182 253244 287098
rect 253204 271176 253256 271182
rect 253204 271118 253256 271124
rect 252744 260840 252796 260846
rect 252744 260782 252796 260788
rect 253020 260840 253072 260846
rect 253020 260782 253072 260788
rect 253032 260166 253060 260782
rect 253020 260160 253072 260166
rect 253020 260102 253072 260108
rect 252650 238368 252706 238377
rect 252650 238303 252706 238312
rect 252664 237425 252692 238303
rect 252650 237416 252706 237425
rect 252650 237351 252706 237360
rect 253202 237416 253258 237425
rect 253202 237351 253258 237360
rect 251822 232656 251878 232665
rect 251822 232591 251878 232600
rect 251362 224768 251418 224777
rect 251362 224703 251418 224712
rect 251180 205624 251232 205630
rect 251180 205566 251232 205572
rect 252468 205624 252520 205630
rect 252468 205566 252520 205572
rect 252480 204950 252508 205566
rect 252468 204944 252520 204950
rect 252468 204886 252520 204892
rect 251180 191140 251232 191146
rect 251180 191082 251232 191088
rect 250718 190632 250774 190641
rect 250718 190567 250774 190576
rect 250628 177336 250680 177342
rect 250628 177278 250680 177284
rect 250732 172417 250760 190567
rect 250718 172408 250774 172417
rect 250718 172343 250774 172352
rect 250626 128752 250682 128761
rect 250626 128687 250682 128696
rect 250640 93809 250668 128687
rect 250718 98696 250774 98705
rect 250718 98631 250774 98640
rect 250626 93800 250682 93809
rect 250626 93735 250682 93744
rect 250732 92478 250760 98631
rect 250720 92472 250772 92478
rect 250720 92414 250772 92420
rect 250536 49088 250588 49094
rect 250536 49030 250588 49036
rect 251192 3602 251220 191082
rect 251824 187740 251876 187746
rect 251824 187682 251876 187688
rect 251836 173913 251864 187682
rect 253216 178702 253244 237351
rect 253296 231192 253348 231198
rect 253296 231134 253348 231140
rect 253308 180130 253336 231134
rect 253952 220833 253980 290119
rect 254044 258738 254072 309130
rect 254122 298344 254178 298353
rect 254122 298279 254178 298288
rect 254136 266354 254164 298279
rect 254124 266348 254176 266354
rect 254124 266290 254176 266296
rect 254032 258732 254084 258738
rect 254032 258674 254084 258680
rect 254044 254590 254072 258674
rect 254032 254584 254084 254590
rect 254032 254526 254084 254532
rect 255332 252482 255360 355263
rect 259458 350704 259514 350713
rect 259458 350639 259514 350648
rect 258170 326904 258226 326913
rect 258170 326839 258226 326848
rect 255412 312588 255464 312594
rect 255412 312530 255464 312536
rect 255424 266286 255452 312530
rect 256790 312488 256846 312497
rect 256790 312423 256846 312432
rect 256700 299532 256752 299538
rect 256700 299474 256752 299480
rect 255962 293992 256018 294001
rect 255962 293927 256018 293936
rect 255412 266280 255464 266286
rect 255412 266222 255464 266228
rect 255424 265674 255452 266222
rect 255412 265668 255464 265674
rect 255412 265610 255464 265616
rect 255320 252476 255372 252482
rect 255320 252418 255372 252424
rect 255332 251870 255360 252418
rect 255320 251864 255372 251870
rect 255320 251806 255372 251812
rect 255320 249824 255372 249830
rect 255320 249766 255372 249772
rect 253938 220824 253994 220833
rect 253938 220759 253994 220768
rect 254582 220824 254638 220833
rect 254582 220759 254638 220768
rect 254596 186998 254624 220759
rect 255332 212537 255360 249766
rect 255318 212528 255374 212537
rect 255318 212463 255374 212472
rect 254584 186992 254636 186998
rect 254584 186934 254636 186940
rect 253296 180124 253348 180130
rect 253296 180066 253348 180072
rect 253204 178696 253256 178702
rect 253204 178638 253256 178644
rect 255976 176254 256004 293927
rect 256712 253910 256740 299474
rect 256804 268394 256832 312423
rect 258080 305040 258132 305046
rect 258080 304982 258132 304988
rect 256792 268388 256844 268394
rect 256792 268330 256844 268336
rect 256804 262886 256832 268330
rect 256792 262880 256844 262886
rect 256792 262822 256844 262828
rect 258092 259418 258120 304982
rect 258184 281518 258212 326839
rect 258722 282160 258778 282169
rect 258722 282095 258778 282104
rect 258172 281512 258224 281518
rect 258172 281454 258224 281460
rect 258080 259412 258132 259418
rect 258080 259354 258132 259360
rect 256700 253904 256752 253910
rect 256700 253846 256752 253852
rect 256884 253904 256936 253910
rect 256884 253846 256936 253852
rect 256896 253230 256924 253846
rect 256884 253224 256936 253230
rect 256884 253166 256936 253172
rect 258080 244316 258132 244322
rect 258080 244258 258132 244264
rect 256700 240168 256752 240174
rect 256700 240110 256752 240116
rect 256712 215286 256740 240110
rect 256700 215280 256752 215286
rect 256700 215222 256752 215228
rect 256712 214810 256740 215222
rect 256700 214804 256752 214810
rect 256700 214746 256752 214752
rect 257344 214804 257396 214810
rect 257344 214746 257396 214752
rect 256054 212528 256110 212537
rect 256054 212463 256110 212472
rect 256068 185881 256096 212463
rect 256054 185872 256110 185881
rect 256054 185807 256110 185816
rect 257356 177410 257384 214746
rect 258092 206990 258120 244258
rect 258736 240854 258764 282095
rect 259368 281512 259420 281518
rect 259368 281454 259420 281460
rect 259380 280838 259408 281454
rect 259368 280832 259420 280838
rect 259368 280774 259420 280780
rect 259368 259412 259420 259418
rect 259368 259354 259420 259360
rect 259380 258738 259408 259354
rect 259368 258732 259420 258738
rect 259368 258674 259420 258680
rect 258724 240848 258776 240854
rect 258724 240790 258776 240796
rect 259472 238513 259500 350639
rect 261484 302320 261536 302326
rect 261484 302262 261536 302268
rect 259458 238504 259514 238513
rect 259458 238439 259514 238448
rect 259472 237969 259500 238439
rect 259458 237960 259514 237969
rect 259458 237895 259514 237904
rect 260104 235272 260156 235278
rect 260104 235214 260156 235220
rect 258816 232552 258868 232558
rect 258816 232494 258868 232500
rect 258722 223000 258778 223009
rect 258722 222935 258778 222944
rect 258080 206984 258132 206990
rect 258080 206926 258132 206932
rect 258736 189825 258764 222935
rect 258828 217326 258856 232494
rect 260116 220153 260144 235214
rect 260102 220144 260158 220153
rect 260102 220079 260158 220088
rect 258816 217320 258868 217326
rect 258816 217262 258868 217268
rect 260102 217288 260158 217297
rect 260102 217223 260158 217232
rect 258816 210452 258868 210458
rect 258816 210394 258868 210400
rect 258722 189816 258778 189825
rect 258722 189751 258778 189760
rect 258828 184385 258856 210394
rect 259368 206984 259420 206990
rect 259368 206926 259420 206932
rect 259380 206378 259408 206926
rect 259368 206372 259420 206378
rect 259368 206314 259420 206320
rect 258814 184376 258870 184385
rect 258814 184311 258870 184320
rect 258078 180840 258134 180849
rect 258078 180775 258134 180784
rect 258092 179382 258120 180775
rect 258080 179376 258132 179382
rect 258080 179318 258132 179324
rect 259366 178256 259422 178265
rect 259366 178191 259422 178200
rect 259380 177993 259408 178191
rect 259736 178084 259788 178090
rect 259736 178026 259788 178032
rect 259366 177984 259422 177993
rect 259366 177919 259422 177928
rect 257344 177404 257396 177410
rect 257344 177346 257396 177352
rect 259748 176633 259776 178026
rect 260116 177449 260144 217223
rect 260102 177440 260158 177449
rect 260102 177375 260158 177384
rect 259734 176624 259790 176633
rect 259734 176559 259790 176568
rect 255964 176248 256016 176254
rect 255964 176190 256016 176196
rect 261496 175953 261524 302262
rect 261574 287328 261630 287337
rect 261574 287263 261630 287272
rect 261588 182918 261616 287263
rect 262232 267034 262260 364375
rect 317418 320784 317474 320793
rect 317418 320719 317474 320728
rect 295984 320204 296036 320210
rect 295984 320146 296036 320152
rect 284944 318844 284996 318850
rect 284944 318786 284996 318792
rect 269764 314696 269816 314702
rect 269764 314638 269816 314644
rect 268384 313336 268436 313342
rect 268384 313278 268436 313284
rect 262956 303680 263008 303686
rect 262956 303622 263008 303628
rect 262864 288448 262916 288454
rect 262864 288390 262916 288396
rect 262220 267028 262272 267034
rect 262220 266970 262272 266976
rect 262232 264217 262260 266970
rect 262218 264208 262274 264217
rect 262218 264143 262274 264152
rect 262220 263628 262272 263634
rect 262220 263570 262272 263576
rect 262232 216578 262260 263570
rect 262220 216572 262272 216578
rect 262220 216514 262272 216520
rect 262232 215354 262260 216514
rect 262220 215348 262272 215354
rect 262220 215290 262272 215296
rect 261576 182912 261628 182918
rect 261576 182854 261628 182860
rect 262876 180198 262904 288390
rect 262968 287745 262996 303622
rect 267004 300960 267056 300966
rect 267004 300902 267056 300908
rect 265624 291236 265676 291242
rect 265624 291178 265676 291184
rect 264244 288516 264296 288522
rect 264244 288458 264296 288464
rect 262954 287736 263010 287745
rect 262954 287671 263010 287680
rect 263966 287192 264022 287201
rect 263966 287127 264022 287136
rect 262956 215348 263008 215354
rect 262956 215290 263008 215296
rect 262864 180192 262916 180198
rect 262864 180134 262916 180140
rect 262968 176594 262996 215290
rect 262956 176588 263008 176594
rect 262956 176530 263008 176536
rect 262220 176248 262272 176254
rect 262220 176190 262272 176196
rect 261482 175944 261538 175953
rect 261482 175879 261538 175888
rect 262232 175817 262260 176190
rect 262218 175808 262274 175817
rect 262218 175743 262274 175752
rect 251822 173904 251878 173913
rect 251822 173839 251878 173848
rect 263980 139754 264008 287127
rect 264060 203584 264112 203590
rect 264060 203526 264112 203532
rect 264072 164529 264100 203526
rect 264256 179058 264284 288458
rect 264336 195288 264388 195294
rect 264336 195230 264388 195236
rect 264348 190454 264376 195230
rect 264348 190426 264468 190454
rect 264256 179030 264376 179058
rect 264150 177576 264206 177585
rect 264150 177511 264206 177520
rect 264164 174321 264192 177511
rect 264348 177342 264376 179030
rect 264244 177336 264296 177342
rect 264244 177278 264296 177284
rect 264336 177336 264388 177342
rect 264336 177278 264388 177284
rect 264256 174729 264284 177278
rect 264334 176896 264390 176905
rect 264334 176831 264390 176840
rect 264348 175166 264376 176831
rect 264440 176662 264468 190426
rect 265072 188352 265124 188358
rect 265072 188294 265124 188300
rect 264980 177404 265032 177410
rect 264980 177346 265032 177352
rect 264886 177304 264942 177313
rect 264886 177239 264942 177248
rect 264428 176656 264480 176662
rect 264428 176598 264480 176604
rect 264428 175364 264480 175370
rect 264428 175306 264480 175312
rect 264336 175160 264388 175166
rect 264336 175102 264388 175108
rect 264242 174720 264298 174729
rect 264242 174655 264298 174664
rect 264150 174312 264206 174321
rect 264150 174247 264206 174256
rect 264440 171465 264468 175306
rect 264900 175114 264928 177239
rect 264992 175273 265020 177346
rect 264978 175264 265034 175273
rect 264978 175199 265034 175208
rect 264900 175086 265020 175114
rect 264426 171456 264482 171465
rect 264426 171391 264482 171400
rect 264992 165578 265020 175086
rect 264152 165572 264204 165578
rect 264152 165514 264204 165520
rect 264980 165572 265032 165578
rect 264980 165514 265032 165520
rect 264058 164520 264114 164529
rect 264058 164455 264114 164464
rect 264164 146305 264192 165514
rect 265084 160585 265112 188294
rect 265256 184272 265308 184278
rect 265256 184214 265308 184220
rect 265162 175944 265218 175953
rect 265162 175879 265218 175888
rect 265176 164801 265204 175879
rect 265162 164792 265218 164801
rect 265162 164727 265218 164736
rect 265070 160576 265126 160585
rect 265070 160511 265126 160520
rect 265072 159384 265124 159390
rect 265072 159326 265124 159332
rect 265084 154465 265112 159326
rect 265070 154456 265126 154465
rect 265070 154391 265126 154400
rect 264886 153776 264942 153785
rect 264886 153711 264942 153720
rect 264900 150521 264928 153711
rect 264886 150512 264942 150521
rect 264886 150447 264942 150456
rect 265268 149161 265296 184214
rect 265636 176633 265664 291178
rect 266360 279472 266412 279478
rect 266360 279414 266412 279420
rect 266372 193225 266400 279414
rect 266450 232656 266506 232665
rect 266450 232591 266506 232600
rect 266358 193216 266414 193225
rect 266358 193151 266414 193160
rect 265622 176624 265678 176633
rect 265622 176559 265678 176568
rect 266360 173800 266412 173806
rect 266358 173768 266360 173777
rect 266412 173768 266414 173777
rect 266358 173703 266414 173712
rect 266360 172440 266412 172446
rect 266358 172408 266360 172417
rect 266412 172408 266414 172417
rect 266358 172343 266414 172352
rect 266360 171012 266412 171018
rect 266360 170954 266412 170960
rect 266372 170513 266400 170954
rect 266358 170504 266414 170513
rect 266358 170439 266414 170448
rect 266360 169720 266412 169726
rect 266360 169662 266412 169668
rect 266372 169561 266400 169662
rect 266358 169552 266414 169561
rect 266358 169487 266414 169496
rect 266360 169040 266412 169046
rect 266358 169008 266360 169017
rect 266412 169008 266414 169017
rect 266358 168943 266414 168952
rect 266360 168020 266412 168026
rect 266360 167962 266412 167968
rect 266372 167657 266400 167962
rect 266358 167648 266414 167657
rect 266358 167583 266414 167592
rect 266360 166388 266412 166394
rect 266360 166330 266412 166336
rect 266372 166161 266400 166330
rect 266358 166152 266414 166161
rect 266358 166087 266414 166096
rect 265346 165608 265402 165617
rect 265346 165543 265402 165552
rect 266360 165572 266412 165578
rect 265360 152561 265388 165543
rect 266360 165514 266412 165520
rect 266372 165209 266400 165514
rect 266358 165200 266414 165209
rect 266358 165135 266414 165144
rect 266360 164212 266412 164218
rect 266360 164154 266412 164160
rect 266372 163441 266400 164154
rect 266358 163432 266414 163441
rect 266358 163367 266414 163376
rect 266360 162580 266412 162586
rect 266360 162522 266412 162528
rect 266372 161945 266400 162522
rect 266358 161936 266414 161945
rect 266358 161871 266414 161880
rect 266360 161424 266412 161430
rect 266360 161366 266412 161372
rect 266372 160993 266400 161366
rect 266358 160984 266414 160993
rect 266358 160919 266414 160928
rect 266464 160041 266492 232591
rect 267016 220289 267044 300902
rect 267740 287088 267792 287094
rect 267740 287030 267792 287036
rect 267002 220280 267058 220289
rect 267002 220215 267058 220224
rect 266544 220108 266596 220114
rect 266544 220050 266596 220056
rect 266556 171134 266584 220050
rect 266636 173868 266688 173874
rect 266636 173810 266688 173816
rect 266648 172825 266676 173810
rect 266634 172816 266690 172825
rect 266634 172751 266690 172760
rect 266636 172508 266688 172514
rect 266636 172450 266688 172456
rect 266648 171873 266676 172450
rect 266634 171864 266690 171873
rect 266634 171799 266690 171808
rect 266556 171106 266676 171134
rect 266544 162852 266596 162858
rect 266544 162794 266596 162800
rect 266556 161537 266584 162794
rect 266542 161528 266598 161537
rect 266542 161463 266598 161472
rect 266542 160168 266598 160177
rect 266542 160103 266598 160112
rect 266450 160032 266506 160041
rect 266450 159967 266506 159976
rect 266360 158704 266412 158710
rect 266360 158646 266412 158652
rect 266372 158137 266400 158646
rect 266358 158128 266414 158137
rect 266358 158063 266414 158072
rect 266360 157344 266412 157350
rect 266360 157286 266412 157292
rect 266372 157185 266400 157286
rect 266358 157176 266414 157185
rect 266358 157111 266414 157120
rect 266556 156913 266584 160103
rect 266648 157729 266676 171106
rect 266728 171080 266780 171086
rect 266728 171022 266780 171028
rect 266740 169969 266768 171022
rect 266726 169960 266782 169969
rect 266726 169895 266782 169904
rect 267002 169144 267058 169153
rect 267002 169079 267058 169088
rect 266726 167648 266782 167657
rect 266726 167583 266782 167592
rect 266740 162897 266768 167583
rect 266726 162888 266782 162897
rect 266726 162823 266782 162832
rect 266818 159352 266874 159361
rect 266818 159287 266874 159296
rect 266728 158024 266780 158030
rect 266728 157966 266780 157972
rect 266634 157720 266690 157729
rect 266634 157655 266690 157664
rect 266542 156904 266598 156913
rect 266542 156839 266598 156848
rect 266450 156768 266506 156777
rect 266450 156703 266506 156712
rect 266360 155916 266412 155922
rect 266360 155858 266412 155864
rect 266372 155825 266400 155858
rect 266358 155816 266414 155825
rect 266358 155751 266414 155760
rect 266360 155372 266412 155378
rect 266360 155314 266412 155320
rect 265716 153944 265768 153950
rect 266372 153921 266400 155314
rect 266464 155281 266492 156703
rect 266450 155272 266506 155281
rect 266450 155207 266506 155216
rect 265716 153886 265768 153892
rect 266358 153912 266414 153921
rect 265346 152552 265402 152561
rect 265346 152487 265402 152496
rect 265254 149152 265310 149161
rect 265254 149087 265310 149096
rect 264244 146328 264296 146334
rect 264150 146296 264206 146305
rect 264244 146270 264296 146276
rect 264150 146231 264206 146240
rect 264150 139768 264206 139777
rect 263980 139726 264150 139754
rect 264150 139703 264206 139712
rect 263980 138922 264100 138938
rect 263980 138916 264112 138922
rect 263980 138910 264060 138916
rect 263980 127922 264008 138910
rect 264060 138858 264112 138864
rect 264256 137306 264284 146270
rect 264334 145616 264390 145625
rect 264334 145551 264390 145560
rect 264348 141681 264376 145551
rect 265624 143608 265676 143614
rect 265624 143550 265676 143556
rect 265438 142080 265494 142089
rect 265438 142015 265494 142024
rect 264334 141672 264390 141681
rect 264334 141607 264390 141616
rect 265452 140865 265480 142015
rect 265438 140856 265494 140865
rect 265438 140791 265494 140800
rect 264072 137278 264284 137306
rect 265438 137320 265494 137329
rect 264072 132494 264100 137278
rect 265438 137255 265494 137264
rect 265452 136785 265480 137255
rect 265438 136776 265494 136785
rect 265438 136711 265494 136720
rect 264072 132466 264284 132494
rect 264150 127936 264206 127945
rect 263980 127894 264150 127922
rect 264150 127871 264206 127880
rect 264256 122834 264284 132466
rect 264886 131472 264942 131481
rect 264886 131407 264942 131416
rect 264796 127696 264848 127702
rect 264796 127638 264848 127644
rect 264072 122806 264284 122834
rect 264072 105369 264100 122806
rect 264244 120216 264296 120222
rect 264244 120158 264296 120164
rect 264058 105360 264114 105369
rect 264058 105295 264114 105304
rect 251824 101448 251876 101454
rect 251824 101390 251876 101396
rect 251836 89690 251864 101390
rect 264060 98048 264112 98054
rect 264060 97990 264112 97996
rect 252192 97980 252244 97986
rect 252192 97922 252244 97928
rect 252204 96694 252232 97922
rect 264072 96830 264100 97990
rect 264060 96824 264112 96830
rect 264060 96766 264112 96772
rect 252192 96688 252244 96694
rect 252192 96630 252244 96636
rect 264150 96656 264206 96665
rect 264150 96591 264206 96600
rect 257804 96076 257856 96082
rect 257804 96018 257856 96024
rect 257896 96076 257948 96082
rect 257896 96018 257948 96024
rect 261024 96076 261076 96082
rect 261024 96018 261076 96024
rect 257816 95849 257844 96018
rect 257908 95985 257936 96018
rect 261036 95985 261064 96018
rect 257894 95976 257950 95985
rect 261022 95976 261078 95985
rect 257894 95911 257950 95920
rect 258724 95940 258776 95946
rect 261022 95911 261078 95920
rect 262862 95976 262918 95985
rect 262862 95911 262918 95920
rect 258724 95882 258776 95888
rect 257802 95840 257858 95849
rect 257802 95775 257858 95784
rect 257344 94512 257396 94518
rect 257344 94454 257396 94460
rect 254582 90536 254638 90545
rect 254582 90471 254638 90480
rect 251824 89684 251876 89690
rect 251824 89626 251876 89632
rect 253204 86352 253256 86358
rect 253204 86294 253256 86300
rect 251824 65544 251876 65550
rect 251824 65486 251876 65492
rect 251836 36650 251864 65486
rect 253216 40730 253244 86294
rect 253204 40724 253256 40730
rect 253204 40666 253256 40672
rect 251824 36644 251876 36650
rect 251824 36586 251876 36592
rect 251272 21412 251324 21418
rect 251272 21354 251324 21360
rect 251180 3596 251232 3602
rect 251180 3538 251232 3544
rect 250444 3528 250496 3534
rect 251284 3482 251312 21354
rect 254596 8974 254624 90471
rect 255964 83564 256016 83570
rect 255964 83506 256016 83512
rect 255318 69728 255374 69737
rect 255318 69663 255374 69672
rect 255332 16574 255360 69663
rect 255410 63608 255466 63617
rect 255410 63543 255466 63552
rect 255424 61577 255452 63543
rect 255410 61568 255466 61577
rect 255410 61503 255466 61512
rect 255332 16546 255912 16574
rect 254584 8968 254636 8974
rect 254584 8910 254636 8916
rect 254674 6216 254730 6225
rect 254674 6151 254730 6160
rect 252376 3596 252428 3602
rect 252376 3538 252428 3544
rect 250444 3470 250496 3476
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 3538
rect 253478 3496 253534 3505
rect 253478 3431 253534 3440
rect 253492 480 253520 3431
rect 254688 480 254716 6151
rect 255884 480 255912 16546
rect 255976 10334 256004 83506
rect 257356 64297 257384 94454
rect 257342 64288 257398 64297
rect 257342 64223 257398 64232
rect 256698 43480 256754 43489
rect 256698 43415 256754 43424
rect 255964 10328 256016 10334
rect 255964 10270 256016 10276
rect 256712 490 256740 43415
rect 258736 22681 258764 95882
rect 260104 93152 260156 93158
rect 260104 93094 260156 93100
rect 258814 91896 258870 91905
rect 258814 91831 258870 91840
rect 258828 39273 258856 91831
rect 260116 39370 260144 93094
rect 260196 87644 260248 87650
rect 260196 87586 260248 87592
rect 260208 44878 260236 87586
rect 262218 68368 262274 68377
rect 262218 68303 262274 68312
rect 260196 44872 260248 44878
rect 260196 44814 260248 44820
rect 260104 39364 260156 39370
rect 260104 39306 260156 39312
rect 258814 39264 258870 39273
rect 258814 39199 258870 39208
rect 259460 31136 259512 31142
rect 259460 31078 259512 31084
rect 258722 22672 258778 22681
rect 258722 22607 258778 22616
rect 258262 3360 258318 3369
rect 258262 3295 258318 3304
rect 256896 598 257108 626
rect 256896 490 256924 598
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256712 462 256924 490
rect 257080 480 257108 598
rect 258276 480 258304 3295
rect 259472 480 259500 31078
rect 262232 16574 262260 68303
rect 262876 36582 262904 95911
rect 263046 95840 263102 95849
rect 263046 95775 263102 95784
rect 262954 94480 263010 94489
rect 262954 94415 263010 94424
rect 262968 67017 262996 94415
rect 263060 84862 263088 95775
rect 264164 94518 264192 96591
rect 264152 94512 264204 94518
rect 264152 94454 264204 94460
rect 263048 84856 263100 84862
rect 263048 84798 263100 84804
rect 262954 67008 263010 67017
rect 262954 66943 263010 66952
rect 262864 36576 262916 36582
rect 262864 36518 262916 36524
rect 263600 26920 263652 26926
rect 263600 26862 263652 26868
rect 263612 16574 263640 26862
rect 264256 24138 264284 120158
rect 264808 120154 264836 127638
rect 264796 120148 264848 120154
rect 264796 120090 264848 120096
rect 264428 104168 264480 104174
rect 264428 104110 264480 104116
rect 264334 97200 264390 97209
rect 264334 97135 264390 97144
rect 264348 80714 264376 97135
rect 264440 89010 264468 104110
rect 264900 99113 264928 131407
rect 265636 102377 265664 143550
rect 265728 126449 265756 153886
rect 266358 153847 266414 153856
rect 266360 153400 266412 153406
rect 266358 153368 266360 153377
rect 266412 153368 266414 153377
rect 266358 153303 266414 153312
rect 266740 152969 266768 157966
rect 266726 152960 266782 152969
rect 266726 152895 266782 152904
rect 266726 152416 266782 152425
rect 266726 152351 266782 152360
rect 266268 151836 266320 151842
rect 266268 151778 266320 151784
rect 266174 148336 266230 148345
rect 266174 148271 266230 148280
rect 265714 126440 265770 126449
rect 265714 126375 265770 126384
rect 265714 123856 265770 123865
rect 265714 123791 265770 123800
rect 265622 102368 265678 102377
rect 265622 102303 265678 102312
rect 265624 100768 265676 100774
rect 265624 100710 265676 100716
rect 264886 99104 264942 99113
rect 264886 99039 264942 99048
rect 264428 89004 264480 89010
rect 264428 88946 264480 88952
rect 264336 80708 264388 80714
rect 264336 80650 264388 80656
rect 264244 24132 264296 24138
rect 264244 24074 264296 24080
rect 262232 16546 262536 16574
rect 263612 16546 264192 16574
rect 261758 14512 261814 14521
rect 261758 14447 261814 14456
rect 260656 6180 260708 6186
rect 260656 6122 260708 6128
rect 260668 480 260696 6122
rect 261772 480 261800 14447
rect 262508 490 262536 16546
rect 262784 598 262996 626
rect 262784 490 262812 598
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 462 262812 490
rect 262968 480 262996 598
rect 264164 480 264192 16546
rect 264980 15972 265032 15978
rect 264980 15914 265032 15920
rect 264992 490 265020 15914
rect 265636 2106 265664 100710
rect 265728 72593 265756 123791
rect 265898 120592 265954 120601
rect 265898 120527 265954 120536
rect 265808 97776 265860 97782
rect 265808 97718 265860 97724
rect 265714 72584 265770 72593
rect 265714 72519 265770 72528
rect 265820 47666 265848 97718
rect 265912 93226 265940 120527
rect 266188 118017 266216 148271
rect 266280 122834 266308 151778
rect 266360 151632 266412 151638
rect 266358 151600 266360 151609
rect 266412 151600 266414 151609
rect 266358 151535 266414 151544
rect 266450 151328 266506 151337
rect 266450 151263 266506 151272
rect 266360 150408 266412 150414
rect 266360 150350 266412 150356
rect 266372 149705 266400 150350
rect 266358 149696 266414 149705
rect 266358 149631 266414 149640
rect 266464 148209 266492 151263
rect 266740 150113 266768 152351
rect 266832 152017 266860 159287
rect 266818 152008 266874 152017
rect 266818 151943 266874 151952
rect 266726 150104 266782 150113
rect 266726 150039 266782 150048
rect 266542 149696 266598 149705
rect 266542 149631 266598 149640
rect 266556 148753 266584 149631
rect 266542 148744 266598 148753
rect 266542 148679 266598 148688
rect 266450 148200 266506 148209
rect 266450 148135 266506 148144
rect 266360 147620 266412 147626
rect 266360 147562 266412 147568
rect 266372 147257 266400 147562
rect 266358 147248 266414 147257
rect 266358 147183 266414 147192
rect 266360 144900 266412 144906
rect 266360 144842 266412 144848
rect 266372 143993 266400 144842
rect 266358 143984 266414 143993
rect 266358 143919 266414 143928
rect 266360 143540 266412 143546
rect 266360 143482 266412 143488
rect 266372 143041 266400 143482
rect 267016 143449 267044 169079
rect 267646 168056 267702 168065
rect 267752 168042 267780 287030
rect 268396 249082 268424 313278
rect 268384 249076 268436 249082
rect 268384 249018 268436 249024
rect 269120 246356 269172 246362
rect 269120 246298 269172 246304
rect 267832 221536 267884 221542
rect 267832 221478 267884 221484
rect 267702 168014 267780 168042
rect 267646 167991 267702 168000
rect 267844 166818 267872 221478
rect 269132 213926 269160 246298
rect 269120 213920 269172 213926
rect 269118 213888 269120 213897
rect 269172 213888 269174 213897
rect 269118 213823 269174 213832
rect 269396 189848 269448 189854
rect 269396 189790 269448 189796
rect 267922 183016 267978 183025
rect 267922 182951 267978 182960
rect 267660 166790 267872 166818
rect 267660 166705 267688 166790
rect 267646 166696 267702 166705
rect 267646 166631 267702 166640
rect 267738 160712 267794 160721
rect 267738 160647 267794 160656
rect 267646 159624 267702 159633
rect 267752 159610 267780 160647
rect 267702 159582 267780 159610
rect 267646 159559 267702 159568
rect 267096 152516 267148 152522
rect 267096 152458 267148 152464
rect 267002 143440 267058 143449
rect 267002 143375 267058 143384
rect 266358 143032 266414 143041
rect 266358 142967 266414 142976
rect 266452 141432 266504 141438
rect 266452 141374 266504 141380
rect 266360 139392 266412 139398
rect 266360 139334 266412 139340
rect 266372 138825 266400 139334
rect 266358 138816 266414 138825
rect 266358 138751 266414 138760
rect 266360 137284 266412 137290
rect 266360 137226 266412 137232
rect 266372 135969 266400 137226
rect 266358 135960 266414 135969
rect 266358 135895 266414 135904
rect 266360 135652 266412 135658
rect 266360 135594 266412 135600
rect 266372 135425 266400 135594
rect 266358 135416 266414 135425
rect 266358 135351 266414 135360
rect 266360 135244 266412 135250
rect 266360 135186 266412 135192
rect 266372 134473 266400 135186
rect 266464 135017 266492 141374
rect 266450 135008 266506 135017
rect 266450 134943 266506 134952
rect 267002 134600 267058 134609
rect 267002 134535 267058 134544
rect 266358 134464 266414 134473
rect 266358 134399 266414 134408
rect 266360 133884 266412 133890
rect 266360 133826 266412 133832
rect 266372 133113 266400 133826
rect 266358 133104 266414 133113
rect 266358 133039 266414 133048
rect 266360 133000 266412 133006
rect 266360 132942 266412 132948
rect 266372 132569 266400 132942
rect 266358 132560 266414 132569
rect 266358 132495 266414 132504
rect 266452 132456 266504 132462
rect 266452 132398 266504 132404
rect 266360 132388 266412 132394
rect 266360 132330 266412 132336
rect 266372 131617 266400 132330
rect 266358 131608 266414 131617
rect 266358 131543 266414 131552
rect 266464 131209 266492 132398
rect 266450 131200 266506 131209
rect 266450 131135 266506 131144
rect 266452 131096 266504 131102
rect 266358 131064 266414 131073
rect 266452 131038 266504 131044
rect 266358 130999 266414 131008
rect 266372 130257 266400 130999
rect 266358 130248 266414 130257
rect 266358 130183 266414 130192
rect 266464 129849 266492 131038
rect 266544 130960 266596 130966
rect 266544 130902 266596 130908
rect 266450 129840 266506 129849
rect 266450 129775 266506 129784
rect 266360 129736 266412 129742
rect 266360 129678 266412 129684
rect 266372 129305 266400 129678
rect 266358 129296 266414 129305
rect 266358 129231 266414 129240
rect 266556 128897 266584 130902
rect 266542 128888 266598 128897
rect 266542 128823 266598 128832
rect 266542 128208 266598 128217
rect 266542 128143 266598 128152
rect 266360 128036 266412 128042
rect 266360 127978 266412 127984
rect 266372 127401 266400 127978
rect 266452 127628 266504 127634
rect 266452 127570 266504 127576
rect 266358 127392 266414 127401
rect 266358 127327 266414 127336
rect 266360 126948 266412 126954
rect 266360 126890 266412 126896
rect 266372 126041 266400 126890
rect 266358 126032 266414 126041
rect 266358 125967 266414 125976
rect 266360 125588 266412 125594
rect 266360 125530 266412 125536
rect 266372 125497 266400 125530
rect 266358 125488 266414 125497
rect 266358 125423 266414 125432
rect 266464 125089 266492 127570
rect 266450 125080 266506 125089
rect 266450 125015 266506 125024
rect 266556 124137 266584 128143
rect 267016 127702 267044 134535
rect 267108 134065 267136 152458
rect 267188 148436 267240 148442
rect 267188 148378 267240 148384
rect 267094 134056 267150 134065
rect 267094 133991 267150 134000
rect 267200 133521 267228 148378
rect 267646 144936 267702 144945
rect 267936 144922 267964 182951
rect 269304 180124 269356 180130
rect 269304 180066 269356 180072
rect 269212 176656 269264 176662
rect 268014 176624 268070 176633
rect 269212 176598 269264 176604
rect 268014 176559 268070 176568
rect 269120 176588 269172 176594
rect 268028 168026 268056 176559
rect 269120 176530 269172 176536
rect 269132 172446 269160 176530
rect 269120 172440 269172 172446
rect 269120 172382 269172 172388
rect 268016 168020 268068 168026
rect 268016 167962 268068 167968
rect 268660 167136 268712 167142
rect 268660 167078 268712 167084
rect 268568 166320 268620 166326
rect 268568 166262 268620 166268
rect 268382 159080 268438 159089
rect 268382 159015 268438 159024
rect 267702 144894 267964 144922
rect 267646 144871 267702 144880
rect 267738 144800 267794 144809
rect 267738 144735 267794 144744
rect 267752 139398 267780 144735
rect 267740 139392 267792 139398
rect 267740 139334 267792 139340
rect 267186 133512 267242 133521
rect 267186 133447 267242 133456
rect 267096 129668 267148 129674
rect 267096 129610 267148 129616
rect 267004 127696 267056 127702
rect 267004 127638 267056 127644
rect 267004 126268 267056 126274
rect 267004 126210 267056 126216
rect 266912 124908 266964 124914
rect 266912 124850 266964 124856
rect 266542 124128 266598 124137
rect 266542 124063 266598 124072
rect 266634 123448 266690 123457
rect 266634 123383 266690 123392
rect 266360 123208 266412 123214
rect 266358 123176 266360 123185
rect 266412 123176 266414 123185
rect 266358 123111 266414 123120
rect 266280 122806 266492 122834
rect 266360 122732 266412 122738
rect 266360 122674 266412 122680
rect 266372 122641 266400 122674
rect 266358 122632 266414 122641
rect 266358 122567 266414 122576
rect 266360 120012 266412 120018
rect 266360 119954 266412 119960
rect 266372 118969 266400 119954
rect 266358 118960 266414 118969
rect 266358 118895 266414 118904
rect 266360 118652 266412 118658
rect 266360 118594 266412 118600
rect 266372 118153 266400 118594
rect 266358 118144 266414 118153
rect 266358 118079 266414 118088
rect 266174 118008 266230 118017
rect 266174 117943 266230 117952
rect 266360 117292 266412 117298
rect 266360 117234 266412 117240
rect 266268 117224 266320 117230
rect 266268 117166 266320 117172
rect 266174 115016 266230 115025
rect 266174 114951 266230 114960
rect 266188 113174 266216 114951
rect 266280 114753 266308 117166
rect 266372 116521 266400 117234
rect 266358 116512 266414 116521
rect 266358 116447 266414 116456
rect 266360 116204 266412 116210
rect 266360 116146 266412 116152
rect 266372 116113 266400 116146
rect 266358 116104 266414 116113
rect 266358 116039 266414 116048
rect 266360 115864 266412 115870
rect 266360 115806 266412 115812
rect 266372 115569 266400 115806
rect 266358 115560 266414 115569
rect 266358 115495 266414 115504
rect 266266 114744 266322 114753
rect 266266 114679 266322 114688
rect 266360 113688 266412 113694
rect 266358 113656 266360 113665
rect 266412 113656 266414 113665
rect 266358 113591 266414 113600
rect 266188 113146 266308 113174
rect 266280 95946 266308 113146
rect 266360 113076 266412 113082
rect 266360 113018 266412 113024
rect 266372 112713 266400 113018
rect 266358 112704 266414 112713
rect 266358 112639 266414 112648
rect 266464 110809 266492 122806
rect 266544 122800 266596 122806
rect 266544 122742 266596 122748
rect 266556 122233 266584 122742
rect 266542 122224 266598 122233
rect 266542 122159 266598 122168
rect 266648 120737 266676 123383
rect 266924 121689 266952 124850
rect 266910 121680 266966 121689
rect 266910 121615 266966 121624
rect 266634 120728 266690 120737
rect 266634 120663 266690 120672
rect 266636 120148 266688 120154
rect 266636 120090 266688 120096
rect 266544 120080 266596 120086
rect 266544 120022 266596 120028
rect 266556 119377 266584 120022
rect 266542 119368 266598 119377
rect 266542 119303 266598 119312
rect 266544 118584 266596 118590
rect 266544 118526 266596 118532
rect 266556 117473 266584 118526
rect 266542 117464 266598 117473
rect 266542 117399 266598 117408
rect 266648 117230 266676 120090
rect 266636 117224 266688 117230
rect 266636 117166 266688 117172
rect 266544 115932 266596 115938
rect 266544 115874 266596 115880
rect 266556 115161 266584 115874
rect 266542 115152 266598 115161
rect 266542 115087 266598 115096
rect 267016 114617 267044 126210
rect 267108 120329 267136 129610
rect 267094 120320 267150 120329
rect 267094 120255 267150 120264
rect 268396 118425 268424 159015
rect 268476 153876 268528 153882
rect 268476 153818 268528 153824
rect 268488 123214 268516 153818
rect 268580 135658 268608 166262
rect 268672 153406 268700 167078
rect 269224 162586 269252 176598
rect 269316 169046 269344 180066
rect 269304 169040 269356 169046
rect 269304 168982 269356 168988
rect 269408 166394 269436 189790
rect 269776 173369 269804 314638
rect 280160 307896 280212 307902
rect 280160 307838 280212 307844
rect 277400 295452 277452 295458
rect 277400 295394 277452 295400
rect 276662 285832 276718 285841
rect 276662 285767 276718 285776
rect 273260 282940 273312 282946
rect 273260 282882 273312 282888
rect 270776 218816 270828 218822
rect 270776 218758 270828 218764
rect 270592 181552 270644 181558
rect 270592 181494 270644 181500
rect 270500 178084 270552 178090
rect 270500 178026 270552 178032
rect 269762 173360 269818 173369
rect 269762 173295 269818 173304
rect 270512 171018 270540 178026
rect 270500 171012 270552 171018
rect 270500 170954 270552 170960
rect 270038 170368 270094 170377
rect 270038 170303 270094 170312
rect 269948 169040 270000 169046
rect 269948 168982 270000 168988
rect 269396 166388 269448 166394
rect 269396 166330 269448 166336
rect 269212 162580 269264 162586
rect 269212 162522 269264 162528
rect 269212 162172 269264 162178
rect 269212 162114 269264 162120
rect 269224 158545 269252 162114
rect 269764 160132 269816 160138
rect 269764 160074 269816 160080
rect 269210 158536 269266 158545
rect 269210 158471 269266 158480
rect 269118 157448 269174 157457
rect 269118 157383 269174 157392
rect 268660 153400 268712 153406
rect 268660 153342 268712 153348
rect 269132 151638 269160 157383
rect 269120 151632 269172 151638
rect 269120 151574 269172 151580
rect 268660 138032 268712 138038
rect 268660 137974 268712 137980
rect 268568 135652 268620 135658
rect 268568 135594 268620 135600
rect 268672 133006 268700 137974
rect 268752 135924 268804 135930
rect 268752 135866 268804 135872
rect 268660 133000 268712 133006
rect 268660 132942 268712 132948
rect 268764 128042 268792 135866
rect 269776 129674 269804 160074
rect 269856 154624 269908 154630
rect 269856 154566 269908 154572
rect 269764 129668 269816 129674
rect 269764 129610 269816 129616
rect 268752 128036 268804 128042
rect 268752 127978 268804 127984
rect 268568 127492 268620 127498
rect 268568 127434 268620 127440
rect 268476 123208 268528 123214
rect 268476 123150 268528 123156
rect 268382 118416 268438 118425
rect 268382 118351 268438 118360
rect 267186 118144 267242 118153
rect 267186 118079 267242 118088
rect 267094 116512 267150 116521
rect 267094 116447 267150 116456
rect 267002 114608 267058 114617
rect 267002 114543 267058 114552
rect 266544 114504 266596 114510
rect 266544 114446 266596 114452
rect 266556 113257 266584 114446
rect 266542 113248 266598 113257
rect 266542 113183 266598 113192
rect 266544 113144 266596 113150
rect 266544 113086 266596 113092
rect 266556 112305 266584 113086
rect 266542 112296 266598 112305
rect 266542 112231 266598 112240
rect 266542 112024 266598 112033
rect 266542 111959 266598 111968
rect 266450 110800 266506 110809
rect 266450 110735 266506 110744
rect 266452 110424 266504 110430
rect 266452 110366 266504 110372
rect 266360 110356 266412 110362
rect 266360 110298 266412 110304
rect 266372 109449 266400 110298
rect 266464 109857 266492 110366
rect 266450 109848 266506 109857
rect 266450 109783 266506 109792
rect 266358 109440 266414 109449
rect 266358 109375 266414 109384
rect 266360 108996 266412 109002
rect 266360 108938 266412 108944
rect 266372 108497 266400 108938
rect 266358 108488 266414 108497
rect 266358 108423 266414 108432
rect 266556 107953 266584 111959
rect 267004 111172 267056 111178
rect 267004 111114 267056 111120
rect 266542 107944 266598 107953
rect 266542 107879 266598 107888
rect 266360 107636 266412 107642
rect 266360 107578 266412 107584
rect 266372 107137 266400 107578
rect 266452 107568 266504 107574
rect 266452 107510 266504 107516
rect 266358 107128 266414 107137
rect 266358 107063 266414 107072
rect 266464 106593 266492 107510
rect 266450 106584 266506 106593
rect 266450 106519 266506 106528
rect 266360 106276 266412 106282
rect 266360 106218 266412 106224
rect 266372 105641 266400 106218
rect 266358 105632 266414 105641
rect 266358 105567 266414 105576
rect 266360 104100 266412 104106
rect 266360 104042 266412 104048
rect 266372 103737 266400 104042
rect 266358 103728 266414 103737
rect 266358 103663 266414 103672
rect 266452 103488 266504 103494
rect 266452 103430 266504 103436
rect 266360 103420 266412 103426
rect 266360 103362 266412 103368
rect 266372 103329 266400 103362
rect 266358 103320 266414 103329
rect 266358 103255 266414 103264
rect 266464 102785 266492 103430
rect 266450 102776 266506 102785
rect 266450 102711 266506 102720
rect 266450 102096 266506 102105
rect 266360 102060 266412 102066
rect 266450 102031 266506 102040
rect 266360 102002 266412 102008
rect 266372 101833 266400 102002
rect 266358 101824 266414 101833
rect 266358 101759 266414 101768
rect 266464 100881 266492 102031
rect 266634 101416 266690 101425
rect 266634 101351 266690 101360
rect 266450 100872 266506 100881
rect 266450 100807 266506 100816
rect 266360 100700 266412 100706
rect 266360 100642 266412 100648
rect 266372 100473 266400 100642
rect 266452 100632 266504 100638
rect 266452 100574 266504 100580
rect 266358 100464 266414 100473
rect 266358 100399 266414 100408
rect 266464 99929 266492 100574
rect 266542 100056 266598 100065
rect 266542 99991 266598 100000
rect 266450 99920 266506 99929
rect 266450 99855 266506 99864
rect 266452 99340 266504 99346
rect 266452 99282 266504 99288
rect 266358 98696 266414 98705
rect 266358 98631 266414 98640
rect 266372 97617 266400 98631
rect 266464 98025 266492 99282
rect 266556 98569 266584 99991
rect 266648 99521 266676 101351
rect 266634 99512 266690 99521
rect 266634 99447 266690 99456
rect 266542 98560 266598 98569
rect 266542 98495 266598 98504
rect 266450 98016 266506 98025
rect 266450 97951 266506 97960
rect 266358 97608 266414 97617
rect 266358 97543 266414 97552
rect 266910 97336 266966 97345
rect 266910 97271 266966 97280
rect 266924 96665 266952 97271
rect 266910 96656 266966 96665
rect 266910 96591 266966 96600
rect 266450 96248 266506 96257
rect 266450 96183 266506 96192
rect 266268 95940 266320 95946
rect 266268 95882 266320 95888
rect 265900 93220 265952 93226
rect 265900 93162 265952 93168
rect 266464 91798 266492 96183
rect 266452 91792 266504 91798
rect 266452 91734 266504 91740
rect 265808 47660 265860 47666
rect 265808 47602 265860 47608
rect 267016 19990 267044 111114
rect 267108 101561 267136 116447
rect 267200 111353 267228 118079
rect 268580 116210 268608 127434
rect 268934 124808 268990 124817
rect 268934 124743 268990 124752
rect 268658 122224 268714 122233
rect 268658 122159 268714 122168
rect 268568 116204 268620 116210
rect 268568 116146 268620 116152
rect 268566 111888 268622 111897
rect 268566 111823 268622 111832
rect 267186 111344 267242 111353
rect 267186 111279 267242 111288
rect 268476 111104 268528 111110
rect 268476 111046 268528 111052
rect 267278 110256 267334 110265
rect 267278 110191 267334 110200
rect 267188 107704 267240 107710
rect 267188 107646 267240 107652
rect 267094 101552 267150 101561
rect 267094 101487 267150 101496
rect 267096 91792 267148 91798
rect 267096 91734 267148 91740
rect 267108 21486 267136 91734
rect 267200 55894 267228 107646
rect 267292 97782 267320 110191
rect 268382 105224 268438 105233
rect 268382 105159 268438 105168
rect 268290 102504 268346 102513
rect 268290 102439 268346 102448
rect 268304 98054 268332 102439
rect 268292 98048 268344 98054
rect 268292 97990 268344 97996
rect 267280 97776 267332 97782
rect 267280 97718 267332 97724
rect 267646 97064 267702 97073
rect 267702 97022 267780 97050
rect 267646 96999 267702 97008
rect 267752 93838 267780 97022
rect 267740 93832 267792 93838
rect 267740 93774 267792 93780
rect 267752 93537 267780 93774
rect 267738 93528 267794 93537
rect 267738 93463 267794 93472
rect 267188 55888 267240 55894
rect 267188 55830 267240 55836
rect 267740 29640 267792 29646
rect 267740 29582 267792 29588
rect 267096 21480 267148 21486
rect 267096 21422 267148 21428
rect 267004 19984 267056 19990
rect 267004 19926 267056 19932
rect 266542 4856 266598 4865
rect 266542 4791 266598 4800
rect 265624 2100 265676 2106
rect 265624 2042 265676 2048
rect 265176 598 265388 626
rect 265176 490 265204 598
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 462 265204 490
rect 265360 480 265388 598
rect 266556 480 266584 4791
rect 267752 480 267780 29582
rect 268396 16574 268424 105159
rect 268488 24206 268516 111046
rect 268580 46306 268608 111823
rect 268672 110265 268700 122159
rect 268948 110537 268976 124743
rect 269764 120760 269816 120766
rect 269764 120702 269816 120708
rect 269028 116612 269080 116618
rect 269028 116554 269080 116560
rect 268934 110528 268990 110537
rect 268934 110463 268990 110472
rect 268658 110256 268714 110265
rect 268658 110191 268714 110200
rect 269040 102241 269068 116554
rect 269026 102232 269082 102241
rect 269026 102167 269082 102176
rect 268658 86184 268714 86193
rect 268658 86119 268714 86128
rect 268672 65550 268700 86119
rect 268660 65544 268712 65550
rect 268660 65486 268712 65492
rect 268568 46300 268620 46306
rect 268568 46242 268620 46248
rect 269120 33788 269172 33794
rect 269120 33730 269172 33736
rect 268476 24200 268528 24206
rect 268476 24142 268528 24148
rect 268304 16546 268424 16574
rect 268304 7614 268332 16546
rect 268382 13152 268438 13161
rect 268382 13087 268438 13096
rect 268292 7608 268344 7614
rect 268292 7550 268344 7556
rect 268396 490 268424 13087
rect 269132 6914 269160 33730
rect 269776 11830 269804 120702
rect 269868 113694 269896 154566
rect 269960 138038 269988 168982
rect 270052 155378 270080 170303
rect 270604 162858 270632 181494
rect 270682 177440 270738 177449
rect 270682 177375 270738 177384
rect 270696 165753 270724 177375
rect 270788 169726 270816 218758
rect 271970 197976 272026 197985
rect 271970 197911 272026 197920
rect 271878 194168 271934 194177
rect 271878 194103 271934 194112
rect 270776 169720 270828 169726
rect 270776 169662 270828 169668
rect 271420 168428 271472 168434
rect 271420 168370 271472 168376
rect 270682 165744 270738 165753
rect 270682 165679 270738 165688
rect 271328 164892 271380 164898
rect 271328 164834 271380 164840
rect 271236 164144 271288 164150
rect 271236 164086 271288 164092
rect 270592 162852 270644 162858
rect 270592 162794 270644 162800
rect 270590 162752 270646 162761
rect 270590 162687 270646 162696
rect 270604 157350 270632 162687
rect 270592 157344 270644 157350
rect 270592 157286 270644 157292
rect 270040 155372 270092 155378
rect 270040 155314 270092 155320
rect 271142 155272 271198 155281
rect 271142 155207 271198 155216
rect 270040 148368 270092 148374
rect 270040 148310 270092 148316
rect 269948 138032 270000 138038
rect 269948 137974 270000 137980
rect 269948 133204 270000 133210
rect 269948 133146 270000 133152
rect 269856 113688 269908 113694
rect 269856 113630 269908 113636
rect 269960 104106 269988 133146
rect 270052 130966 270080 148310
rect 270040 130960 270092 130966
rect 270040 130902 270092 130908
rect 270040 129056 270092 129062
rect 270040 128998 270092 129004
rect 269948 104100 270000 104106
rect 269948 104042 270000 104048
rect 269854 102232 269910 102241
rect 269854 102167 269910 102176
rect 269764 11824 269816 11830
rect 269764 11766 269816 11772
rect 269868 11762 269896 102167
rect 270052 102066 270080 128998
rect 271156 115870 271184 155207
rect 271248 144906 271276 164086
rect 271236 144900 271288 144906
rect 271236 144842 271288 144848
rect 271236 141500 271288 141506
rect 271236 141442 271288 141448
rect 271144 115864 271196 115870
rect 271144 115806 271196 115812
rect 270222 109168 270278 109177
rect 270222 109103 270278 109112
rect 270130 103864 270186 103873
rect 270130 103799 270186 103808
rect 270040 102060 270092 102066
rect 270040 102002 270092 102008
rect 270144 86358 270172 103799
rect 270236 102377 270264 109103
rect 271248 103426 271276 141442
rect 271340 126954 271368 164834
rect 271432 131102 271460 168370
rect 271892 159390 271920 194103
rect 271984 173806 272012 197911
rect 272064 180192 272116 180198
rect 272064 180134 272116 180140
rect 271972 173800 272024 173806
rect 271972 173742 272024 173748
rect 271970 165608 272026 165617
rect 272076 165578 272104 180134
rect 272156 177336 272208 177342
rect 272156 177278 272208 177284
rect 272168 168609 272196 177278
rect 272706 170096 272762 170105
rect 272706 170031 272762 170040
rect 272154 168600 272210 168609
rect 272154 168535 272210 168544
rect 272616 167068 272668 167074
rect 272616 167010 272668 167016
rect 271970 165543 272026 165552
rect 272064 165572 272116 165578
rect 271880 159384 271932 159390
rect 271880 159326 271932 159332
rect 271984 144809 272012 165543
rect 272064 165514 272116 165520
rect 272522 157584 272578 157593
rect 272522 157519 272578 157528
rect 271970 144800 272026 144809
rect 271970 144735 272026 144744
rect 271420 131096 271472 131102
rect 271420 131038 271472 131044
rect 271786 129976 271842 129985
rect 271786 129911 271842 129920
rect 271328 126948 271380 126954
rect 271328 126890 271380 126896
rect 271418 115832 271474 115841
rect 271418 115767 271474 115776
rect 271326 107672 271382 107681
rect 271326 107607 271382 107616
rect 271236 103420 271288 103426
rect 271236 103362 271288 103368
rect 270222 102368 270278 102377
rect 270222 102303 270278 102312
rect 271234 101008 271290 101017
rect 271234 100943 271290 100952
rect 271144 95260 271196 95266
rect 271144 95202 271196 95208
rect 270132 86352 270184 86358
rect 270132 86294 270184 86300
rect 269856 11756 269908 11762
rect 269856 11698 269908 11704
rect 271156 7682 271184 95202
rect 271248 25566 271276 100943
rect 271340 43518 271368 107607
rect 271432 100881 271460 115767
rect 271512 102196 271564 102202
rect 271512 102138 271564 102144
rect 271418 100872 271474 100881
rect 271418 100807 271474 100816
rect 271524 90545 271552 102138
rect 271800 96529 271828 129911
rect 272536 117298 272564 157519
rect 272628 126993 272656 167010
rect 272720 130665 272748 170031
rect 273272 143546 273300 282882
rect 274640 271176 274692 271182
rect 274640 271118 274692 271124
rect 273352 204944 273404 204950
rect 273352 204886 273404 204892
rect 273364 172514 273392 204886
rect 273444 178696 273496 178702
rect 273444 178638 273496 178644
rect 273352 172508 273404 172514
rect 273352 172450 273404 172456
rect 273456 171134 273484 178638
rect 273904 172576 273956 172582
rect 273904 172518 273956 172524
rect 273364 171106 273484 171134
rect 273364 164150 273392 171106
rect 273442 164248 273498 164257
rect 273442 164183 273498 164192
rect 273352 164144 273404 164150
rect 273352 164086 273404 164092
rect 273456 155961 273484 164183
rect 273442 155952 273498 155961
rect 273442 155887 273498 155896
rect 273260 143540 273312 143546
rect 273260 143482 273312 143488
rect 272800 142180 272852 142186
rect 272800 142122 272852 142128
rect 272706 130656 272762 130665
rect 272706 130591 272762 130600
rect 272812 127498 272840 142122
rect 273916 133890 273944 172518
rect 273994 164656 274050 164665
rect 273994 164591 274050 164600
rect 273904 133884 273956 133890
rect 273904 133826 273956 133832
rect 274008 127634 274036 164591
rect 274652 158710 274680 271118
rect 274732 265668 274784 265674
rect 274732 265610 274784 265616
rect 274744 159361 274772 265610
rect 276020 260228 276072 260234
rect 276020 260170 276072 260176
rect 276032 223582 276060 260170
rect 276020 223576 276072 223582
rect 276018 223544 276020 223553
rect 276072 223544 276074 223553
rect 276018 223479 276074 223488
rect 276032 223453 276060 223479
rect 276020 202224 276072 202230
rect 276020 202166 276072 202172
rect 274822 176896 274878 176905
rect 274822 176831 274878 176840
rect 274836 161430 274864 176831
rect 276032 167142 276060 202166
rect 276112 186992 276164 186998
rect 276112 186934 276164 186940
rect 276020 167136 276072 167142
rect 276020 167078 276072 167084
rect 275282 162072 275338 162081
rect 275282 162007 275338 162016
rect 274824 161424 274876 161430
rect 274824 161366 274876 161372
rect 274730 159352 274786 159361
rect 274730 159287 274786 159296
rect 274640 158704 274692 158710
rect 274640 158646 274692 158652
rect 274088 145716 274140 145722
rect 274088 145658 274140 145664
rect 274100 132394 274128 145658
rect 274180 142860 274232 142866
rect 274180 142802 274232 142808
rect 274088 132388 274140 132394
rect 274088 132330 274140 132336
rect 273996 127628 274048 127634
rect 273996 127570 274048 127576
rect 272800 127492 272852 127498
rect 272800 127434 272852 127440
rect 272614 126984 272670 126993
rect 272614 126919 272670 126928
rect 272708 125656 272760 125662
rect 272708 125598 272760 125604
rect 272524 117292 272576 117298
rect 272524 117234 272576 117240
rect 272616 116000 272668 116006
rect 272616 115942 272668 115948
rect 272628 111178 272656 115942
rect 272616 111172 272668 111178
rect 272616 111114 272668 111120
rect 272522 111072 272578 111081
rect 272522 111007 272578 111016
rect 272062 100872 272118 100881
rect 272062 100807 272118 100816
rect 272076 100774 272104 100807
rect 272064 100768 272116 100774
rect 272064 100710 272116 100716
rect 271786 96520 271842 96529
rect 271786 96455 271842 96464
rect 271510 90536 271566 90545
rect 271510 90471 271566 90480
rect 271328 43512 271380 43518
rect 271328 43454 271380 43460
rect 271328 32496 271380 32502
rect 271328 32438 271380 32444
rect 271236 25560 271288 25566
rect 271236 25502 271288 25508
rect 271144 7676 271196 7682
rect 271144 7618 271196 7624
rect 269132 6886 270080 6914
rect 268672 598 268884 626
rect 268672 490 268700 598
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 462 268700 490
rect 268856 480 268884 598
rect 270052 480 270080 6886
rect 271236 3528 271288 3534
rect 271236 3470 271288 3476
rect 271248 480 271276 3470
rect 271340 3369 271368 32438
rect 271420 28348 271472 28354
rect 271420 28290 271472 28296
rect 271432 3534 271460 28290
rect 272536 13190 272564 111007
rect 272616 99408 272668 99414
rect 272616 99350 272668 99356
rect 272628 42158 272656 99350
rect 272720 69698 272748 125598
rect 274086 124672 274142 124681
rect 274086 124607 274142 124616
rect 272800 123480 272852 123486
rect 272800 123422 272852 123428
rect 272812 100638 272840 123422
rect 273258 117872 273314 117881
rect 273258 117807 273314 117816
rect 273168 113824 273220 113830
rect 273272 113801 273300 117807
rect 273168 113766 273220 113772
rect 273258 113792 273314 113801
rect 273180 104825 273208 113766
rect 273258 113727 273314 113736
rect 273994 109848 274050 109857
rect 273994 109783 274050 109792
rect 273166 104816 273222 104825
rect 273166 104751 273222 104760
rect 272892 104236 272944 104242
rect 272892 104178 272944 104184
rect 272800 100632 272852 100638
rect 272800 100574 272852 100580
rect 272904 87650 272932 104178
rect 273904 98660 273956 98666
rect 273904 98602 273956 98608
rect 272892 87644 272944 87650
rect 272892 87586 272944 87592
rect 272708 69692 272760 69698
rect 272708 69634 272760 69640
rect 273260 50448 273312 50454
rect 273260 50390 273312 50396
rect 272616 42152 272668 42158
rect 272616 42094 272668 42100
rect 272524 13184 272576 13190
rect 272524 13126 272576 13132
rect 271420 3528 271472 3534
rect 271420 3470 271472 3476
rect 272432 3528 272484 3534
rect 272432 3470 272484 3476
rect 271326 3360 271382 3369
rect 271326 3295 271382 3304
rect 272444 480 272472 3470
rect 273272 490 273300 50390
rect 273916 30977 273944 98602
rect 274008 53106 274036 109783
rect 274100 71058 274128 124607
rect 274192 118590 274220 142802
rect 274272 133272 274324 133278
rect 274272 133214 274324 133220
rect 274180 118584 274232 118590
rect 274180 118526 274232 118532
rect 274178 104000 274234 104009
rect 274178 103935 274234 103944
rect 274088 71052 274140 71058
rect 274088 70994 274140 71000
rect 274192 61402 274220 103935
rect 274284 99346 274312 133214
rect 274548 131164 274600 131170
rect 274548 131106 274600 131112
rect 274560 121689 274588 131106
rect 275296 125594 275324 162007
rect 275376 158296 275428 158302
rect 275376 158238 275428 158244
rect 275388 132462 275416 158238
rect 276124 158030 276152 186934
rect 276676 182918 276704 285767
rect 276204 182912 276256 182918
rect 276204 182854 276256 182860
rect 276664 182912 276716 182918
rect 276664 182854 276716 182860
rect 276216 170241 276244 182854
rect 276664 173936 276716 173942
rect 276664 173878 276716 173884
rect 276202 170232 276258 170241
rect 276202 170167 276258 170176
rect 276112 158024 276164 158030
rect 275558 157992 275614 158001
rect 276112 157966 276164 157972
rect 275558 157927 275614 157936
rect 275468 150476 275520 150482
rect 275468 150418 275520 150424
rect 275376 132456 275428 132462
rect 275376 132398 275428 132404
rect 275284 125588 275336 125594
rect 275284 125530 275336 125536
rect 275284 122868 275336 122874
rect 275284 122810 275336 122816
rect 274546 121680 274602 121689
rect 274546 121615 274602 121624
rect 274546 121544 274602 121553
rect 274546 121479 274602 121488
rect 274560 107522 274588 121479
rect 274560 107494 274680 107522
rect 274272 99340 274324 99346
rect 274272 99282 274324 99288
rect 274652 91798 274680 107494
rect 274640 91792 274692 91798
rect 274640 91734 274692 91740
rect 275296 77994 275324 122810
rect 275376 113212 275428 113218
rect 275376 113154 275428 113160
rect 275284 77988 275336 77994
rect 275284 77930 275336 77936
rect 275388 68241 275416 113154
rect 275480 110362 275508 150418
rect 275572 147626 275600 157927
rect 275560 147620 275612 147626
rect 275560 147562 275612 147568
rect 275560 144220 275612 144226
rect 275560 144162 275612 144168
rect 275572 114510 275600 144162
rect 276676 135250 276704 173878
rect 276846 166424 276902 166433
rect 276846 166359 276902 166368
rect 276756 162920 276808 162926
rect 276756 162862 276808 162868
rect 276768 151201 276796 162862
rect 276754 151192 276810 151201
rect 276754 151127 276810 151136
rect 276664 135244 276716 135250
rect 276664 135186 276716 135192
rect 275650 131744 275706 131753
rect 275650 131679 275706 131688
rect 275664 121553 275692 131679
rect 276860 129742 276888 166359
rect 277412 164218 277440 295394
rect 278044 240848 278096 240854
rect 278044 240790 278096 240796
rect 278056 210458 278084 240790
rect 278044 210452 278096 210458
rect 278044 210394 278096 210400
rect 277492 209092 277544 209098
rect 277492 209034 277544 209040
rect 277504 166569 277532 209034
rect 278780 206372 278832 206378
rect 278780 206314 278832 206320
rect 277584 184204 277636 184210
rect 277584 184146 277636 184152
rect 277596 170377 277624 184146
rect 278320 171148 278372 171154
rect 278320 171090 278372 171096
rect 277582 170368 277638 170377
rect 277582 170303 277638 170312
rect 277490 166560 277546 166569
rect 277490 166495 277546 166504
rect 278136 165164 278188 165170
rect 278136 165106 278188 165112
rect 277400 164212 277452 164218
rect 277400 164154 277452 164160
rect 278042 160440 278098 160449
rect 278042 160375 278098 160384
rect 277032 158024 277084 158030
rect 277032 157966 277084 157972
rect 276940 146940 276992 146946
rect 276940 146882 276992 146888
rect 276848 129736 276900 129742
rect 276848 129678 276900 129684
rect 276756 128376 276808 128382
rect 276756 128318 276808 128324
rect 275650 121544 275706 121553
rect 275650 121479 275706 121488
rect 276662 117464 276718 117473
rect 276662 117399 276718 117408
rect 275560 114504 275612 114510
rect 275560 114446 275612 114452
rect 275558 110800 275614 110809
rect 275558 110735 275614 110744
rect 275468 110356 275520 110362
rect 275468 110298 275520 110304
rect 275572 84930 275600 110735
rect 275560 84924 275612 84930
rect 275560 84866 275612 84872
rect 275374 68232 275430 68241
rect 275374 68167 275430 68176
rect 274180 61396 274232 61402
rect 274180 61338 274232 61344
rect 273996 53100 274048 53106
rect 273996 53042 274048 53048
rect 276020 39432 276072 39438
rect 276020 39374 276072 39380
rect 273902 30968 273958 30977
rect 273902 30903 273958 30912
rect 274822 3360 274878 3369
rect 274822 3295 274878 3304
rect 273456 598 273668 626
rect 273456 490 273484 598
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 462 273484 490
rect 273640 480 273668 598
rect 274836 480 274864 3295
rect 276032 480 276060 39374
rect 276676 22778 276704 117399
rect 276768 49026 276796 128318
rect 276952 107574 276980 146882
rect 277044 145722 277072 157966
rect 277032 145716 277084 145722
rect 277032 145658 277084 145664
rect 277124 137352 277176 137358
rect 277124 137294 277176 137300
rect 277032 129804 277084 129810
rect 277032 129746 277084 129752
rect 277044 115025 277072 129746
rect 277136 126274 277164 137294
rect 277124 126268 277176 126274
rect 277124 126210 277176 126216
rect 277306 126032 277362 126041
rect 277306 125967 277362 125976
rect 277320 118017 277348 125967
rect 278056 120057 278084 160375
rect 278148 152425 278176 165106
rect 278226 153912 278282 153921
rect 278226 153847 278282 153856
rect 278134 152416 278190 152425
rect 278134 152351 278190 152360
rect 278136 150544 278188 150550
rect 278136 150486 278188 150492
rect 278042 120048 278098 120057
rect 278042 119983 278098 119992
rect 277306 118008 277362 118017
rect 277306 117943 277362 117952
rect 277030 115016 277086 115025
rect 277030 114951 277086 114960
rect 277030 113792 277086 113801
rect 277030 113727 277086 113736
rect 276940 107568 276992 107574
rect 276940 107510 276992 107516
rect 276846 106312 276902 106321
rect 276846 106247 276902 106256
rect 276860 58585 276888 106247
rect 277044 98841 277072 113727
rect 278044 110492 278096 110498
rect 278044 110434 278096 110440
rect 277030 98832 277086 98841
rect 277030 98767 277086 98776
rect 276940 98728 276992 98734
rect 276940 98670 276992 98676
rect 276952 83570 276980 98670
rect 276940 83564 276992 83570
rect 276940 83506 276992 83512
rect 276846 58576 276902 58585
rect 276846 58511 276902 58520
rect 276756 49020 276808 49026
rect 276756 48962 276808 48968
rect 278056 22846 278084 110434
rect 278148 110430 278176 150486
rect 278240 113082 278268 153847
rect 278332 132433 278360 171090
rect 278792 167385 278820 206314
rect 278870 187096 278926 187105
rect 278870 187031 278926 187040
rect 278778 167376 278834 167385
rect 278778 167311 278834 167320
rect 278778 157448 278834 157457
rect 278778 157383 278834 157392
rect 278792 150414 278820 157383
rect 278884 156913 278912 187031
rect 279514 172816 279570 172825
rect 279514 172751 279570 172760
rect 279424 158772 279476 158778
rect 279424 158714 279476 158720
rect 278870 156904 278926 156913
rect 278870 156839 278926 156848
rect 278780 150408 278832 150414
rect 278780 150350 278832 150356
rect 278318 132424 278374 132433
rect 278318 132359 278374 132368
rect 278320 130416 278372 130422
rect 278320 130358 278372 130364
rect 278228 113076 278280 113082
rect 278228 113018 278280 113024
rect 278136 110424 278188 110430
rect 278136 110366 278188 110372
rect 278228 109064 278280 109070
rect 278228 109006 278280 109012
rect 278136 102264 278188 102270
rect 278136 102206 278188 102212
rect 278148 86290 278176 102206
rect 278136 86284 278188 86290
rect 278136 86226 278188 86232
rect 278240 75206 278268 109006
rect 278332 95266 278360 130358
rect 279436 118658 279464 158714
rect 279528 148442 279556 172751
rect 280172 171086 280200 307838
rect 280802 301064 280858 301073
rect 280802 300999 280858 301008
rect 280252 270564 280304 270570
rect 280252 270506 280304 270512
rect 280264 173874 280292 270506
rect 280816 244934 280844 300999
rect 282920 283892 282972 283898
rect 282920 283834 282972 283840
rect 282184 276684 282236 276690
rect 282184 276626 282236 276632
rect 280804 244928 280856 244934
rect 280804 244870 280856 244876
rect 280342 232520 280398 232529
rect 280342 232455 280398 232464
rect 280252 173868 280304 173874
rect 280252 173810 280304 173816
rect 280160 171080 280212 171086
rect 280160 171022 280212 171028
rect 279608 169788 279660 169794
rect 279608 169730 279660 169736
rect 279620 158302 279648 169730
rect 279608 158296 279660 158302
rect 279608 158238 279660 158244
rect 279608 155984 279660 155990
rect 279608 155926 279660 155932
rect 279516 148436 279568 148442
rect 279516 148378 279568 148384
rect 279620 142186 279648 155926
rect 280356 155922 280384 232455
rect 282092 221468 282144 221474
rect 282092 221410 282144 221416
rect 281540 220176 281592 220182
rect 281540 220118 281592 220124
rect 280896 171216 280948 171222
rect 280896 171158 280948 171164
rect 280804 167136 280856 167142
rect 280804 167078 280856 167084
rect 280344 155916 280396 155922
rect 280344 155858 280396 155864
rect 279700 147688 279752 147694
rect 279700 147630 279752 147636
rect 279608 142180 279660 142186
rect 279608 142122 279660 142128
rect 279608 138032 279660 138038
rect 279608 137974 279660 137980
rect 279424 118652 279476 118658
rect 279424 118594 279476 118600
rect 278504 117496 278556 117502
rect 278504 117438 278556 117444
rect 278412 111852 278464 111858
rect 278412 111794 278464 111800
rect 278424 102202 278452 111794
rect 278516 111110 278544 117438
rect 279516 117360 279568 117366
rect 279516 117302 279568 117308
rect 279422 115832 279478 115841
rect 279422 115767 279478 115776
rect 278504 111104 278556 111110
rect 278504 111046 278556 111052
rect 278412 102196 278464 102202
rect 278412 102138 278464 102144
rect 278320 95260 278372 95266
rect 278320 95202 278372 95208
rect 278228 75200 278280 75206
rect 278228 75142 278280 75148
rect 278778 25528 278834 25537
rect 278778 25463 278834 25472
rect 278044 22840 278096 22846
rect 278044 22782 278096 22788
rect 276664 22772 276716 22778
rect 276664 22714 276716 22720
rect 276110 19952 276166 19961
rect 276110 19887 276166 19896
rect 276124 16574 276152 19887
rect 278792 16574 278820 25463
rect 276124 16546 276704 16574
rect 278792 16546 279096 16574
rect 276676 490 276704 16546
rect 278318 4040 278374 4049
rect 278318 3975 278374 3984
rect 276952 598 277164 626
rect 276952 490 276980 598
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 462 276980 490
rect 277136 480 277164 598
rect 278332 480 278360 3975
rect 279068 490 279096 16546
rect 279436 6254 279464 115767
rect 279528 28286 279556 117302
rect 279620 55865 279648 137974
rect 279712 107642 279740 147630
rect 280066 147112 280122 147121
rect 280066 147047 280122 147056
rect 279790 143848 279846 143857
rect 279790 143783 279846 143792
rect 279804 116521 279832 143783
rect 280080 143585 280108 147047
rect 280066 143576 280122 143585
rect 280066 143511 280122 143520
rect 280816 138718 280844 167078
rect 280908 158030 280936 171158
rect 281552 167657 281580 220118
rect 282104 220114 282132 221410
rect 282092 220108 282144 220114
rect 282092 220050 282144 220056
rect 281632 208412 281684 208418
rect 281632 208354 281684 208360
rect 281538 167648 281594 167657
rect 281538 167583 281594 167592
rect 281644 165170 281672 208354
rect 282196 177342 282224 276626
rect 282184 177336 282236 177342
rect 282184 177278 282236 177284
rect 282276 172644 282328 172650
rect 282276 172586 282328 172592
rect 282182 168464 282238 168473
rect 282182 168399 282238 168408
rect 281632 165164 281684 165170
rect 281632 165106 281684 165112
rect 281080 158840 281132 158846
rect 281080 158782 281132 158788
rect 280896 158024 280948 158030
rect 280896 157966 280948 157972
rect 280988 149116 281040 149122
rect 280988 149058 281040 149064
rect 280804 138712 280856 138718
rect 280804 138654 280856 138660
rect 280896 138100 280948 138106
rect 280896 138042 280948 138048
rect 280804 125724 280856 125730
rect 280804 125666 280856 125672
rect 279790 116512 279846 116521
rect 279790 116447 279846 116456
rect 279700 107636 279752 107642
rect 279700 107578 279752 107584
rect 279700 100768 279752 100774
rect 279700 100710 279752 100716
rect 279712 84833 279740 100710
rect 279698 84824 279754 84833
rect 279698 84759 279754 84768
rect 279606 55856 279662 55865
rect 279606 55791 279662 55800
rect 280816 32434 280844 125666
rect 280908 87553 280936 138042
rect 281000 109002 281028 149058
rect 281092 120018 281120 158782
rect 281172 155168 281224 155174
rect 281172 155110 281224 155116
rect 281184 137358 281212 155110
rect 281172 137352 281224 137358
rect 281172 137294 281224 137300
rect 282196 128353 282224 168399
rect 282288 152522 282316 172586
rect 282932 166297 282960 283834
rect 284956 235278 284984 318786
rect 294602 314800 294658 314809
rect 294602 314735 294658 314744
rect 288440 313404 288492 313410
rect 288440 313346 288492 313352
rect 286416 306468 286468 306474
rect 286416 306410 286468 306416
rect 286324 280832 286376 280838
rect 286324 280774 286376 280780
rect 284944 235272 284996 235278
rect 284944 235214 284996 235220
rect 283010 222320 283066 222329
rect 283010 222255 283066 222264
rect 282918 166288 282974 166297
rect 282918 166223 282974 166232
rect 282552 164484 282604 164490
rect 282552 164426 282604 164432
rect 282460 161560 282512 161566
rect 282460 161502 282512 161508
rect 282276 152516 282328 152522
rect 282276 152458 282328 152464
rect 282274 148744 282330 148753
rect 282274 148679 282330 148688
rect 282182 128344 282238 128353
rect 282182 128279 282238 128288
rect 281080 120012 281132 120018
rect 281080 119954 281132 119960
rect 282182 115968 282238 115977
rect 282182 115903 282238 115912
rect 281446 113384 281502 113393
rect 281446 113319 281502 113328
rect 280988 108996 281040 109002
rect 280988 108938 281040 108944
rect 280988 106412 281040 106418
rect 280988 106354 281040 106360
rect 280894 87544 280950 87553
rect 280894 87479 280950 87488
rect 281000 57254 281028 106354
rect 281460 106185 281488 113319
rect 281446 106176 281502 106185
rect 281446 106111 281502 106120
rect 281080 104984 281132 104990
rect 281080 104926 281132 104932
rect 281092 60081 281120 104926
rect 281540 102332 281592 102338
rect 281540 102274 281592 102280
rect 281552 98666 281580 102274
rect 281540 98660 281592 98666
rect 281540 98602 281592 98608
rect 281078 60072 281134 60081
rect 281078 60007 281134 60016
rect 280988 57248 281040 57254
rect 280988 57190 281040 57196
rect 282196 46209 282224 115903
rect 282288 106282 282316 148679
rect 282368 142180 282420 142186
rect 282368 142122 282420 142128
rect 282276 106276 282328 106282
rect 282276 106218 282328 106224
rect 282274 103592 282330 103601
rect 282274 103527 282330 103536
rect 282182 46200 282238 46209
rect 282182 46135 282238 46144
rect 282288 37942 282316 103527
rect 282380 100706 282408 142122
rect 282472 122738 282500 161502
rect 282564 142769 282592 164426
rect 283024 158001 283052 222255
rect 286336 215966 286364 280774
rect 286428 243574 286456 306410
rect 287702 302424 287758 302433
rect 287702 302359 287758 302368
rect 287716 250510 287744 302359
rect 287704 250504 287756 250510
rect 287704 250446 287756 250452
rect 286416 243568 286468 243574
rect 286416 243510 286468 243516
rect 286508 242956 286560 242962
rect 286508 242898 286560 242904
rect 286324 215960 286376 215966
rect 286324 215902 286376 215908
rect 284300 194608 284352 194614
rect 284300 194550 284352 194556
rect 283104 187740 283156 187746
rect 283104 187682 283156 187688
rect 283116 162178 283144 187682
rect 283748 174072 283800 174078
rect 283748 174014 283800 174020
rect 283656 165640 283708 165646
rect 283656 165582 283708 165588
rect 283104 162172 283156 162178
rect 283104 162114 283156 162120
rect 283010 157992 283066 158001
rect 283010 157927 283066 157936
rect 283564 156052 283616 156058
rect 283564 155994 283616 156000
rect 282550 142760 282606 142769
rect 282550 142695 282606 142704
rect 282828 124228 282880 124234
rect 282828 124170 282880 124176
rect 282460 122732 282512 122738
rect 282460 122674 282512 122680
rect 282458 122224 282514 122233
rect 282458 122159 282514 122168
rect 282472 113830 282500 122159
rect 282840 117502 282868 124170
rect 282828 117496 282880 117502
rect 282828 117438 282880 117444
rect 283576 117201 283604 155994
rect 283668 153950 283696 165582
rect 283656 153944 283708 153950
rect 283656 153886 283708 153892
rect 283656 151904 283708 151910
rect 283656 151846 283708 151852
rect 283562 117192 283618 117201
rect 283562 117127 283618 117136
rect 282460 113824 282512 113830
rect 282460 113766 282512 113772
rect 282920 110560 282972 110566
rect 282920 110502 282972 110508
rect 282458 109032 282514 109041
rect 282458 108967 282514 108976
rect 282472 102270 282500 108967
rect 282932 104242 282960 110502
rect 283668 110401 283696 151846
rect 283760 137290 283788 174014
rect 284312 160721 284340 194550
rect 285680 193928 285732 193934
rect 285680 193870 285732 193876
rect 285218 174448 285274 174457
rect 285218 174383 285274 174392
rect 284942 168600 284998 168609
rect 284942 168535 284998 168544
rect 284298 160712 284354 160721
rect 284298 160647 284354 160656
rect 283840 157956 283892 157962
rect 283840 157898 283892 157904
rect 283852 138689 283880 157898
rect 284956 148374 284984 168535
rect 285128 161492 285180 161498
rect 285128 161434 285180 161440
rect 285034 155952 285090 155961
rect 285034 155887 285090 155896
rect 284944 148368 284996 148374
rect 284944 148310 284996 148316
rect 284944 144968 284996 144974
rect 284944 144910 284996 144916
rect 284300 139868 284352 139874
rect 284300 139810 284352 139816
rect 283838 138680 283894 138689
rect 283838 138615 283894 138624
rect 283748 137284 283800 137290
rect 283748 137226 283800 137232
rect 283840 136672 283892 136678
rect 283840 136614 283892 136620
rect 283852 122097 283880 136614
rect 284312 133210 284340 139810
rect 284300 133204 284352 133210
rect 284300 133146 284352 133152
rect 283932 127016 283984 127022
rect 283932 126958 283984 126964
rect 283838 122088 283894 122097
rect 283838 122023 283894 122032
rect 283748 121508 283800 121514
rect 283748 121450 283800 121456
rect 283654 110392 283710 110401
rect 283654 110327 283710 110336
rect 283564 109132 283616 109138
rect 283564 109074 283616 109080
rect 282920 104236 282972 104242
rect 282920 104178 282972 104184
rect 282918 102504 282974 102513
rect 282918 102439 282974 102448
rect 282460 102264 282512 102270
rect 282460 102206 282512 102212
rect 282368 100700 282420 100706
rect 282368 100642 282420 100648
rect 282932 98734 282960 102439
rect 282920 98728 282972 98734
rect 282920 98670 282972 98676
rect 282458 98288 282514 98297
rect 282458 98223 282514 98232
rect 282368 98116 282420 98122
rect 282368 98058 282420 98064
rect 282380 46238 282408 98058
rect 282472 91905 282500 98223
rect 282458 91896 282514 91905
rect 282458 91831 282514 91840
rect 283576 51746 283604 109074
rect 283760 104174 283788 121450
rect 283944 113801 283972 126958
rect 283930 113792 283986 113801
rect 283930 113727 283986 113736
rect 284024 113280 284076 113286
rect 284024 113222 284076 113228
rect 284036 105505 284064 113222
rect 284298 112704 284354 112713
rect 284298 112639 284354 112648
rect 284312 109721 284340 112639
rect 284298 109712 284354 109721
rect 284298 109647 284354 109656
rect 284022 105496 284078 105505
rect 284022 105431 284078 105440
rect 283840 104916 283892 104922
rect 283840 104858 283892 104864
rect 283748 104168 283800 104174
rect 283748 104110 283800 104116
rect 283656 98184 283708 98190
rect 283656 98126 283708 98132
rect 283564 51740 283616 51746
rect 283564 51682 283616 51688
rect 282368 46232 282420 46238
rect 282368 46174 282420 46180
rect 283668 43450 283696 98126
rect 283852 93158 283880 104858
rect 284956 103494 284984 144910
rect 285048 115938 285076 155887
rect 285140 124914 285168 161434
rect 285232 141438 285260 174383
rect 285692 162761 285720 193870
rect 285770 184376 285826 184385
rect 285770 184311 285826 184320
rect 285678 162752 285734 162761
rect 285678 162687 285734 162696
rect 285784 156777 285812 184311
rect 286520 184210 286548 242898
rect 287702 238232 287758 238241
rect 287702 238167 287758 238176
rect 286508 184204 286560 184210
rect 286508 184146 286560 184152
rect 287610 173632 287666 173641
rect 287610 173567 287666 173576
rect 287624 172650 287652 173567
rect 287612 172644 287664 172650
rect 287612 172586 287664 172592
rect 287242 172272 287298 172281
rect 287242 172207 287298 172216
rect 286414 170096 286470 170105
rect 286414 170031 286470 170040
rect 286322 162888 286378 162897
rect 286322 162823 286378 162832
rect 285770 156768 285826 156777
rect 285770 156703 285826 156712
rect 285220 141432 285272 141438
rect 285220 141374 285272 141380
rect 285220 132524 285272 132530
rect 285220 132466 285272 132472
rect 285128 124908 285180 124914
rect 285128 124850 285180 124856
rect 285128 118720 285180 118726
rect 285128 118662 285180 118668
rect 285036 115932 285088 115938
rect 285036 115874 285088 115880
rect 285140 111858 285168 118662
rect 285232 116618 285260 132466
rect 286336 122806 286364 162823
rect 286428 131073 286456 170031
rect 287256 169046 287284 172207
rect 287244 169040 287296 169046
rect 287244 168982 287296 168988
rect 287426 164520 287482 164529
rect 287426 164455 287482 164464
rect 287440 163441 287468 164455
rect 287426 163432 287482 163441
rect 287426 163367 287482 163376
rect 287150 161936 287206 161945
rect 287150 161871 287206 161880
rect 286506 160304 286562 160313
rect 286506 160239 286562 160248
rect 286414 131064 286470 131073
rect 286414 130999 286470 131008
rect 286414 123312 286470 123321
rect 286414 123247 286470 123256
rect 286324 122800 286376 122806
rect 286324 122742 286376 122748
rect 285220 116612 285272 116618
rect 285220 116554 285272 116560
rect 285588 116068 285640 116074
rect 285588 116010 285640 116016
rect 285220 114572 285272 114578
rect 285220 114514 285272 114520
rect 285128 111852 285180 111858
rect 285128 111794 285180 111800
rect 285128 106480 285180 106486
rect 285128 106422 285180 106428
rect 284944 103488 284996 103494
rect 284944 103430 284996 103436
rect 285036 102264 285088 102270
rect 285036 102206 285088 102212
rect 284300 102196 284352 102202
rect 284300 102138 284352 102144
rect 284116 99476 284168 99482
rect 284116 99418 284168 99424
rect 283930 98696 283986 98705
rect 283930 98631 283986 98640
rect 283840 93152 283892 93158
rect 283840 93094 283892 93100
rect 283944 59945 283972 98631
rect 284128 98025 284156 99418
rect 284114 98016 284170 98025
rect 284114 97951 284170 97960
rect 284312 94489 284340 102138
rect 284944 100836 284996 100842
rect 284944 100778 284996 100784
rect 284298 94480 284354 94489
rect 284298 94415 284354 94424
rect 284956 82113 284984 100778
rect 284942 82104 284998 82113
rect 284942 82039 284998 82048
rect 284298 66872 284354 66881
rect 284298 66807 284354 66816
rect 283930 59936 283986 59945
rect 283930 59871 283986 59880
rect 283656 43444 283708 43450
rect 283656 43386 283708 43392
rect 282276 37936 282328 37942
rect 282276 37878 282328 37884
rect 280804 32428 280856 32434
rect 280804 32370 280856 32376
rect 279516 28280 279568 28286
rect 279516 28222 279568 28228
rect 281540 18692 281592 18698
rect 281540 18634 281592 18640
rect 280802 10296 280858 10305
rect 280802 10231 280858 10240
rect 279424 6248 279476 6254
rect 279424 6190 279476 6196
rect 280710 3360 280766 3369
rect 280710 3295 280766 3304
rect 279344 598 279556 626
rect 279344 490 279372 598
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 462 279372 490
rect 279528 480 279556 598
rect 280724 480 280752 3295
rect 280816 3126 280844 10231
rect 280804 3120 280856 3126
rect 280804 3062 280856 3068
rect 281552 490 281580 18634
rect 283104 3120 283156 3126
rect 283104 3062 283156 3068
rect 281736 598 281948 626
rect 281736 490 281764 598
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281552 462 281764 490
rect 281920 480 281948 598
rect 283116 480 283144 3062
rect 284312 480 284340 66807
rect 285048 62801 285076 102206
rect 285140 71097 285168 106422
rect 285232 102338 285260 114514
rect 285220 102332 285272 102338
rect 285220 102274 285272 102280
rect 285600 101017 285628 116010
rect 286322 108760 286378 108769
rect 286322 108695 286378 108704
rect 285586 101008 285642 101017
rect 285586 100943 285642 100952
rect 285126 71088 285182 71097
rect 285126 71023 285182 71032
rect 285034 62792 285090 62801
rect 285034 62727 285090 62736
rect 286336 54534 286364 108695
rect 286428 80753 286456 123247
rect 286520 120086 286548 160239
rect 287164 157962 287192 161871
rect 287518 161120 287574 161129
rect 287518 161055 287574 161064
rect 287532 160138 287560 161055
rect 287520 160132 287572 160138
rect 287520 160074 287572 160080
rect 287426 158944 287482 158953
rect 287426 158879 287482 158888
rect 287440 158778 287468 158879
rect 287428 158772 287480 158778
rect 287428 158714 287480 158720
rect 287152 157956 287204 157962
rect 287152 157898 287204 157904
rect 287716 157457 287744 238167
rect 287978 175672 288034 175681
rect 287978 175607 288034 175616
rect 287794 175264 287850 175273
rect 287794 175199 287850 175208
rect 287808 174078 287836 175199
rect 287886 174856 287942 174865
rect 287886 174791 287942 174800
rect 287796 174072 287848 174078
rect 287796 174014 287848 174020
rect 287796 173392 287848 173398
rect 287796 173334 287848 173340
rect 287808 164937 287836 173334
rect 287900 166326 287928 174791
rect 287992 173398 288020 175607
rect 288346 174040 288402 174049
rect 288346 173975 288402 173984
rect 288360 173942 288388 173975
rect 288348 173936 288400 173942
rect 288348 173878 288400 173884
rect 287980 173392 288032 173398
rect 287980 173334 288032 173340
rect 288346 172680 288402 172689
rect 288346 172615 288402 172624
rect 288360 172582 288388 172615
rect 288348 172576 288400 172582
rect 288348 172518 288400 172524
rect 288254 171864 288310 171873
rect 288254 171799 288310 171808
rect 288268 171154 288296 171799
rect 288346 171456 288402 171465
rect 288346 171391 288402 171400
rect 288360 171222 288388 171391
rect 288348 171216 288400 171222
rect 288348 171158 288400 171164
rect 288256 171148 288308 171154
rect 288256 171090 288308 171096
rect 288346 171048 288402 171057
rect 288346 170983 288402 170992
rect 288360 169794 288388 170983
rect 288348 169788 288400 169794
rect 288348 169730 288400 169736
rect 288162 169688 288218 169697
rect 288162 169623 288218 169632
rect 288176 168434 288204 169623
rect 288254 169280 288310 169289
rect 288254 169215 288310 169224
rect 288164 168428 288216 168434
rect 288164 168370 288216 168376
rect 287978 167920 288034 167929
rect 287978 167855 288034 167864
rect 287992 167142 288020 167855
rect 287980 167136 288032 167142
rect 287980 167078 288032 167084
rect 288268 166433 288296 169215
rect 288346 167104 288402 167113
rect 288346 167039 288348 167048
rect 288400 167039 288402 167048
rect 288348 167010 288400 167016
rect 288346 166696 288402 166705
rect 288346 166631 288402 166640
rect 288254 166424 288310 166433
rect 288254 166359 288310 166368
rect 287888 166320 287940 166326
rect 287888 166262 287940 166268
rect 288254 166288 288310 166297
rect 288254 166223 288310 166232
rect 288070 165880 288126 165889
rect 288070 165815 288126 165824
rect 287794 164928 287850 164937
rect 287794 164863 287850 164872
rect 287886 163704 287942 163713
rect 287886 163639 287942 163648
rect 287702 157448 287758 157457
rect 287702 157383 287758 157392
rect 287704 155236 287756 155242
rect 287704 155178 287756 155184
rect 286598 154864 286654 154873
rect 286598 154799 286654 154808
rect 286508 120080 286560 120086
rect 286508 120022 286560 120028
rect 286612 114481 286640 154799
rect 287242 148608 287298 148617
rect 287242 148543 287298 148552
rect 287256 146946 287284 148543
rect 287716 147121 287744 155178
rect 287794 154592 287850 154601
rect 287794 154527 287850 154536
rect 287702 147112 287758 147121
rect 287702 147047 287758 147056
rect 287426 146976 287482 146985
rect 287244 146940 287296 146946
rect 287426 146911 287482 146920
rect 287244 146882 287296 146888
rect 287440 145761 287468 146911
rect 287426 145752 287482 145761
rect 287426 145687 287482 145696
rect 287426 145208 287482 145217
rect 287426 145143 287482 145152
rect 287440 144974 287468 145143
rect 287428 144968 287480 144974
rect 287428 144910 287480 144916
rect 287702 144392 287758 144401
rect 287702 144327 287758 144336
rect 287426 141264 287482 141273
rect 287426 141199 287482 141208
rect 287150 133648 287206 133657
rect 287150 133583 287206 133592
rect 287164 128353 287192 133583
rect 287440 133278 287468 141199
rect 287428 133272 287480 133278
rect 287428 133214 287480 133220
rect 287716 129062 287744 144327
rect 287808 144226 287836 154527
rect 287900 153882 287928 163639
rect 288084 162081 288112 165815
rect 288268 164898 288296 166223
rect 288360 165646 288388 166631
rect 288348 165640 288400 165646
rect 288348 165582 288400 165588
rect 288256 164892 288308 164898
rect 288256 164834 288308 164840
rect 288162 164112 288218 164121
rect 288162 164047 288218 164056
rect 288176 162926 288204 164047
rect 288254 163296 288310 163305
rect 288254 163231 288310 163240
rect 288164 162920 288216 162926
rect 288164 162862 288216 162868
rect 288070 162072 288126 162081
rect 288070 162007 288126 162016
rect 288268 161566 288296 163231
rect 288346 162344 288402 162353
rect 288346 162279 288402 162288
rect 288256 161560 288308 161566
rect 288256 161502 288308 161508
rect 288360 161498 288388 162279
rect 288348 161492 288400 161498
rect 288348 161434 288400 161440
rect 288346 159760 288402 159769
rect 288346 159695 288402 159704
rect 288360 158846 288388 159695
rect 288348 158840 288400 158846
rect 288348 158782 288400 158788
rect 288254 158536 288310 158545
rect 288254 158471 288310 158480
rect 288162 157176 288218 157185
rect 288162 157111 288218 157120
rect 288070 156768 288126 156777
rect 288070 156703 288126 156712
rect 287978 155952 288034 155961
rect 287978 155887 288034 155896
rect 287992 155174 288020 155887
rect 288084 155281 288112 156703
rect 288176 155990 288204 157111
rect 288164 155984 288216 155990
rect 288164 155926 288216 155932
rect 288070 155272 288126 155281
rect 288070 155207 288126 155216
rect 287980 155168 288032 155174
rect 287980 155110 288032 155116
rect 288268 154986 288296 158471
rect 288346 158128 288402 158137
rect 288346 158063 288402 158072
rect 288360 156058 288388 158063
rect 288452 156641 288480 313346
rect 291844 293276 291896 293282
rect 291844 293218 291896 293224
rect 290462 284472 290518 284481
rect 290462 284407 290518 284416
rect 288532 260908 288584 260914
rect 288532 260850 288584 260856
rect 288438 156632 288494 156641
rect 288438 156567 288494 156576
rect 288348 156052 288400 156058
rect 288348 155994 288400 156000
rect 288544 155242 288572 260850
rect 288624 211200 288676 211206
rect 288624 211142 288676 211148
rect 288532 155236 288584 155242
rect 288532 155178 288584 155184
rect 288346 155136 288402 155145
rect 288346 155071 288402 155080
rect 287992 154958 288296 154986
rect 287888 153876 287940 153882
rect 287888 153818 287940 153824
rect 287992 151814 288020 154958
rect 288360 154630 288388 155071
rect 288348 154624 288400 154630
rect 288348 154566 288400 154572
rect 288254 152552 288310 152561
rect 288254 152487 288310 152496
rect 288268 151842 288296 152487
rect 288346 152008 288402 152017
rect 288346 151943 288402 151952
rect 288360 151910 288388 151943
rect 288348 151904 288400 151910
rect 288348 151846 288400 151852
rect 287900 151786 288020 151814
rect 288256 151836 288308 151842
rect 287796 144220 287848 144226
rect 287796 144162 287848 144168
rect 287900 142866 287928 151786
rect 288256 151778 288308 151784
rect 288346 151600 288402 151609
rect 288346 151535 288402 151544
rect 287978 151192 288034 151201
rect 287978 151127 288034 151136
rect 287992 150482 288020 151127
rect 288254 150784 288310 150793
rect 288254 150719 288310 150728
rect 287980 150476 288032 150482
rect 287980 150418 288032 150424
rect 288268 149841 288296 150719
rect 288360 150550 288388 151535
rect 288348 150544 288400 150550
rect 288348 150486 288400 150492
rect 288346 150376 288402 150385
rect 288346 150311 288402 150320
rect 288254 149832 288310 149841
rect 288254 149767 288310 149776
rect 288360 149122 288388 150311
rect 288348 149116 288400 149122
rect 288348 149058 288400 149064
rect 288346 149016 288402 149025
rect 288346 148951 288402 148960
rect 288360 147694 288388 148951
rect 288530 148744 288586 148753
rect 288530 148679 288586 148688
rect 288544 147937 288572 148679
rect 288530 147928 288586 147937
rect 288530 147863 288586 147872
rect 288348 147688 288400 147694
rect 288348 147630 288400 147636
rect 288346 147384 288402 147393
rect 288346 147319 288402 147328
rect 288360 146334 288388 147319
rect 288348 146328 288400 146334
rect 288348 146270 288400 146276
rect 288070 146024 288126 146033
rect 288070 145959 288126 145968
rect 287978 143032 288034 143041
rect 287978 142967 288034 142976
rect 287888 142860 287940 142866
rect 287888 142802 287940 142808
rect 287886 142624 287942 142633
rect 287886 142559 287942 142568
rect 287794 139632 287850 139641
rect 287794 139567 287850 139576
rect 287704 129056 287756 129062
rect 287704 128998 287756 129004
rect 287150 128344 287206 128353
rect 287150 128279 287206 128288
rect 287150 124536 287206 124545
rect 287150 124471 287206 124480
rect 286690 121680 286746 121689
rect 286690 121615 286746 121624
rect 286598 114472 286654 114481
rect 286598 114407 286654 114416
rect 286506 112160 286562 112169
rect 286506 112095 286562 112104
rect 286520 90370 286548 112095
rect 286704 111081 286732 121615
rect 287164 120766 287192 124471
rect 287702 123720 287758 123729
rect 287702 123655 287758 123664
rect 287152 120760 287204 120766
rect 287152 120702 287204 120708
rect 287610 119368 287666 119377
rect 287610 119303 287666 119312
rect 286966 118960 287022 118969
rect 286966 118895 287022 118904
rect 286782 113248 286838 113257
rect 286782 113183 286838 113192
rect 286690 111072 286746 111081
rect 286690 111007 286746 111016
rect 286796 98122 286824 113183
rect 286980 112033 287008 118895
rect 287624 118726 287652 119303
rect 287612 118720 287664 118726
rect 287612 118662 287664 118668
rect 287426 116376 287482 116385
rect 287426 116311 287482 116320
rect 287440 116074 287468 116311
rect 287428 116068 287480 116074
rect 287428 116010 287480 116016
rect 287610 113792 287666 113801
rect 287610 113727 287666 113736
rect 287624 113218 287652 113727
rect 287612 113212 287664 113218
rect 287612 113154 287664 113160
rect 286966 112024 287022 112033
rect 286966 111959 287022 111968
rect 287610 101824 287666 101833
rect 287610 101759 287666 101768
rect 287624 100842 287652 101759
rect 287612 100836 287664 100842
rect 287612 100778 287664 100784
rect 286784 98116 286836 98122
rect 286784 98058 286836 98064
rect 286598 97608 286654 97617
rect 286598 97543 286654 97552
rect 286508 90364 286560 90370
rect 286508 90306 286560 90312
rect 286414 80744 286470 80753
rect 286414 80679 286470 80688
rect 286612 77897 286640 97543
rect 287716 82249 287744 123655
rect 287808 109041 287836 139567
rect 287900 123486 287928 142559
rect 287992 142186 288020 142967
rect 287980 142180 288032 142186
rect 287980 142122 288032 142128
rect 288084 139874 288112 145959
rect 288254 145616 288310 145625
rect 288254 145551 288310 145560
rect 288162 144800 288218 144809
rect 288162 144735 288218 144744
rect 288176 143614 288204 144735
rect 288164 143608 288216 143614
rect 288164 143550 288216 143556
rect 288268 141506 288296 145551
rect 288256 141500 288308 141506
rect 288256 141442 288308 141448
rect 288636 140049 288664 211142
rect 290476 180130 290504 284407
rect 291856 189689 291884 293218
rect 293224 258732 293276 258738
rect 293224 258674 293276 258680
rect 291934 235240 291990 235249
rect 291934 235175 291990 235184
rect 291842 189680 291898 189689
rect 291842 189615 291898 189624
rect 290464 180124 290516 180130
rect 290464 180066 290516 180072
rect 291948 177313 291976 235175
rect 292028 202156 292080 202162
rect 292028 202098 292080 202104
rect 292040 178770 292068 202098
rect 293236 180198 293264 258674
rect 293224 180192 293276 180198
rect 293224 180134 293276 180140
rect 292028 178764 292080 178770
rect 292028 178706 292080 178712
rect 294616 177449 294644 314735
rect 294696 210452 294748 210458
rect 294696 210394 294748 210400
rect 294708 188358 294736 210394
rect 294696 188352 294748 188358
rect 294696 188294 294748 188300
rect 295996 180033 296024 320146
rect 305000 317484 305052 317490
rect 305000 317426 305052 317432
rect 304264 311908 304316 311914
rect 304264 311850 304316 311856
rect 301226 299704 301282 299713
rect 301226 299639 301282 299648
rect 297364 294636 297416 294642
rect 297364 294578 297416 294584
rect 296074 214704 296130 214713
rect 296074 214639 296130 214648
rect 296088 181558 296116 214639
rect 296076 181552 296128 181558
rect 297376 181529 297404 294578
rect 300124 285728 300176 285734
rect 300124 285670 300176 285676
rect 298744 280220 298796 280226
rect 298744 280162 298796 280168
rect 297456 198076 297508 198082
rect 297456 198018 297508 198024
rect 296076 181494 296128 181500
rect 297362 181520 297418 181529
rect 297362 181455 297418 181464
rect 295982 180024 296038 180033
rect 295982 179959 296038 179968
rect 297468 178129 297496 198018
rect 297454 178120 297510 178129
rect 297454 178055 297510 178064
rect 294602 177440 294658 177449
rect 294602 177375 294658 177384
rect 291934 177304 291990 177313
rect 291934 177239 291990 177248
rect 298756 176934 298784 280162
rect 298836 220108 298888 220114
rect 298836 220050 298888 220056
rect 298848 187134 298876 220050
rect 298836 187128 298888 187134
rect 298836 187070 298888 187076
rect 298744 176928 298796 176934
rect 298744 176870 298796 176876
rect 300136 176254 300164 285670
rect 300216 196716 300268 196722
rect 300216 196658 300268 196664
rect 300228 176594 300256 196658
rect 301240 190454 301268 299639
rect 302882 291272 302938 291281
rect 302882 291207 302938 291216
rect 302240 245676 302292 245682
rect 302240 245618 302292 245624
rect 301504 238060 301556 238066
rect 301504 238002 301556 238008
rect 301240 190426 301360 190454
rect 301044 181484 301096 181490
rect 301044 181426 301096 181432
rect 300858 176760 300914 176769
rect 300858 176695 300914 176704
rect 300216 176588 300268 176594
rect 300216 176530 300268 176536
rect 300124 176248 300176 176254
rect 300124 176190 300176 176196
rect 300872 176089 300900 176695
rect 300858 176080 300914 176089
rect 300858 176015 300914 176024
rect 298190 175944 298246 175953
rect 298190 175879 298246 175888
rect 298204 175846 298232 175879
rect 298192 175840 298244 175846
rect 298192 175782 298244 175788
rect 289174 167512 289230 167521
rect 289174 167447 289230 167456
rect 288714 164656 288770 164665
rect 288714 164591 288770 164600
rect 288728 164490 288756 164591
rect 288716 164484 288768 164490
rect 288716 164426 288768 164432
rect 289082 153776 289138 153785
rect 289082 153711 289138 153720
rect 288622 140040 288678 140049
rect 288622 139975 288678 139984
rect 288072 139868 288124 139874
rect 288072 139810 288124 139816
rect 288254 139224 288310 139233
rect 288254 139159 288310 139168
rect 288268 138106 288296 139159
rect 288346 138272 288402 138281
rect 288346 138207 288402 138216
rect 288256 138100 288308 138106
rect 288256 138042 288308 138048
rect 288360 138038 288388 138207
rect 288348 138032 288400 138038
rect 288348 137974 288400 137980
rect 288346 137456 288402 137465
rect 288346 137391 288402 137400
rect 288360 136678 288388 137391
rect 288348 136672 288400 136678
rect 288348 136614 288400 136620
rect 288346 133104 288402 133113
rect 288346 133039 288402 133048
rect 288360 132530 288388 133039
rect 288348 132524 288400 132530
rect 288348 132466 288400 132472
rect 288346 132288 288402 132297
rect 288346 132223 288402 132232
rect 288360 131170 288388 132223
rect 288348 131164 288400 131170
rect 288348 131106 288400 131112
rect 288346 130520 288402 130529
rect 288346 130455 288402 130464
rect 288360 129810 288388 130455
rect 288348 129804 288400 129810
rect 288348 129746 288400 129752
rect 288070 129704 288126 129713
rect 288070 129639 288126 129648
rect 287978 129296 288034 129305
rect 287978 129231 288034 129240
rect 287992 128382 288020 129231
rect 287980 128376 288032 128382
rect 287980 128318 288032 128324
rect 287978 127936 288034 127945
rect 287978 127871 288034 127880
rect 287992 127022 288020 127871
rect 287980 127016 288032 127022
rect 287980 126958 288032 126964
rect 288084 124817 288112 129639
rect 288162 127528 288218 127537
rect 288162 127463 288218 127472
rect 288070 124808 288126 124817
rect 288070 124743 288126 124752
rect 287978 124128 288034 124137
rect 287978 124063 288034 124072
rect 287888 123480 287940 123486
rect 287888 123422 287940 123428
rect 287992 122874 288020 124063
rect 287980 122868 288032 122874
rect 287980 122810 288032 122816
rect 288176 122834 288204 127463
rect 288254 126304 288310 126313
rect 288254 126239 288310 126248
rect 288268 125730 288296 126239
rect 288346 125896 288402 125905
rect 288346 125831 288402 125840
rect 288256 125724 288308 125730
rect 288256 125666 288308 125672
rect 288360 125662 288388 125831
rect 288348 125656 288400 125662
rect 288348 125598 288400 125604
rect 288346 125352 288402 125361
rect 288346 125287 288402 125296
rect 288360 124234 288388 125287
rect 288348 124228 288400 124234
rect 288348 124170 288400 124176
rect 288530 123856 288586 123865
rect 288530 123791 288586 123800
rect 288544 123049 288572 123791
rect 288530 123040 288586 123049
rect 288530 122975 288586 122984
rect 288176 122806 288388 122834
rect 288254 121544 288310 121553
rect 288254 121479 288256 121488
rect 288308 121479 288310 121488
rect 288256 121450 288308 121456
rect 288254 121136 288310 121145
rect 288254 121071 288310 121080
rect 288268 120154 288296 121071
rect 288256 120148 288308 120154
rect 288256 120090 288308 120096
rect 288254 117736 288310 117745
rect 288254 117671 288310 117680
rect 288268 117366 288296 117671
rect 288256 117360 288308 117366
rect 288256 117302 288308 117308
rect 288162 117192 288218 117201
rect 288162 117127 288218 117136
rect 288176 116006 288204 117127
rect 288164 116000 288216 116006
rect 288164 115942 288216 115948
rect 288070 115152 288126 115161
rect 288070 115087 288126 115096
rect 287978 114200 288034 114209
rect 287978 114135 288034 114144
rect 287992 113286 288020 114135
rect 287980 113280 288032 113286
rect 287980 113222 288032 113228
rect 287886 113112 287942 113121
rect 287886 113047 287942 113056
rect 287794 109032 287850 109041
rect 287794 108967 287850 108976
rect 287900 98190 287928 113047
rect 287978 111616 288034 111625
rect 287978 111551 288034 111560
rect 287992 110566 288020 111551
rect 287980 110560 288032 110566
rect 287980 110502 288032 110508
rect 287978 107400 288034 107409
rect 287978 107335 288034 107344
rect 287992 106486 288020 107335
rect 287980 106480 288032 106486
rect 287980 106422 288032 106428
rect 287978 105632 288034 105641
rect 287978 105567 288034 105576
rect 287992 104990 288020 105567
rect 287980 104984 288032 104990
rect 287980 104926 288032 104932
rect 288084 103514 288112 115087
rect 288254 114608 288310 114617
rect 288254 114543 288256 114552
rect 288308 114543 288310 114552
rect 288256 114514 288308 114520
rect 288360 112033 288388 122806
rect 289096 113150 289124 153711
rect 289188 135930 289216 167447
rect 301056 151814 301084 181426
rect 301136 176248 301188 176254
rect 301136 176190 301188 176196
rect 301148 161474 301176 176190
rect 301332 170649 301360 190426
rect 301412 178764 301464 178770
rect 301412 178706 301464 178712
rect 301424 175273 301452 178706
rect 301516 178702 301544 238002
rect 301596 235272 301648 235278
rect 301596 235214 301648 235220
rect 301608 184278 301636 235214
rect 301686 189816 301742 189825
rect 301686 189751 301742 189760
rect 301596 184272 301648 184278
rect 301596 184214 301648 184220
rect 301504 178696 301556 178702
rect 301504 178638 301556 178644
rect 301700 176633 301728 189751
rect 301686 176624 301742 176633
rect 301686 176559 301742 176568
rect 301410 175264 301466 175273
rect 301410 175199 301466 175208
rect 301412 175160 301464 175166
rect 301412 175102 301464 175108
rect 301424 174457 301452 175102
rect 301410 174448 301466 174457
rect 301410 174383 301466 174392
rect 301318 170640 301374 170649
rect 301318 170575 301374 170584
rect 301148 161446 301360 161474
rect 301332 160857 301360 161446
rect 301318 160848 301374 160857
rect 301318 160783 301374 160792
rect 301056 151786 301360 151814
rect 301332 150657 301360 151786
rect 301318 150648 301374 150657
rect 301318 150583 301374 150592
rect 289358 138680 289414 138689
rect 289358 138615 289414 138624
rect 289266 136232 289322 136241
rect 289266 136167 289322 136176
rect 289176 135924 289228 135930
rect 289176 135866 289228 135872
rect 289174 131064 289230 131073
rect 289174 130999 289230 131008
rect 289084 113144 289136 113150
rect 289084 113086 289136 113092
rect 288346 112024 288402 112033
rect 288346 111959 288402 111968
rect 288254 111208 288310 111217
rect 288254 111143 288310 111152
rect 288268 110498 288296 111143
rect 288256 110492 288308 110498
rect 288256 110434 288308 110440
rect 288254 110392 288310 110401
rect 288254 110327 288310 110336
rect 288268 109138 288296 110327
rect 288346 109576 288402 109585
rect 288346 109511 288402 109520
rect 288256 109132 288308 109138
rect 288256 109074 288308 109080
rect 288360 109070 288388 109511
rect 288348 109064 288400 109070
rect 288348 109006 288400 109012
rect 288346 108624 288402 108633
rect 288346 108559 288402 108568
rect 288360 107710 288388 108559
rect 289082 108216 289138 108225
rect 289082 108151 289138 108160
rect 288348 107704 288400 107710
rect 288348 107646 288400 107652
rect 288346 106992 288402 107001
rect 288346 106927 288402 106936
rect 288360 106418 288388 106927
rect 288348 106412 288400 106418
rect 288348 106354 288400 106360
rect 288346 106040 288402 106049
rect 288346 105975 288402 105984
rect 288360 104922 288388 105975
rect 288348 104916 288400 104922
rect 288348 104858 288400 104864
rect 288530 104000 288586 104009
rect 288530 103935 288586 103944
rect 288544 103601 288572 103935
rect 288530 103592 288586 103601
rect 288530 103527 288586 103536
rect 287992 103486 288112 103514
rect 287992 102513 288020 103486
rect 288346 103456 288402 103465
rect 288346 103391 288402 103400
rect 288254 102640 288310 102649
rect 288254 102575 288310 102584
rect 287978 102504 288034 102513
rect 287978 102439 288034 102448
rect 288268 102202 288296 102575
rect 288360 102270 288388 103391
rect 288348 102264 288400 102270
rect 288348 102206 288400 102212
rect 288256 102196 288308 102202
rect 288256 102138 288308 102144
rect 288346 101280 288402 101289
rect 288346 101215 288402 101224
rect 288360 100774 288388 101215
rect 288348 100768 288400 100774
rect 288348 100710 288400 100716
rect 288254 100464 288310 100473
rect 288254 100399 288310 100408
rect 288268 99482 288296 100399
rect 288346 99648 288402 99657
rect 288346 99583 288402 99592
rect 288256 99476 288308 99482
rect 288256 99418 288308 99424
rect 288360 99414 288388 99583
rect 288348 99408 288400 99414
rect 288348 99350 288400 99356
rect 288530 98832 288586 98841
rect 288530 98767 288586 98776
rect 288544 98297 288572 98767
rect 288530 98288 288586 98297
rect 288530 98223 288586 98232
rect 287888 98184 287940 98190
rect 287888 98126 287940 98132
rect 287794 98016 287850 98025
rect 287794 97951 287850 97960
rect 287702 82240 287758 82249
rect 287702 82175 287758 82184
rect 287808 78033 287836 97951
rect 287886 97472 287942 97481
rect 287886 97407 287942 97416
rect 287900 86193 287928 97407
rect 288348 97300 288400 97306
rect 288348 97242 288400 97248
rect 288360 97073 288388 97242
rect 288346 97064 288402 97073
rect 288346 96999 288402 97008
rect 287886 86184 287942 86193
rect 287886 86119 287942 86128
rect 287794 78024 287850 78033
rect 287794 77959 287850 77968
rect 286598 77888 286654 77897
rect 286598 77823 286654 77832
rect 286324 54528 286376 54534
rect 286324 54470 286376 54476
rect 289096 50386 289124 108151
rect 289188 79393 289216 130999
rect 289280 130422 289308 136167
rect 289268 130416 289320 130422
rect 289372 130393 289400 138615
rect 289450 136640 289506 136649
rect 289450 136575 289506 136584
rect 289268 130358 289320 130364
rect 289358 130384 289414 130393
rect 289358 130319 289414 130328
rect 289464 122233 289492 136575
rect 302252 125225 302280 245618
rect 302896 188465 302924 291207
rect 303620 261520 303672 261526
rect 303620 261462 303672 261468
rect 302882 188456 302938 188465
rect 302882 188391 302938 188400
rect 302332 188352 302384 188358
rect 302332 188294 302384 188300
rect 302344 185842 302372 188294
rect 302424 187128 302476 187134
rect 302424 187070 302476 187076
rect 302332 185836 302384 185842
rect 302332 185778 302384 185784
rect 302330 185736 302386 185745
rect 302330 185671 302386 185680
rect 302344 161809 302372 185671
rect 302436 182170 302464 187070
rect 302424 182164 302476 182170
rect 302424 182106 302476 182112
rect 302514 178120 302570 178129
rect 302514 178055 302570 178064
rect 302424 177336 302476 177342
rect 302424 177278 302476 177284
rect 302330 161800 302386 161809
rect 302330 161735 302386 161744
rect 302436 159497 302464 177278
rect 302528 168745 302556 178055
rect 303632 172553 303660 261462
rect 304276 202337 304304 311850
rect 304354 213344 304410 213353
rect 304354 213279 304410 213288
rect 304262 202328 304318 202337
rect 304262 202263 304318 202272
rect 304264 200796 304316 200802
rect 304264 200738 304316 200744
rect 304276 183025 304304 200738
rect 304368 183530 304396 213279
rect 304448 185836 304500 185842
rect 304448 185778 304500 185784
rect 304356 183524 304408 183530
rect 304356 183466 304408 183472
rect 304262 183016 304318 183025
rect 304262 182951 304318 182960
rect 303804 182912 303856 182918
rect 303804 182854 303856 182860
rect 303712 182164 303764 182170
rect 303712 182106 303764 182112
rect 303618 172544 303674 172553
rect 303618 172479 303674 172488
rect 302514 168736 302570 168745
rect 302514 168671 302570 168680
rect 302422 159488 302478 159497
rect 302422 159423 302478 159432
rect 303620 158704 303672 158710
rect 303620 158646 303672 158652
rect 303632 158001 303660 158646
rect 303618 157992 303674 158001
rect 303618 157927 303674 157936
rect 303620 155916 303672 155922
rect 303620 155858 303672 155864
rect 303632 155009 303660 155858
rect 303618 155000 303674 155009
rect 303618 154935 303674 154944
rect 303620 154488 303672 154494
rect 303620 154430 303672 154436
rect 303632 154193 303660 154430
rect 303618 154184 303674 154193
rect 303618 154119 303674 154128
rect 303724 151201 303752 182106
rect 303816 160018 303844 182854
rect 304460 180033 304488 185778
rect 304446 180024 304502 180033
rect 304446 179959 304502 179968
rect 303896 172508 303948 172514
rect 303896 172450 303948 172456
rect 303908 171737 303936 172450
rect 303894 171728 303950 171737
rect 303894 171663 303950 171672
rect 304906 170912 304962 170921
rect 305012 170898 305040 317426
rect 315946 310584 316002 310593
rect 315946 310519 316002 310528
rect 315960 306649 315988 310519
rect 315946 306640 316002 306649
rect 315946 306575 316002 306584
rect 315946 306368 316002 306377
rect 315946 306303 316002 306312
rect 315960 296857 315988 306303
rect 315946 296848 316002 296857
rect 315946 296783 316002 296792
rect 315946 296712 316002 296721
rect 315946 296647 316002 296656
rect 313278 292904 313334 292913
rect 313278 292839 313334 292848
rect 309138 289912 309194 289921
rect 309138 289847 309194 289856
rect 307022 284064 307078 284073
rect 307022 283999 307078 284008
rect 306656 260160 306708 260166
rect 306656 260102 306708 260108
rect 305092 254584 305144 254590
rect 305092 254526 305144 254532
rect 304962 170870 305040 170898
rect 304906 170847 304962 170856
rect 303896 169720 303948 169726
rect 303896 169662 303948 169668
rect 303908 169425 303936 169662
rect 303894 169416 303950 169425
rect 303894 169351 303950 169360
rect 303896 168360 303948 168366
rect 303896 168302 303948 168308
rect 303908 167113 303936 168302
rect 303894 167104 303950 167113
rect 303894 167039 303950 167048
rect 303896 167000 303948 167006
rect 303896 166942 303948 166948
rect 303908 166433 303936 166942
rect 303894 166424 303950 166433
rect 303894 166359 303950 166368
rect 304264 166320 304316 166326
rect 304264 166262 304316 166268
rect 303896 165572 303948 165578
rect 303896 165514 303948 165520
rect 303908 164937 303936 165514
rect 303894 164928 303950 164937
rect 303894 164863 303950 164872
rect 303896 164212 303948 164218
rect 303896 164154 303948 164160
rect 303908 164121 303936 164154
rect 303894 164112 303950 164121
rect 303894 164047 303950 164056
rect 303896 163328 303948 163334
rect 303894 163296 303896 163305
rect 303948 163296 303950 163305
rect 303894 163231 303950 163240
rect 303896 162852 303948 162858
rect 303896 162794 303948 162800
rect 303908 162625 303936 162794
rect 303894 162616 303950 162625
rect 303894 162551 303950 162560
rect 303896 161424 303948 161430
rect 303896 161366 303948 161372
rect 303908 161129 303936 161366
rect 303894 161120 303950 161129
rect 303894 161055 303950 161064
rect 303816 159990 303936 160018
rect 303804 159928 303856 159934
rect 303804 159870 303856 159876
rect 303816 158817 303844 159870
rect 303802 158808 303858 158817
rect 303802 158743 303858 158752
rect 303804 157344 303856 157350
rect 303802 157312 303804 157321
rect 303856 157312 303858 157321
rect 303802 157247 303858 157256
rect 303908 156505 303936 159990
rect 303894 156496 303950 156505
rect 303894 156431 303950 156440
rect 303804 155848 303856 155854
rect 303804 155790 303856 155796
rect 303816 155689 303844 155790
rect 303802 155680 303858 155689
rect 303802 155615 303858 155624
rect 303804 154556 303856 154562
rect 303804 154498 303856 154504
rect 303816 153513 303844 154498
rect 303802 153504 303858 153513
rect 303802 153439 303858 153448
rect 303804 153196 303856 153202
rect 303804 153138 303856 153144
rect 303816 152697 303844 153138
rect 303896 153128 303948 153134
rect 303896 153070 303948 153076
rect 303802 152688 303858 152697
rect 303802 152623 303858 152632
rect 303908 151881 303936 153070
rect 303894 151872 303950 151881
rect 303894 151807 303950 151816
rect 303710 151192 303766 151201
rect 303710 151127 303766 151136
rect 303804 150408 303856 150414
rect 303804 150350 303856 150356
rect 303816 149705 303844 150350
rect 303802 149696 303858 149705
rect 303802 149631 303858 149640
rect 303804 149048 303856 149054
rect 303804 148990 303856 148996
rect 303816 148889 303844 148990
rect 303802 148880 303858 148889
rect 303802 148815 303858 148824
rect 303712 147620 303764 147626
rect 303712 147562 303764 147568
rect 303724 147393 303752 147562
rect 303710 147384 303766 147393
rect 303710 147319 303766 147328
rect 303804 146260 303856 146266
rect 303804 146202 303856 146208
rect 303816 145897 303844 146202
rect 303802 145888 303858 145897
rect 303712 145852 303764 145858
rect 303802 145823 303858 145832
rect 303712 145794 303764 145800
rect 303724 145081 303752 145794
rect 303710 145072 303766 145081
rect 303710 145007 303766 145016
rect 303804 144900 303856 144906
rect 303804 144842 303856 144848
rect 303816 144265 303844 144842
rect 303802 144256 303858 144265
rect 303802 144191 303858 144200
rect 303988 144220 304040 144226
rect 303988 144162 304040 144168
rect 303804 142112 303856 142118
rect 304000 142089 304028 144162
rect 303804 142054 303856 142060
rect 303986 142080 304042 142089
rect 303816 141273 303844 142054
rect 303986 142015 304042 142024
rect 303802 141264 303858 141273
rect 303802 141199 303858 141208
rect 303620 139868 303672 139874
rect 303620 139810 303672 139816
rect 303632 139777 303660 139810
rect 303618 139768 303674 139777
rect 303618 139703 303674 139712
rect 303804 139392 303856 139398
rect 303804 139334 303856 139340
rect 303816 138281 303844 139334
rect 304276 138961 304304 166262
rect 305104 151814 305132 254526
rect 306472 198008 306524 198014
rect 306472 197950 306524 197956
rect 305184 189780 305236 189786
rect 305184 189722 305236 189728
rect 305012 151786 305132 151814
rect 304906 148064 304962 148073
rect 305012 148050 305040 151786
rect 304962 148022 305040 148050
rect 304906 147999 304962 148008
rect 304262 138952 304318 138961
rect 304262 138887 304318 138896
rect 303802 138272 303858 138281
rect 303802 138207 303858 138216
rect 303804 137964 303856 137970
rect 303804 137906 303856 137912
rect 303816 137465 303844 137906
rect 303802 137456 303858 137465
rect 303802 137391 303858 137400
rect 303620 136604 303672 136610
rect 303620 136546 303672 136552
rect 303632 135969 303660 136546
rect 303618 135960 303674 135969
rect 303618 135895 303674 135904
rect 303712 135244 303764 135250
rect 303712 135186 303764 135192
rect 303724 134473 303752 135186
rect 304724 134564 304776 134570
rect 304724 134506 304776 134512
rect 303710 134464 303766 134473
rect 303710 134399 303766 134408
rect 303896 133884 303948 133890
rect 303896 133826 303948 133832
rect 303804 133816 303856 133822
rect 303804 133758 303856 133764
rect 303816 133657 303844 133758
rect 303802 133648 303858 133657
rect 303802 133583 303858 133592
rect 303908 132841 303936 133826
rect 303894 132832 303950 132841
rect 303894 132767 303950 132776
rect 303804 132456 303856 132462
rect 303804 132398 303856 132404
rect 303816 132161 303844 132398
rect 303896 132388 303948 132394
rect 303896 132330 303948 132336
rect 303802 132152 303858 132161
rect 303802 132087 303858 132096
rect 303908 131345 303936 132330
rect 303894 131336 303950 131345
rect 303894 131271 303950 131280
rect 303804 131096 303856 131102
rect 303804 131038 303856 131044
rect 303816 130665 303844 131038
rect 303802 130656 303858 130665
rect 303802 130591 303858 130600
rect 304264 130416 304316 130422
rect 304264 130358 304316 130364
rect 303804 129736 303856 129742
rect 303804 129678 303856 129684
rect 303816 129033 303844 129678
rect 303802 129024 303858 129033
rect 303802 128959 303858 128968
rect 303802 128344 303858 128353
rect 303802 128279 303804 128288
rect 303856 128279 303858 128288
rect 303804 128250 303856 128256
rect 303620 128240 303672 128246
rect 303620 128182 303672 128188
rect 303632 127537 303660 128182
rect 303618 127528 303674 127537
rect 303618 127463 303674 127472
rect 303712 125588 303764 125594
rect 303712 125530 303764 125536
rect 302238 125216 302294 125225
rect 302238 125151 302294 125160
rect 303724 124545 303752 125530
rect 303710 124536 303766 124545
rect 303710 124471 303766 124480
rect 303712 124160 303764 124166
rect 303712 124102 303764 124108
rect 303724 123049 303752 124102
rect 303804 124092 303856 124098
rect 303804 124034 303856 124040
rect 303816 123729 303844 124034
rect 303802 123720 303858 123729
rect 303802 123655 303858 123664
rect 303710 123040 303766 123049
rect 303710 122975 303766 122984
rect 303620 122800 303672 122806
rect 303620 122742 303672 122748
rect 303632 122233 303660 122742
rect 289450 122224 289506 122233
rect 289450 122159 289506 122168
rect 303618 122224 303674 122233
rect 303618 122159 303674 122168
rect 289266 121952 289322 121961
rect 289266 121887 289322 121896
rect 289174 79384 289230 79393
rect 289174 79319 289230 79328
rect 289280 75177 289308 121887
rect 303804 121440 303856 121446
rect 303802 121408 303804 121417
rect 303856 121408 303858 121417
rect 303802 121343 303858 121352
rect 303804 120080 303856 120086
rect 303804 120022 303856 120028
rect 303816 119241 303844 120022
rect 303802 119232 303858 119241
rect 303802 119167 303858 119176
rect 303896 118652 303948 118658
rect 303896 118594 303948 118600
rect 303804 118448 303856 118454
rect 303802 118416 303804 118425
rect 303856 118416 303858 118425
rect 303802 118351 303858 118360
rect 303908 117609 303936 118594
rect 303894 117600 303950 117609
rect 303894 117535 303950 117544
rect 303804 117292 303856 117298
rect 303804 117234 303856 117240
rect 289726 116784 289782 116793
rect 289726 116719 289782 116728
rect 289740 95130 289768 116719
rect 303816 116113 303844 117234
rect 303802 116104 303858 116113
rect 303802 116039 303858 116048
rect 303804 115932 303856 115938
rect 303804 115874 303856 115880
rect 303620 115456 303672 115462
rect 303618 115424 303620 115433
rect 303672 115424 303674 115433
rect 303618 115359 303674 115368
rect 303816 114617 303844 115874
rect 303802 114608 303858 114617
rect 303802 114543 303858 114552
rect 303804 114504 303856 114510
rect 303804 114446 303856 114452
rect 303816 113801 303844 114446
rect 303802 113792 303858 113801
rect 303802 113727 303858 113736
rect 303804 113144 303856 113150
rect 303802 113112 303804 113121
rect 303856 113112 303858 113121
rect 303802 113047 303858 113056
rect 303712 112804 303764 112810
rect 303712 112746 303764 112752
rect 303724 112305 303752 112746
rect 303710 112296 303766 112305
rect 303710 112231 303766 112240
rect 303712 111784 303764 111790
rect 303712 111726 303764 111732
rect 303724 110809 303752 111726
rect 303804 111716 303856 111722
rect 303804 111658 303856 111664
rect 303816 111625 303844 111658
rect 303802 111616 303858 111625
rect 303802 111551 303858 111560
rect 303710 110800 303766 110809
rect 303710 110735 303766 110744
rect 303804 108996 303856 109002
rect 303804 108938 303856 108944
rect 303816 107817 303844 108938
rect 304276 108497 304304 130358
rect 304736 126041 304764 134506
rect 305196 129849 305224 189722
rect 305276 183524 305328 183530
rect 305276 183466 305328 183472
rect 305288 177410 305316 183466
rect 305276 177404 305328 177410
rect 305276 177346 305328 177352
rect 305276 176928 305328 176934
rect 305276 176870 305328 176876
rect 305288 139874 305316 176870
rect 305276 139868 305328 139874
rect 305276 139810 305328 139816
rect 305182 129840 305238 129849
rect 305182 129775 305238 129784
rect 304722 126032 304778 126041
rect 304722 125967 304778 125976
rect 304354 123448 304410 123457
rect 304354 123383 304410 123392
rect 304262 108488 304318 108497
rect 304262 108423 304318 108432
rect 303802 107808 303858 107817
rect 303802 107743 303858 107752
rect 303804 107636 303856 107642
rect 303804 107578 303856 107584
rect 303816 107001 303844 107578
rect 303802 106992 303858 107001
rect 303802 106927 303858 106936
rect 303710 105496 303766 105505
rect 303710 105431 303766 105440
rect 303724 103514 303752 105431
rect 303804 104848 303856 104854
rect 303804 104790 303856 104796
rect 303816 104009 303844 104790
rect 304368 104689 304396 123383
rect 306484 115462 306512 197950
rect 306564 176588 306616 176594
rect 306564 176530 306616 176536
rect 306576 159934 306604 176530
rect 306564 159928 306616 159934
rect 306564 159870 306616 159876
rect 306472 115456 306524 115462
rect 306472 115398 306524 115404
rect 306668 112810 306696 260102
rect 307036 177342 307064 283999
rect 307760 224324 307812 224330
rect 307760 224266 307812 224272
rect 307024 177336 307076 177342
rect 307024 177278 307076 177284
rect 307772 113150 307800 224266
rect 308404 206304 308456 206310
rect 308404 206246 308456 206252
rect 307942 202192 307998 202201
rect 307942 202127 307998 202136
rect 307850 182880 307906 182889
rect 307850 182815 307906 182824
rect 307864 118454 307892 182815
rect 307956 163334 307984 202127
rect 308036 181552 308088 181558
rect 308036 181494 308088 181500
rect 307944 163328 307996 163334
rect 307944 163270 307996 163276
rect 308048 145858 308076 181494
rect 308416 181490 308444 206246
rect 308404 181484 308456 181490
rect 308404 181426 308456 181432
rect 308036 145852 308088 145858
rect 308036 145794 308088 145800
rect 307852 118448 307904 118454
rect 307852 118390 307904 118396
rect 307760 113144 307812 113150
rect 307760 113086 307812 113092
rect 306656 112804 306708 112810
rect 306656 112746 306708 112752
rect 309152 107642 309180 289847
rect 309230 285968 309286 285977
rect 309230 285903 309286 285912
rect 309244 123457 309272 285903
rect 312176 269816 312228 269822
rect 312176 269758 312228 269764
rect 310520 244928 310572 244934
rect 310520 244870 310572 244876
rect 309416 187060 309468 187066
rect 309416 187002 309468 187008
rect 309322 177304 309378 177313
rect 309322 177239 309378 177248
rect 309336 143585 309364 177239
rect 309428 165578 309456 187002
rect 309416 165572 309468 165578
rect 309416 165514 309468 165520
rect 309322 143576 309378 143585
rect 309322 143511 309378 143520
rect 309230 123448 309286 123457
rect 309230 123383 309286 123392
rect 310532 115938 310560 244870
rect 311992 207664 312044 207670
rect 311992 207606 312044 207612
rect 310612 192500 310664 192506
rect 310612 192442 310664 192448
rect 310624 136610 310652 192442
rect 310796 185700 310848 185706
rect 310796 185642 310848 185648
rect 310704 180192 310756 180198
rect 310704 180134 310756 180140
rect 310716 158710 310744 180134
rect 310808 167006 310836 185642
rect 311900 177404 311952 177410
rect 311900 177346 311952 177352
rect 311912 169726 311940 177346
rect 311900 169720 311952 169726
rect 311900 169662 311952 169668
rect 310796 167000 310848 167006
rect 310796 166942 310848 166948
rect 310704 158704 310756 158710
rect 310704 158646 310756 158652
rect 310612 136604 310664 136610
rect 310612 136546 310664 136552
rect 312004 118658 312032 207606
rect 312084 184204 312136 184210
rect 312084 184146 312136 184152
rect 312096 153134 312124 184146
rect 312084 153128 312136 153134
rect 312084 153070 312136 153076
rect 312188 134570 312216 269758
rect 312176 134564 312228 134570
rect 312176 134506 312228 134512
rect 311992 118652 312044 118658
rect 311992 118594 312044 118600
rect 310520 115932 310572 115938
rect 310520 115874 310572 115880
rect 313292 111722 313320 292839
rect 315960 287201 315988 296647
rect 315946 287192 316002 287201
rect 315946 287127 316002 287136
rect 315946 287056 316002 287065
rect 315946 286991 316002 287000
rect 313924 284368 313976 284374
rect 313924 284310 313976 284316
rect 313372 225072 313424 225078
rect 313372 225014 313424 225020
rect 313384 128246 313412 225014
rect 313464 184272 313516 184278
rect 313464 184214 313516 184220
rect 313476 134609 313504 184214
rect 313556 180124 313608 180130
rect 313556 180066 313608 180072
rect 313568 157350 313596 180066
rect 313936 179926 313964 284310
rect 315960 277545 315988 286991
rect 315946 277536 316002 277545
rect 315946 277471 316002 277480
rect 315946 277400 316002 277409
rect 315946 277335 316002 277344
rect 315960 267889 315988 277335
rect 315946 267880 316002 267889
rect 315946 267815 316002 267824
rect 315946 267744 316002 267753
rect 315946 267679 316002 267688
rect 315960 248441 315988 267679
rect 315946 248432 316002 248441
rect 315946 248367 316002 248376
rect 315946 248296 316002 248305
rect 315946 248231 316002 248240
rect 315960 238785 315988 248231
rect 315946 238776 316002 238785
rect 315946 238711 316002 238720
rect 315946 238640 316002 238649
rect 315946 238575 316002 238584
rect 314660 231872 314712 231878
rect 314660 231814 314712 231820
rect 313924 179920 313976 179926
rect 313924 179862 313976 179868
rect 313556 157344 313608 157350
rect 313556 157286 313608 157292
rect 313462 134600 313518 134609
rect 313462 134535 313518 134544
rect 313372 128240 313424 128246
rect 313372 128182 313424 128188
rect 314672 117298 314700 231814
rect 315960 229129 315988 238575
rect 316038 233880 316094 233889
rect 316038 233815 316094 233824
rect 315946 229120 316002 229129
rect 315946 229055 316002 229064
rect 315946 228984 316002 228993
rect 315946 228919 316002 228928
rect 315960 219473 315988 228919
rect 315946 219464 316002 219473
rect 315946 219399 316002 219408
rect 315946 219328 316002 219337
rect 315946 219263 316002 219272
rect 315960 209817 315988 219263
rect 315946 209808 316002 209817
rect 315946 209743 316002 209752
rect 315946 209672 316002 209681
rect 315946 209607 316002 209616
rect 314752 200864 314804 200870
rect 314752 200806 314804 200812
rect 314660 117292 314712 117298
rect 314660 117234 314712 117240
rect 313280 111716 313332 111722
rect 313280 111658 313332 111664
rect 309140 107636 309192 107642
rect 309140 107578 309192 107584
rect 314764 104854 314792 200806
rect 315960 200161 315988 209607
rect 315946 200152 316002 200161
rect 315946 200087 316002 200096
rect 315946 200016 316002 200025
rect 315946 199951 316002 199960
rect 314844 196648 314896 196654
rect 314844 196590 314896 196596
rect 314856 139398 314884 196590
rect 315960 190505 315988 199951
rect 315946 190496 316002 190505
rect 315946 190431 316002 190440
rect 315946 190360 316002 190369
rect 315946 190295 316002 190304
rect 314934 183016 314990 183025
rect 314934 182951 314990 182960
rect 314844 139392 314896 139398
rect 314844 139334 314896 139340
rect 314948 129742 314976 182951
rect 315960 180849 315988 190295
rect 315946 180840 316002 180849
rect 315946 180775 316002 180784
rect 315946 180704 316002 180713
rect 315946 180639 316002 180648
rect 315960 171193 315988 180639
rect 315946 171184 316002 171193
rect 315946 171119 316002 171128
rect 315946 171048 316002 171057
rect 315946 170983 316002 170992
rect 315960 161537 315988 170983
rect 315946 161528 316002 161537
rect 315946 161463 316002 161472
rect 315946 161392 316002 161401
rect 315946 161327 316002 161336
rect 315960 151881 315988 161327
rect 315946 151872 316002 151881
rect 315946 151807 316002 151816
rect 315946 151736 316002 151745
rect 315946 151671 316002 151680
rect 315960 142225 315988 151671
rect 315946 142216 316002 142225
rect 315946 142151 316002 142160
rect 315946 142080 316002 142089
rect 315946 142015 316002 142024
rect 315960 132569 315988 142015
rect 315946 132560 316002 132569
rect 315946 132495 316002 132504
rect 315946 132424 316002 132433
rect 315946 132359 316002 132368
rect 314936 129736 314988 129742
rect 314936 129678 314988 129684
rect 315960 122913 315988 132359
rect 315946 122904 316002 122913
rect 315946 122839 316002 122848
rect 315946 122768 316002 122777
rect 315946 122703 316002 122712
rect 315960 119377 315988 122703
rect 315946 119368 316002 119377
rect 315946 119303 316002 119312
rect 316052 114510 316080 233815
rect 316224 228404 316276 228410
rect 316224 228346 316276 228352
rect 316132 215960 316184 215966
rect 316132 215902 316184 215908
rect 316144 144226 316172 215902
rect 316236 172514 316264 228346
rect 316316 177336 316368 177342
rect 316316 177278 316368 177284
rect 316224 172508 316276 172514
rect 316224 172450 316276 172456
rect 316328 150414 316356 177278
rect 316316 150408 316368 150414
rect 316316 150350 316368 150356
rect 316132 144220 316184 144226
rect 316132 144162 316184 144168
rect 316040 114504 316092 114510
rect 316040 114446 316092 114452
rect 314752 104848 314804 104854
rect 314752 104790 314804 104796
rect 304354 104680 304410 104689
rect 304354 104615 304410 104624
rect 303802 104000 303858 104009
rect 303802 103935 303858 103944
rect 303724 103486 303844 103514
rect 303618 103184 303674 103193
rect 303618 103119 303674 103128
rect 303632 101538 303660 103119
rect 303712 102128 303764 102134
rect 303712 102070 303764 102076
rect 303724 101697 303752 102070
rect 303710 101688 303766 101697
rect 303710 101623 303766 101632
rect 303632 101510 303752 101538
rect 301318 100600 301374 100609
rect 301148 100558 301318 100586
rect 290924 96008 290976 96014
rect 290924 95950 290976 95956
rect 289728 95124 289780 95130
rect 289728 95066 289780 95072
rect 289818 94888 289874 94897
rect 289818 94823 289874 94832
rect 289832 76809 289860 94823
rect 290936 93770 290964 95950
rect 291106 95704 291162 95713
rect 291162 95662 291240 95690
rect 291106 95639 291162 95648
rect 290924 93764 290976 93770
rect 290924 93706 290976 93712
rect 289818 76800 289874 76809
rect 289818 76735 289874 76744
rect 289266 75168 289322 75177
rect 289266 75103 289322 75112
rect 289818 72448 289874 72457
rect 289818 72383 289874 72392
rect 289084 50380 289136 50386
rect 289084 50322 289136 50328
rect 287060 35284 287112 35290
rect 287060 35226 287112 35232
rect 285678 24168 285734 24177
rect 285678 24103 285734 24112
rect 285692 16574 285720 24103
rect 287072 16574 287100 35226
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 284944 10396 284996 10402
rect 284944 10338 284996 10344
rect 284956 490 284984 10338
rect 285232 598 285444 626
rect 285232 490 285260 598
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 462 285260 490
rect 285416 480 285444 598
rect 286612 480 286640 16546
rect 287348 490 287376 16546
rect 288990 11656 289046 11665
rect 288990 11591 289046 11600
rect 287624 598 287836 626
rect 287624 490 287652 598
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 462 287652 490
rect 287808 480 287836 598
rect 289004 480 289032 11591
rect 289832 490 289860 72383
rect 291212 42090 291240 95662
rect 291292 95124 291344 95130
rect 291292 95066 291344 95072
rect 291200 42084 291252 42090
rect 291200 42026 291252 42032
rect 291200 40792 291252 40798
rect 291200 40734 291252 40740
rect 291212 3482 291240 40734
rect 291304 4826 291332 95066
rect 295996 93838 296024 96084
rect 295984 93832 296036 93838
rect 295984 93774 296036 93780
rect 299478 91760 299534 91769
rect 299478 91695 299534 91704
rect 298742 89040 298798 89049
rect 298742 88975 298798 88984
rect 295984 83496 296036 83502
rect 295984 83438 296036 83444
rect 295340 25628 295392 25634
rect 295340 25570 295392 25576
rect 295352 16574 295380 25570
rect 295352 16546 295656 16574
rect 292578 13016 292634 13025
rect 292578 12951 292634 12960
rect 291292 4820 291344 4826
rect 291292 4762 291344 4768
rect 291212 3454 291424 3482
rect 290016 598 290228 626
rect 290016 490 290044 598
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289832 462 290044 490
rect 290200 480 290228 598
rect 291396 480 291424 3454
rect 292592 480 292620 12951
rect 294878 3496 294934 3505
rect 293684 3460 293736 3466
rect 294878 3431 294934 3440
rect 293684 3402 293736 3408
rect 293696 480 293724 3402
rect 294892 480 294920 3431
rect 295628 490 295656 16546
rect 295996 3466 296024 83438
rect 296718 26888 296774 26897
rect 296718 26823 296774 26832
rect 296732 16574 296760 26823
rect 296732 16546 297312 16574
rect 295984 3460 296036 3466
rect 295984 3402 296036 3408
rect 295904 598 296116 626
rect 295904 490 295932 598
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 462 295932 490
rect 296088 480 296116 598
rect 297284 480 297312 16546
rect 298098 11656 298154 11665
rect 298098 11591 298154 11600
rect 298112 490 298140 11591
rect 298756 3330 298784 88975
rect 299492 3482 299520 91695
rect 301148 89690 301176 100558
rect 301318 100535 301374 100544
rect 301502 99648 301558 99657
rect 301502 99583 301558 99592
rect 301410 97336 301466 97345
rect 301410 97271 301466 97280
rect 301318 96656 301374 96665
rect 301318 96591 301374 96600
rect 301332 95169 301360 96591
rect 301318 95160 301374 95169
rect 301318 95095 301374 95104
rect 301424 95033 301452 97271
rect 301516 95198 301544 99583
rect 303618 99376 303674 99385
rect 303618 99311 303674 99320
rect 302238 98560 302294 98569
rect 302238 98495 302294 98504
rect 301504 95192 301556 95198
rect 301504 95134 301556 95140
rect 301410 95024 301466 95033
rect 301410 94959 301466 94968
rect 302252 93673 302280 98495
rect 302238 93664 302294 93673
rect 302238 93599 302294 93608
rect 303632 92478 303660 99311
rect 303620 92472 303672 92478
rect 303620 92414 303672 92420
rect 303724 91050 303752 101510
rect 303816 93770 303844 103486
rect 303896 96620 303948 96626
rect 303896 96562 303948 96568
rect 303908 96393 303936 96562
rect 303894 96384 303950 96393
rect 303894 96319 303950 96328
rect 303804 93764 303856 93770
rect 303804 93706 303856 93712
rect 303712 91044 303764 91050
rect 303712 90986 303764 90992
rect 304262 90400 304318 90409
rect 304262 90335 304318 90344
rect 301136 89684 301188 89690
rect 301136 89626 301188 89632
rect 299570 73808 299626 73817
rect 299570 73743 299626 73752
rect 299584 3602 299612 73743
rect 304276 6186 304304 90335
rect 311898 65512 311954 65521
rect 311898 65447 311954 65456
rect 307758 33824 307814 33833
rect 307758 33759 307814 33768
rect 304264 6180 304316 6186
rect 304264 6122 304316 6128
rect 303160 4888 303212 4894
rect 303160 4830 303212 4836
rect 299572 3596 299624 3602
rect 299572 3538 299624 3544
rect 300768 3596 300820 3602
rect 300768 3538 300820 3544
rect 299492 3454 299704 3482
rect 298744 3324 298796 3330
rect 298744 3266 298796 3272
rect 298296 598 298508 626
rect 298296 490 298324 598
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 462 298324 490
rect 298480 480 298508 598
rect 299676 480 299704 3454
rect 300780 480 300808 3538
rect 301964 3324 302016 3330
rect 301964 3266 302016 3272
rect 301976 480 302004 3266
rect 303172 480 303200 4830
rect 307772 3534 307800 33759
rect 310518 29608 310574 29617
rect 310518 29543 310574 29552
rect 310532 16574 310560 29543
rect 311912 16574 311940 65447
rect 310532 16546 311480 16574
rect 311912 16546 312216 16574
rect 310242 8936 310298 8945
rect 310242 8871 310298 8880
rect 307760 3528 307812 3534
rect 309048 3528 309100 3534
rect 307760 3470 307812 3476
rect 307942 3496 307998 3505
rect 304356 3460 304408 3466
rect 304356 3402 304408 3408
rect 306748 3460 306800 3466
rect 309048 3470 309100 3476
rect 307942 3431 307998 3440
rect 306748 3402 306800 3408
rect 304368 480 304396 3402
rect 305552 2168 305604 2174
rect 305552 2110 305604 2116
rect 305564 480 305592 2110
rect 306760 480 306788 3402
rect 307956 480 307984 3431
rect 309060 480 309088 3470
rect 310256 480 310284 8871
rect 311452 480 311480 16546
rect 312188 490 312216 16546
rect 314660 14476 314712 14482
rect 314660 14418 314712 14424
rect 313830 7032 313886 7041
rect 313830 6967 313886 6976
rect 312464 598 312676 626
rect 312464 490 312492 598
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 462 312492 490
rect 312648 480 312676 598
rect 313844 480 313872 6967
rect 314672 490 314700 14418
rect 317326 4040 317382 4049
rect 317326 3975 317382 3984
rect 316224 3324 316276 3330
rect 316224 3266 316276 3272
rect 314856 598 315068 626
rect 314856 490 314884 598
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 462 314884 490
rect 315040 480 315068 598
rect 316236 480 316264 3266
rect 317340 480 317368 3975
rect 317432 3466 317460 320719
rect 324412 307828 324464 307834
rect 324412 307770 324464 307776
rect 322940 257372 322992 257378
rect 322940 257314 322992 257320
rect 317512 250504 317564 250510
rect 317512 250446 317564 250452
rect 317524 132394 317552 250446
rect 321652 243568 321704 243574
rect 321652 243510 321704 243516
rect 320272 241528 320324 241534
rect 320272 241470 320324 241476
rect 318892 231124 318944 231130
rect 318892 231066 318944 231072
rect 317602 213208 317658 213217
rect 317602 213143 317658 213152
rect 317616 162858 317644 213143
rect 318798 203552 318854 203561
rect 318798 203487 318854 203496
rect 317696 179920 317748 179926
rect 317696 179862 317748 179868
rect 317604 162852 317656 162858
rect 317604 162794 317656 162800
rect 317708 146266 317736 179862
rect 317696 146260 317748 146266
rect 317696 146202 317748 146208
rect 317512 132388 317564 132394
rect 317512 132330 317564 132336
rect 318812 16574 318840 203487
rect 318904 120086 318932 231066
rect 318982 220144 319038 220153
rect 318982 220079 319038 220088
rect 318996 130422 319024 220079
rect 320178 191040 320234 191049
rect 320178 190975 320234 190984
rect 319076 178696 319128 178702
rect 319076 178638 319128 178644
rect 319088 161430 319116 178638
rect 319076 161424 319128 161430
rect 319076 161366 319128 161372
rect 318984 130416 319036 130422
rect 318984 130358 319036 130364
rect 318892 120080 318944 120086
rect 318892 120022 318944 120028
rect 318812 16546 319760 16574
rect 317420 3460 317472 3466
rect 317420 3402 317472 3408
rect 318522 2000 318578 2009
rect 318522 1935 318578 1944
rect 318536 480 318564 1935
rect 319732 480 319760 16546
rect 320192 3330 320220 190975
rect 320284 149054 320312 241470
rect 321560 234660 321612 234666
rect 321560 234602 321612 234608
rect 320364 199504 320416 199510
rect 320364 199446 320416 199452
rect 320272 149048 320324 149054
rect 320272 148990 320324 148996
rect 320376 121446 320404 199446
rect 320454 181520 320510 181529
rect 320454 181455 320510 181464
rect 320468 168366 320496 181455
rect 320456 168360 320508 168366
rect 320456 168302 320508 168308
rect 320364 121440 320416 121446
rect 320364 121382 320416 121388
rect 321572 109002 321600 234602
rect 321664 133822 321692 243510
rect 322202 195256 322258 195265
rect 322202 195191 322258 195200
rect 321744 181484 321796 181490
rect 321744 181426 321796 181432
rect 321756 155854 321784 181426
rect 321744 155848 321796 155854
rect 321744 155790 321796 155796
rect 321652 133816 321704 133822
rect 321652 133758 321704 133764
rect 321560 108996 321612 109002
rect 321560 108938 321612 108944
rect 322216 3534 322244 195191
rect 322952 142118 322980 257314
rect 324318 218648 324374 218657
rect 324318 218583 324374 218592
rect 323030 205048 323086 205057
rect 323030 204983 323086 204992
rect 322940 142112 322992 142118
rect 322940 142054 322992 142060
rect 323044 102134 323072 204983
rect 323124 182844 323176 182850
rect 323124 182786 323176 182792
rect 323136 144906 323164 182786
rect 323214 180024 323270 180033
rect 323214 179959 323270 179968
rect 323228 166326 323256 179959
rect 323216 166320 323268 166326
rect 323216 166262 323268 166268
rect 323124 144900 323176 144906
rect 323124 144842 323176 144848
rect 323032 102128 323084 102134
rect 323032 102070 323084 102076
rect 324332 3534 324360 218583
rect 324424 122806 324452 307770
rect 324962 300928 325018 300937
rect 324962 300863 325018 300872
rect 324502 184240 324558 184249
rect 324502 184175 324558 184184
rect 324516 153202 324544 184175
rect 324504 153196 324556 153202
rect 324504 153138 324556 153144
rect 324412 122800 324464 122806
rect 324412 122742 324464 122748
rect 324976 78674 325004 300863
rect 325700 272536 325752 272542
rect 325700 272478 325752 272484
rect 325712 124098 325740 272478
rect 325790 230616 325846 230625
rect 325790 230551 325846 230560
rect 325700 124092 325752 124098
rect 325700 124034 325752 124040
rect 325804 111790 325832 230551
rect 325884 192568 325936 192574
rect 325884 192510 325936 192516
rect 325896 164218 325924 192510
rect 325884 164212 325936 164218
rect 325884 164154 325936 164160
rect 325792 111784 325844 111790
rect 325792 111726 325844 111732
rect 324964 78668 325016 78674
rect 324964 78610 325016 78616
rect 325700 78668 325752 78674
rect 325700 78610 325752 78616
rect 324410 47560 324466 47569
rect 324410 47495 324466 47504
rect 322204 3528 322256 3534
rect 320914 3496 320970 3505
rect 320914 3431 320970 3440
rect 322110 3496 322166 3505
rect 322204 3470 322256 3476
rect 323308 3528 323360 3534
rect 323308 3470 323360 3476
rect 324320 3528 324372 3534
rect 324320 3470 324372 3476
rect 322110 3431 322166 3440
rect 320180 3324 320232 3330
rect 320180 3266 320232 3272
rect 320928 480 320956 3431
rect 322124 480 322152 3431
rect 323320 480 323348 3470
rect 324424 480 324452 47495
rect 325712 16574 325740 78610
rect 327092 16574 327120 368455
rect 327172 273964 327224 273970
rect 327172 273906 327224 273912
rect 327184 132462 327212 273906
rect 328458 267064 328514 267073
rect 328458 266999 328514 267008
rect 327264 253224 327316 253230
rect 327264 253166 327316 253172
rect 327172 132456 327224 132462
rect 327172 132398 327224 132404
rect 327276 124166 327304 253166
rect 327354 186960 327410 186969
rect 327354 186895 327410 186904
rect 327368 147626 327396 186895
rect 327356 147620 327408 147626
rect 327356 147562 327408 147568
rect 328472 125594 328500 266999
rect 329932 242208 329984 242214
rect 329932 242150 329984 242156
rect 328552 229764 328604 229770
rect 328552 229706 328604 229712
rect 328564 137970 328592 229706
rect 329838 200696 329894 200705
rect 329838 200631 329894 200640
rect 328552 137964 328604 137970
rect 328552 137906 328604 137912
rect 328460 125588 328512 125594
rect 328460 125530 328512 125536
rect 327264 124160 327316 124166
rect 327264 124102 327316 124108
rect 329852 16574 329880 200631
rect 329944 131102 329972 242150
rect 329932 131096 329984 131102
rect 329932 131038 329984 131044
rect 325712 16546 326384 16574
rect 327092 16546 328040 16574
rect 329852 16546 330432 16574
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 325620 480 325648 3470
rect 326356 490 326384 16546
rect 326632 598 326844 626
rect 326632 490 326660 598
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 462 326660 490
rect 326816 480 326844 598
rect 328012 480 328040 16546
rect 329194 4856 329250 4865
rect 329194 4791 329250 4800
rect 329208 480 329236 4791
rect 330404 480 330432 16546
rect 331232 490 331260 372574
rect 582378 365120 582434 365129
rect 582378 365055 582434 365064
rect 580172 352572 580224 352578
rect 580172 352514 580224 352520
rect 580184 351937 580212 352514
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 340878 350568 340934 350577
rect 340878 350503 340934 350512
rect 338118 343768 338174 343777
rect 338118 343703 338174 343712
rect 335360 335368 335412 335374
rect 335360 335310 335412 335316
rect 333978 325000 334034 325009
rect 333978 324935 334034 324944
rect 331312 267776 331364 267782
rect 331312 267718 331364 267724
rect 331324 155922 331352 267718
rect 331404 233300 331456 233306
rect 331404 233242 331456 233248
rect 331312 155916 331364 155922
rect 331312 155858 331364 155864
rect 331416 133890 331444 233242
rect 332690 228304 332746 228313
rect 332690 228239 332746 228248
rect 332598 207632 332654 207641
rect 332598 207567 332654 207576
rect 331404 133884 331456 133890
rect 331404 133826 331456 133832
rect 332612 3534 332640 207567
rect 332704 154494 332732 228239
rect 332692 154488 332744 154494
rect 332692 154430 332744 154436
rect 333992 16574 334020 324935
rect 334072 249076 334124 249082
rect 334072 249018 334124 249024
rect 334084 96626 334112 249018
rect 334072 96620 334124 96626
rect 334072 96562 334124 96568
rect 333992 16546 334664 16574
rect 332600 3528 332652 3534
rect 332600 3470 332652 3476
rect 333888 3528 333940 3534
rect 333888 3470 333940 3476
rect 332692 2984 332744 2990
rect 332692 2926 332744 2932
rect 331416 598 331628 626
rect 331416 490 331444 598
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 462 331444 490
rect 331600 480 331628 598
rect 332704 480 332732 2926
rect 333900 480 333928 3470
rect 334636 490 334664 16546
rect 335372 2990 335400 335310
rect 335544 217320 335596 217326
rect 335544 217262 335596 217268
rect 335450 211848 335506 211857
rect 335450 211783 335506 211792
rect 335464 16574 335492 211783
rect 335556 154562 335584 217262
rect 336738 215384 336794 215393
rect 336738 215319 336794 215328
rect 335544 154556 335596 154562
rect 335544 154498 335596 154504
rect 336752 128314 336780 215319
rect 336740 128308 336792 128314
rect 336740 128250 336792 128256
rect 335464 16546 336320 16574
rect 335360 2984 335412 2990
rect 335360 2926 335412 2932
rect 334912 598 335124 626
rect 334912 490 334940 598
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 462 334940 490
rect 335096 480 335124 598
rect 336292 480 336320 16546
rect 338132 3534 338160 343703
rect 339498 338192 339554 338201
rect 339498 338127 339554 338136
rect 338672 4820 338724 4826
rect 338672 4762 338724 4768
rect 337476 3528 337528 3534
rect 337476 3470 337528 3476
rect 338120 3528 338172 3534
rect 338120 3470 338172 3476
rect 337488 480 337516 3470
rect 338684 480 338712 4762
rect 339512 490 339540 338127
rect 339590 309224 339646 309233
rect 339590 309159 339646 309168
rect 339604 135250 339632 309159
rect 339592 135244 339644 135250
rect 339592 135186 339644 135192
rect 340892 16574 340920 350503
rect 582392 345681 582420 365055
rect 582378 345672 582434 345681
rect 582378 345607 582434 345616
rect 357440 340944 357492 340950
rect 357440 340886 357492 340892
rect 353298 222864 353354 222873
rect 353298 222799 353354 222808
rect 342258 214568 342314 214577
rect 342258 214503 342314 214512
rect 342272 16574 342300 214503
rect 345018 206272 345074 206281
rect 345018 206207 345074 206216
rect 345032 16574 345060 206207
rect 351918 199336 351974 199345
rect 351918 199271 351974 199280
rect 347044 17332 347096 17338
rect 347044 17274 347096 17280
rect 340892 16546 341012 16574
rect 342272 16546 342944 16574
rect 345032 16546 345336 16574
rect 339696 598 339908 626
rect 339696 490 339724 598
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 462 339724 490
rect 339880 480 339908 598
rect 340984 480 341012 16546
rect 342168 6180 342220 6186
rect 342168 6122 342220 6128
rect 342180 480 342208 6122
rect 342916 490 342944 16546
rect 344558 3360 344614 3369
rect 344558 3295 344614 3304
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 480 344600 3295
rect 345308 490 345336 16546
rect 346952 3324 347004 3330
rect 346952 3266 347004 3272
rect 345584 598 345796 626
rect 345584 490 345612 598
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 462 345612 490
rect 345768 480 345796 598
rect 346964 480 346992 3266
rect 347056 3126 347084 17274
rect 351642 3632 351698 3641
rect 351642 3567 351698 3576
rect 350448 3528 350500 3534
rect 348054 3496 348110 3505
rect 350448 3470 350500 3476
rect 348054 3431 348110 3440
rect 347044 3120 347096 3126
rect 347044 3062 347096 3068
rect 348068 480 348096 3431
rect 349252 3120 349304 3126
rect 349252 3062 349304 3068
rect 349264 480 349292 3062
rect 350460 480 350488 3470
rect 351656 480 351684 3567
rect 351932 3330 351960 199271
rect 353312 3534 353340 222799
rect 356058 221504 356114 221513
rect 356058 221439 356114 221448
rect 353300 3528 353352 3534
rect 353300 3470 353352 3476
rect 356072 3369 356100 221439
rect 357452 3505 357480 340886
rect 582378 334112 582434 334121
rect 582378 334047 582434 334056
rect 360200 325712 360252 325718
rect 360200 325654 360252 325660
rect 358818 196616 358874 196625
rect 358818 196551 358874 196560
rect 358832 3641 358860 196551
rect 360212 4826 360240 325654
rect 574742 299568 574798 299577
rect 574742 299503 574798 299512
rect 522304 251864 522356 251870
rect 522304 251806 522356 251812
rect 522316 167006 522344 251806
rect 574756 179382 574784 299503
rect 580262 272232 580318 272241
rect 580262 272167 580318 272176
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 240145 580212 245511
rect 580276 240786 580304 272167
rect 580264 240780 580316 240786
rect 580264 240722 580316 240728
rect 580170 240136 580226 240145
rect 580170 240071 580226 240080
rect 580908 225072 580960 225078
rect 580908 225014 580960 225020
rect 574744 179376 574796 179382
rect 574744 179318 574796 179324
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 522304 167000 522356 167006
rect 522304 166942 522356 166948
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580920 126041 580948 225014
rect 580906 126032 580962 126041
rect 580906 125967 580962 125976
rect 582392 16574 582420 334047
rect 582564 296744 582616 296750
rect 582564 296686 582616 296692
rect 582472 295384 582524 295390
rect 582472 295326 582524 295332
rect 582484 19825 582512 295326
rect 582576 73001 582604 296686
rect 582668 276010 582696 471407
rect 583022 418296 583078 418305
rect 583022 418231 583078 418240
rect 582838 378448 582894 378457
rect 582838 378383 582894 378392
rect 582746 298752 582802 298761
rect 582746 298687 582802 298696
rect 582656 276004 582708 276010
rect 582656 275946 582708 275952
rect 582656 262880 582708 262886
rect 582656 262822 582708 262828
rect 582668 232393 582696 262822
rect 582760 237289 582788 298687
rect 582852 282878 582880 378383
rect 582930 302288 582986 302297
rect 582930 302223 582986 302232
rect 582840 282872 582892 282878
rect 582840 282814 582892 282820
rect 582838 237960 582894 237969
rect 582838 237895 582894 237904
rect 582746 237280 582802 237289
rect 582746 237215 582802 237224
rect 582654 232384 582710 232393
rect 582654 232319 582710 232328
rect 582656 226364 582708 226370
rect 582656 226306 582708 226312
rect 582562 72992 582618 73001
rect 582562 72927 582618 72936
rect 582470 19816 582526 19825
rect 582470 19751 582526 19760
rect 582392 16546 582604 16574
rect 360200 4820 360252 4826
rect 360200 4762 360252 4768
rect 358818 3632 358874 3641
rect 358818 3567 358874 3576
rect 582196 3528 582248 3534
rect 357438 3496 357494 3505
rect 582196 3470 582248 3476
rect 582576 3482 582604 16546
rect 582668 6633 582696 226306
rect 582748 224256 582800 224262
rect 582748 224198 582800 224204
rect 582760 33153 582788 224198
rect 582852 46345 582880 237895
rect 582944 112849 582972 302223
rect 583036 289105 583064 418231
rect 583390 404968 583446 404977
rect 583390 404903 583446 404912
rect 583298 325272 583354 325281
rect 583298 325207 583354 325216
rect 583114 312080 583170 312089
rect 583114 312015 583170 312024
rect 583022 289096 583078 289105
rect 583022 289031 583078 289040
rect 583022 284336 583078 284345
rect 583022 284271 583078 284280
rect 583036 258913 583064 284271
rect 583128 266354 583156 312015
rect 583208 294024 583260 294030
rect 583208 293966 583260 293972
rect 583116 266348 583168 266354
rect 583116 266290 583168 266296
rect 583114 264208 583170 264217
rect 583114 264143 583170 264152
rect 583022 258904 583078 258913
rect 583022 258839 583078 258848
rect 583024 225004 583076 225010
rect 583024 224946 583076 224952
rect 582930 112840 582986 112849
rect 582930 112775 582986 112784
rect 583036 59673 583064 224946
rect 583128 99521 583156 264143
rect 583220 139369 583248 293966
rect 583312 247722 583340 325207
rect 583404 291825 583432 404903
rect 583482 305008 583538 305017
rect 583482 304943 583538 304952
rect 583390 291816 583446 291825
rect 583390 291751 583446 291760
rect 583392 278044 583444 278050
rect 583392 277986 583444 277992
rect 583300 247716 583352 247722
rect 583300 247658 583352 247664
rect 583298 229800 583354 229809
rect 583298 229735 583354 229744
rect 583206 139360 583262 139369
rect 583206 139295 583262 139304
rect 583114 99512 583170 99521
rect 583114 99447 583170 99456
rect 583312 86193 583340 229735
rect 583404 152697 583432 277986
rect 583496 219337 583524 304943
rect 583666 303648 583722 303657
rect 583666 303583 583722 303592
rect 583576 278792 583628 278798
rect 583576 278734 583628 278740
rect 583588 225078 583616 278734
rect 583576 225072 583628 225078
rect 583576 225014 583628 225020
rect 583482 219328 583538 219337
rect 583482 219263 583538 219272
rect 583482 208992 583538 209001
rect 583482 208927 583538 208936
rect 583390 152688 583446 152697
rect 583390 152623 583446 152632
rect 583298 86184 583354 86193
rect 583298 86119 583354 86128
rect 583022 59664 583078 59673
rect 583022 59599 583078 59608
rect 582838 46336 582894 46345
rect 582838 46271 582894 46280
rect 582746 33144 582802 33153
rect 582746 33079 582802 33088
rect 582654 6624 582710 6633
rect 582654 6559 582710 6568
rect 583496 3534 583524 208927
rect 583574 203008 583630 203017
rect 583574 202943 583630 202952
rect 583484 3528 583536 3534
rect 357438 3431 357494 3440
rect 356058 3360 356114 3369
rect 351920 3324 351972 3330
rect 356058 3295 356114 3304
rect 351920 3266 351972 3272
rect 581000 3052 581052 3058
rect 581000 2994 581052 3000
rect 581012 480 581040 2994
rect 582208 480 582236 3470
rect 582576 3454 583432 3482
rect 583484 3470 583536 3476
rect 583404 480 583432 3454
rect 583588 3058 583616 202943
rect 583680 193089 583708 303583
rect 583760 298172 583812 298178
rect 583760 298114 583812 298120
rect 583772 206281 583800 298114
rect 583758 206272 583814 206281
rect 583758 206207 583814 206216
rect 583666 193080 583722 193089
rect 583666 193015 583722 193024
rect 583576 3052 583628 3058
rect 583576 2994 583628 3000
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 2778 658144 2834 658200
rect 2778 579944 2834 580000
rect 3238 566888 3294 566944
rect 3514 671200 3570 671256
rect 3514 632068 3516 632088
rect 3516 632068 3568 632088
rect 3568 632068 3570 632088
rect 3514 632032 3570 632068
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 3514 553852 3570 553888
rect 3514 553832 3516 553852
rect 3516 553832 3568 553852
rect 3568 553832 3570 553852
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 2778 501744 2834 501800
rect 3330 475632 3386 475688
rect 2778 462596 2834 462632
rect 2778 462576 2780 462596
rect 2780 462576 2832 462596
rect 2832 462576 2834 462596
rect 3146 449520 3202 449576
rect 3422 423580 3424 423600
rect 3424 423580 3476 423600
rect 3476 423580 3478 423600
rect 3422 423544 3478 423580
rect 3422 410488 3478 410544
rect 2778 397432 2834 397488
rect 7562 382880 7618 382936
rect 3146 371320 3202 371376
rect 3422 358400 3478 358456
rect 3146 345344 3202 345400
rect 7562 327256 7618 327312
rect 4066 319232 4122 319288
rect 3422 306176 3478 306232
rect 2778 293120 2834 293176
rect 3422 267144 3478 267200
rect 3422 254088 3478 254144
rect 3422 241032 3478 241088
rect 4802 222264 4858 222320
rect 3330 214920 3386 214976
rect 3514 206216 3570 206272
rect 3422 201864 3478 201920
rect 3238 162832 3294 162888
rect 3514 188808 3570 188864
rect 3514 149776 3570 149832
rect 3514 136720 3570 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 4066 76472 4122 76528
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 2778 45500 2780 45520
rect 2780 45500 2832 45520
rect 2832 45500 2834 45520
rect 2778 45464 2834 45500
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 6826 18536 6882 18592
rect 53654 590688 53710 590744
rect 17222 391176 17278 391232
rect 33782 386960 33838 387016
rect 17222 328480 17278 328536
rect 16486 77832 16542 77888
rect 13726 69536 13782 69592
rect 15106 53080 15162 53136
rect 21362 326168 21418 326224
rect 36542 197920 36598 197976
rect 22006 83408 22062 83464
rect 19246 68176 19302 68232
rect 17866 48864 17922 48920
rect 34426 82048 34482 82104
rect 22742 77968 22798 78024
rect 19430 3304 19486 3360
rect 26146 59880 26202 59936
rect 24766 21256 24822 21312
rect 33046 55936 33102 55992
rect 29642 37848 29698 37904
rect 28906 30912 28962 30968
rect 33782 39208 33838 39264
rect 35806 79464 35862 79520
rect 38566 46144 38622 46200
rect 41326 66816 41382 66872
rect 42706 44784 42762 44840
rect 43994 239400 44050 239456
rect 48134 62736 48190 62792
rect 43902 25472 43958 25528
rect 46846 22616 46902 22672
rect 50894 239536 50950 239592
rect 50802 227568 50858 227624
rect 50894 79328 50950 79384
rect 52090 236544 52146 236600
rect 53654 445984 53710 446040
rect 55034 445848 55090 445904
rect 53562 224848 53618 224904
rect 53746 289992 53802 290048
rect 55034 219136 55090 219192
rect 54942 198600 54998 198656
rect 53746 72392 53802 72448
rect 53746 64096 53802 64152
rect 52366 33768 52422 33824
rect 48226 1944 48282 2000
rect 56322 231104 56378 231160
rect 56414 217912 56470 217968
rect 61934 590824 61990 590880
rect 58990 357992 59046 358048
rect 57794 241440 57850 241496
rect 56506 71168 56562 71224
rect 55126 29552 55182 29608
rect 57794 35128 57850 35184
rect 66074 581576 66130 581632
rect 61934 393252 61936 393272
rect 61936 393252 61988 393272
rect 61988 393252 61990 393272
rect 61934 393216 61990 393252
rect 59082 230424 59138 230480
rect 59174 75248 59230 75304
rect 57886 32408 57942 32464
rect 60462 237904 60518 237960
rect 60554 216552 60610 216608
rect 61658 313384 61714 313440
rect 65982 572872 66038 572928
rect 65522 564440 65578 564496
rect 66810 588240 66866 588296
rect 66258 586508 66260 586528
rect 66260 586508 66312 586528
rect 66312 586508 66314 586528
rect 66258 586472 66314 586508
rect 66810 582412 66866 582448
rect 66810 582392 66812 582412
rect 66812 582392 66864 582412
rect 66864 582392 66866 582412
rect 66810 579692 66866 579728
rect 66810 579672 66812 579692
rect 66812 579672 66864 579692
rect 66864 579672 66866 579692
rect 66902 575592 66958 575648
rect 67454 575320 67510 575376
rect 66442 571784 66498 571840
rect 67362 570152 67418 570208
rect 66902 568792 66958 568848
rect 66902 567432 66958 567488
rect 66810 564340 66812 564360
rect 66812 564340 66864 564360
rect 66864 564340 66866 564360
rect 66810 564304 66866 564340
rect 66810 561740 66866 561776
rect 66810 561720 66812 561740
rect 66812 561720 66864 561740
rect 66864 561720 66866 561740
rect 66534 560496 66590 560552
rect 66534 559136 66590 559192
rect 66902 556280 66958 556336
rect 66626 554920 66682 554976
rect 66534 553696 66590 553752
rect 66442 549616 66498 549672
rect 66534 548256 66590 548312
rect 66626 547576 66682 547632
rect 66166 546352 66222 546408
rect 66810 544040 66866 544096
rect 66810 542680 66866 542736
rect 65982 448568 66038 448624
rect 64602 385600 64658 385656
rect 63222 362208 63278 362264
rect 64786 350784 64842 350840
rect 64602 337320 64658 337376
rect 61842 193160 61898 193216
rect 63314 223488 63370 223544
rect 63222 199960 63278 200016
rect 62026 69672 62082 69728
rect 60646 65456 60702 65512
rect 59266 54440 59322 54496
rect 62026 50224 62082 50280
rect 64694 335552 64750 335608
rect 65982 388864 66038 388920
rect 66534 437688 66590 437744
rect 66810 435240 66866 435296
rect 66442 433064 66498 433120
rect 66810 430888 66866 430944
rect 66810 428440 66866 428496
rect 66810 426264 66866 426320
rect 66810 424088 66866 424144
rect 66810 421912 66866 421968
rect 67086 541728 67142 541784
rect 67546 566752 67602 566808
rect 67730 589872 67786 589928
rect 72974 699760 73030 699816
rect 72422 590960 72478 591016
rect 71042 590824 71098 590880
rect 73618 590688 73674 590744
rect 77022 590688 77078 590744
rect 75642 588784 75698 588840
rect 83462 592048 83518 592104
rect 82542 590824 82598 590880
rect 81346 590552 81402 590608
rect 82634 590688 82690 590744
rect 83738 590960 83794 591016
rect 86866 590960 86922 591016
rect 86958 588784 87014 588840
rect 88982 590552 89038 590608
rect 88062 588512 88118 588568
rect 67730 585792 67786 585848
rect 88982 582936 89038 582992
rect 67730 578312 67786 578368
rect 67638 558864 67694 558920
rect 67454 552200 67510 552256
rect 66994 439864 67050 439920
rect 66902 419500 66904 419520
rect 66904 419500 66956 419520
rect 66956 419500 66958 419520
rect 66902 419464 66958 419500
rect 66442 417288 66498 417344
rect 66810 415112 66866 415168
rect 66258 406156 66314 406192
rect 66258 406136 66260 406156
rect 66260 406136 66312 406156
rect 66312 406136 66314 406156
rect 66258 403688 66314 403744
rect 66258 401548 66260 401568
rect 66260 401548 66312 401568
rect 66312 401548 66314 401568
rect 66258 401512 66314 401548
rect 66442 399336 66498 399392
rect 66994 396888 67050 396944
rect 66810 392536 66866 392592
rect 66166 388320 66222 388376
rect 66074 360848 66130 360904
rect 66074 312024 66130 312080
rect 67178 326712 67234 326768
rect 66902 324808 66958 324864
rect 66810 323720 66866 323776
rect 66442 320456 66498 320512
rect 66810 319368 66866 319424
rect 66902 318280 66958 318336
rect 66810 317500 66812 317520
rect 66812 317500 66864 317520
rect 66864 317500 66866 317520
rect 66810 317464 66866 317500
rect 67454 412664 67510 412720
rect 67362 338408 67418 338464
rect 67362 326984 67418 327040
rect 67362 321544 67418 321600
rect 67270 316376 67326 316432
rect 66810 315288 66866 315344
rect 66902 314200 66958 314256
rect 66810 313112 66866 313168
rect 66442 310936 66498 310992
rect 66810 309848 66866 309904
rect 66718 307944 66774 308000
rect 66902 305768 66958 305824
rect 66902 304680 66958 304736
rect 66258 303628 66260 303648
rect 66260 303628 66312 303648
rect 66312 303628 66314 303648
rect 66258 303592 66314 303628
rect 66810 302504 66866 302560
rect 66810 301416 66866 301472
rect 66258 300600 66314 300656
rect 66810 299512 66866 299568
rect 66442 296248 66498 296304
rect 66258 294092 66314 294128
rect 66258 294072 66260 294092
rect 66260 294072 66312 294092
rect 66312 294072 66314 294092
rect 66902 292984 66958 293040
rect 66810 292168 66866 292224
rect 66810 289992 66866 290048
rect 66258 288904 66314 288960
rect 66810 287816 66866 287872
rect 66810 285676 66812 285696
rect 66812 285676 66864 285696
rect 66864 285676 66866 285696
rect 66810 285640 66866 285676
rect 66626 283736 66682 283792
rect 66350 282648 66406 282704
rect 66810 280472 66866 280528
rect 66626 279384 66682 279440
rect 66258 277208 66314 277264
rect 66166 276120 66222 276176
rect 66074 256264 66130 256320
rect 64694 234504 64750 234560
rect 64602 219272 64658 219328
rect 66810 272040 66866 272096
rect 66810 270952 66866 271008
rect 66442 269864 66498 269920
rect 66442 267708 66498 267744
rect 66442 267688 66444 267708
rect 66444 267688 66496 267708
rect 66496 267688 66498 267708
rect 66994 286728 67050 286784
rect 67086 284552 67142 284608
rect 67546 394712 67602 394768
rect 67822 576952 67878 577008
rect 68650 540776 68706 540832
rect 69662 535472 69718 535528
rect 70674 535472 70730 535528
rect 67822 445712 67878 445768
rect 68466 445712 68522 445768
rect 72422 448568 72478 448624
rect 71778 447208 71834 447264
rect 76746 538056 76802 538112
rect 76470 536696 76526 536752
rect 75918 535472 75974 535528
rect 76746 535472 76802 535528
rect 81438 461488 81494 461544
rect 82082 457408 82138 457464
rect 78678 445848 78734 445904
rect 84750 536016 84806 536072
rect 82726 456184 82782 456240
rect 84106 460128 84162 460184
rect 82082 445848 82138 445904
rect 86866 462848 86922 462904
rect 86222 449112 86278 449168
rect 85578 445984 85634 446040
rect 87050 457408 87106 457464
rect 88890 567248 88946 567284
rect 88890 567228 88892 567248
rect 88892 567228 88944 567248
rect 88944 567228 88946 567248
rect 89626 456048 89682 456104
rect 89902 585792 89958 585848
rect 89810 560088 89866 560144
rect 91098 581576 91154 581632
rect 91098 578856 91154 578912
rect 91098 577496 91154 577552
rect 91926 584568 91982 584624
rect 91834 583652 91836 583672
rect 91836 583652 91888 583672
rect 91888 583652 91890 583672
rect 91834 583616 91890 583652
rect 91190 576680 91246 576736
rect 91098 575048 91154 575104
rect 91098 573416 91154 573472
rect 91190 572056 91246 572112
rect 91098 571396 91154 571432
rect 91098 571376 91100 571396
rect 91100 571376 91152 571396
rect 91152 571376 91154 571396
rect 91098 570016 91154 570072
rect 92202 568656 92258 568712
rect 91098 565836 91100 565856
rect 91100 565836 91152 565856
rect 91152 565836 91154 565856
rect 91098 565800 91154 565836
rect 91742 564440 91798 564496
rect 91098 563100 91154 563136
rect 91098 563080 91100 563100
rect 91100 563080 91152 563100
rect 91152 563080 91154 563100
rect 91098 560904 91154 560960
rect 89994 545264 90050 545320
rect 91190 558184 91246 558240
rect 91190 556824 91246 556880
rect 91190 555464 91246 555520
rect 91190 552880 91246 552936
rect 91190 552084 91246 552120
rect 91190 552064 91192 552084
rect 91192 552064 91244 552084
rect 91244 552064 91246 552084
rect 91190 549344 91246 549400
rect 91282 547848 91338 547904
rect 91190 544040 91246 544096
rect 91190 542428 91246 542464
rect 91190 542408 91192 542428
rect 91192 542408 91244 542428
rect 91244 542408 91246 542428
rect 91190 541320 91246 541376
rect 91190 539708 91246 539744
rect 91190 539688 91192 539708
rect 91192 539688 91244 539708
rect 91244 539688 91246 539708
rect 91374 546488 91430 546544
rect 91006 458768 91062 458824
rect 91834 560088 91890 560144
rect 91742 451832 91798 451888
rect 91558 448568 91614 448624
rect 90132 444488 90188 444544
rect 93766 469784 93822 469840
rect 93122 460128 93178 460184
rect 95146 467064 95202 467120
rect 95882 455504 95938 455560
rect 95238 446392 95294 446448
rect 93858 445712 93914 445768
rect 94502 445712 94558 445768
rect 98642 588648 98698 588704
rect 97906 580896 97962 580952
rect 97906 580216 97962 580272
rect 101402 588784 101458 588840
rect 100666 462848 100722 462904
rect 98734 461488 98790 461544
rect 96618 445712 96674 445768
rect 97354 445712 97410 445768
rect 104254 459584 104310 459640
rect 104162 450472 104218 450528
rect 102138 445712 102194 445768
rect 107014 590824 107070 590880
rect 105542 445984 105598 446040
rect 106922 456048 106978 456104
rect 110418 592048 110474 592104
rect 108394 447752 108450 447808
rect 112442 590960 112498 591016
rect 110418 445712 110474 445768
rect 111154 445712 111210 445768
rect 109038 444624 109094 444680
rect 118698 585656 118754 585712
rect 116398 445848 116454 445904
rect 113178 445712 113234 445768
rect 114098 445712 114154 445768
rect 117318 445712 117374 445768
rect 123482 582936 123538 582992
rect 119020 444624 119076 444680
rect 68650 444216 68706 444272
rect 67730 442040 67786 442096
rect 67454 309032 67510 309088
rect 120630 419328 120686 419384
rect 120630 416744 120686 416800
rect 67822 410488 67878 410544
rect 68374 408312 68430 408368
rect 67822 389816 67878 389872
rect 69938 390360 69994 390416
rect 71870 390360 71926 390416
rect 72054 389000 72110 389056
rect 73066 389000 73122 389056
rect 70306 347928 70362 347984
rect 69386 331200 69442 331256
rect 68282 329024 68338 329080
rect 67638 322632 67694 322688
rect 68650 327120 68706 327176
rect 68558 326440 68614 326496
rect 70674 332560 70730 332616
rect 72974 334192 73030 334248
rect 74538 388864 74594 388920
rect 76562 387096 76618 387152
rect 74998 341400 75054 341456
rect 75734 327120 75790 327176
rect 70030 327004 70086 327040
rect 79966 388320 80022 388376
rect 76654 366288 76710 366344
rect 77942 355408 77998 355464
rect 77206 342352 77262 342408
rect 92754 390904 92810 390960
rect 85486 389000 85542 389056
rect 81346 369008 81402 369064
rect 79966 367648 80022 367704
rect 80702 339496 80758 339552
rect 84014 383016 84070 383072
rect 84106 374584 84162 374640
rect 83462 353504 83518 353560
rect 84014 353504 84070 353560
rect 85762 352552 85818 352608
rect 85578 351056 85634 351112
rect 85762 345072 85818 345128
rect 84106 330520 84162 330576
rect 83646 327664 83702 327720
rect 86314 333240 86370 333296
rect 89810 390360 89866 390416
rect 91282 390360 91338 390416
rect 90362 389000 90418 389056
rect 89626 358808 89682 358864
rect 88982 352552 89038 352608
rect 89442 338272 89498 338328
rect 87142 336776 87198 336832
rect 102598 390904 102654 390960
rect 110418 390904 110474 390960
rect 111154 390904 111210 390960
rect 100666 390496 100722 390552
rect 93766 388320 93822 388376
rect 91006 371320 91062 371376
rect 97354 390360 97410 390416
rect 95882 389000 95938 389056
rect 94502 369824 94558 369880
rect 93214 350648 93270 350704
rect 93766 350648 93822 350704
rect 90822 331336 90878 331392
rect 92754 334328 92810 334384
rect 98826 390360 98882 390416
rect 98642 368328 98698 368384
rect 100114 389816 100170 389872
rect 98642 367104 98698 367160
rect 95146 340992 95202 341048
rect 97906 339768 97962 339824
rect 98642 333240 98698 333296
rect 98550 332696 98606 332752
rect 99286 330384 99342 330440
rect 93858 327256 93914 327312
rect 77298 327120 77354 327176
rect 83922 327120 83978 327176
rect 105082 390360 105138 390416
rect 102598 389000 102654 389056
rect 105542 389000 105598 389056
rect 102046 360168 102102 360224
rect 101402 346432 101458 346488
rect 100758 341400 100814 341456
rect 102782 342216 102838 342272
rect 106554 390360 106610 390416
rect 105634 386960 105690 387016
rect 108026 390360 108082 390416
rect 108302 389272 108358 389328
rect 108302 388320 108358 388376
rect 108302 385600 108358 385656
rect 109498 390360 109554 390416
rect 107842 363024 107898 363080
rect 106922 352008 106978 352064
rect 105542 346976 105598 347032
rect 106186 342488 106242 342544
rect 107750 335416 107806 335472
rect 106922 330384 106978 330440
rect 114098 389272 114154 389328
rect 111798 389000 111854 389056
rect 112626 389000 112682 389056
rect 115938 390360 115994 390416
rect 112442 356632 112498 356688
rect 112442 353640 112498 353696
rect 110418 347792 110474 347848
rect 111706 347792 111762 347848
rect 108762 334056 108818 334112
rect 109958 331064 110014 331120
rect 111706 343712 111762 343768
rect 111798 339632 111854 339688
rect 113086 349152 113142 349208
rect 112442 335960 112498 336016
rect 114466 343848 114522 343904
rect 118698 389408 118754 389464
rect 117778 389172 117780 389192
rect 117780 389172 117832 389192
rect 117832 389172 117834 389192
rect 117778 389136 117834 389172
rect 120262 390360 120318 390416
rect 119342 386280 119398 386336
rect 117318 365608 117374 365664
rect 117318 364384 117374 364440
rect 116582 355272 116638 355328
rect 115938 349696 115994 349752
rect 115294 346568 115350 346624
rect 115294 331064 115350 331120
rect 115018 328480 115074 328536
rect 120814 419464 120870 419520
rect 120722 411032 120778 411088
rect 121182 410488 121238 410544
rect 123114 450472 123170 450528
rect 122746 430888 122802 430944
rect 121642 428440 121698 428496
rect 121550 396888 121606 396944
rect 121458 392536 121514 392592
rect 119434 374584 119490 374640
rect 121366 364520 121422 364576
rect 120722 360304 120778 360360
rect 119434 357448 119490 357504
rect 118606 340856 118662 340912
rect 123022 447752 123078 447808
rect 122930 424088 122986 424144
rect 123114 433064 123170 433120
rect 123114 428440 123170 428496
rect 123022 417288 123078 417344
rect 123022 412664 123078 412720
rect 122930 394712 122986 394768
rect 122838 378664 122894 378720
rect 123482 447616 123538 447672
rect 124126 439864 124182 439920
rect 124862 536696 124918 536752
rect 123666 437688 123722 437744
rect 123850 433064 123906 433120
rect 123206 421912 123262 421968
rect 124126 415148 124128 415168
rect 124128 415148 124180 415168
rect 124180 415148 124182 415168
rect 124126 415112 124182 415148
rect 124126 408312 124182 408368
rect 124126 406156 124182 406192
rect 124126 406136 124128 406156
rect 124128 406136 124180 406156
rect 124180 406136 124182 406156
rect 124034 403688 124090 403744
rect 124126 401548 124128 401568
rect 124128 401548 124180 401568
rect 124180 401548 124182 401568
rect 124126 401512 124182 401548
rect 123666 399336 123722 399392
rect 123666 394712 123722 394768
rect 121458 353368 121514 353424
rect 122746 353368 122802 353424
rect 122102 328480 122158 328536
rect 128266 446256 128322 446312
rect 128266 445848 128322 445904
rect 124862 345616 124918 345672
rect 125506 338136 125562 338192
rect 128266 363568 128322 363624
rect 126978 362208 127034 362264
rect 125690 357312 125746 357368
rect 126886 357312 126942 357368
rect 125690 356088 125746 356144
rect 129002 536016 129058 536072
rect 128542 446256 128598 446312
rect 128450 348372 128452 348392
rect 128452 348372 128504 348392
rect 128504 348372 128506 348392
rect 128450 348336 128506 348372
rect 129830 352552 129886 352608
rect 129830 351872 129886 351928
rect 130474 447208 130530 447264
rect 130474 365744 130530 365800
rect 130382 349832 130438 349888
rect 154118 702480 154174 702536
rect 582378 697176 582434 697232
rect 580262 670656 580318 670712
rect 580170 590960 580226 591016
rect 580170 589872 580226 589928
rect 580262 577632 580318 577688
rect 133786 401648 133842 401704
rect 131118 355272 131174 355328
rect 129738 329160 129794 329216
rect 132038 331472 132094 331528
rect 131486 329840 131542 329896
rect 137282 444488 137338 444544
rect 136638 388728 136694 388784
rect 579802 537784 579858 537840
rect 582470 683848 582526 683904
rect 582562 644000 582618 644056
rect 582378 536016 582434 536072
rect 582654 630808 582710 630864
rect 582746 617480 582802 617536
rect 582746 564304 582802 564360
rect 582470 524456 582526 524512
rect 580170 511284 580226 511320
rect 580170 511264 580172 511284
rect 580172 511264 580224 511284
rect 580224 511264 580226 511284
rect 582378 484608 582434 484664
rect 142158 425584 142214 425640
rect 137926 368464 137982 368520
rect 135902 355544 135958 355600
rect 136546 350512 136602 350568
rect 134522 349696 134578 349752
rect 133142 337320 133198 337376
rect 132590 336912 132646 336968
rect 132682 330112 132738 330168
rect 134154 330248 134210 330304
rect 133326 329976 133382 330032
rect 139398 337048 139454 337104
rect 145562 377304 145618 377360
rect 144918 353776 144974 353832
rect 145562 353776 145618 353832
rect 144826 353640 144882 353696
rect 144826 352552 144882 352608
rect 143446 332832 143502 332888
rect 144826 341128 144882 341184
rect 146206 340892 146208 340912
rect 146208 340892 146260 340912
rect 146260 340892 146262 340912
rect 146206 340856 146262 340892
rect 145378 335960 145434 336016
rect 146206 328480 146262 328536
rect 150346 340856 150402 340912
rect 147586 329976 147642 330032
rect 70030 326984 70032 327004
rect 70032 326984 70084 327004
rect 70084 326984 70086 327004
rect 142894 326984 142950 327040
rect 149058 329024 149114 329080
rect 148276 327664 148332 327720
rect 151174 356632 151230 356688
rect 151082 329024 151138 329080
rect 150714 327528 150770 327584
rect 152462 355408 152518 355464
rect 153842 346976 153898 347032
rect 153934 335552 153990 335608
rect 153658 328616 153714 328672
rect 151726 328480 151782 328536
rect 152830 327528 152886 327584
rect 154394 327256 154450 327312
rect 153106 326984 153162 327040
rect 154394 327020 154396 327040
rect 154396 327020 154448 327040
rect 154448 327020 154450 327040
rect 154394 326984 154450 327020
rect 68650 326168 68706 326224
rect 67638 309032 67694 309088
rect 67546 298424 67602 298480
rect 67546 295160 67602 295216
rect 67454 281560 67510 281616
rect 67362 278296 67418 278352
rect 67362 275304 67418 275360
rect 67086 274216 67142 274272
rect 66994 273128 67050 273184
rect 66810 265784 66866 265840
rect 66810 264696 66866 264752
rect 66442 263608 66498 263664
rect 66810 262520 66866 262576
rect 66810 261432 66866 261488
rect 66810 258440 66866 258496
rect 66442 257352 66498 257408
rect 66994 255992 67050 256048
rect 66442 255176 66498 255232
rect 66626 253000 66682 253056
rect 66810 248920 66866 248976
rect 66810 247832 66866 247888
rect 67270 246744 67326 246800
rect 67178 244568 67234 244624
rect 67178 241304 67234 241360
rect 67546 260344 67602 260400
rect 67270 221448 67326 221504
rect 66166 202816 66222 202872
rect 67730 306856 67786 306912
rect 154854 326848 154910 326904
rect 154670 276936 154726 276992
rect 155866 356632 155922 356688
rect 156142 349696 156198 349752
rect 155958 345616 156014 345672
rect 155958 318008 156014 318064
rect 154854 295568 154910 295624
rect 154762 264696 154818 264752
rect 155222 290400 155278 290456
rect 154854 261976 154910 262032
rect 68098 258712 68154 258768
rect 67914 250824 67970 250880
rect 67730 250008 67786 250064
rect 67638 233144 67694 233200
rect 69754 241868 69810 241904
rect 69754 241848 69756 241868
rect 69756 241848 69808 241868
rect 69808 241848 69810 241868
rect 69662 241712 69718 241768
rect 67730 226072 67786 226128
rect 70306 238584 70362 238640
rect 69662 216416 69718 216472
rect 71686 240352 71742 240408
rect 71778 234368 71834 234424
rect 74446 239536 74502 239592
rect 73158 238448 73214 238504
rect 73802 237904 73858 237960
rect 73802 220632 73858 220688
rect 75182 213832 75238 213888
rect 77206 239400 77262 239456
rect 77114 212336 77170 212392
rect 74538 205536 74594 205592
rect 79322 225936 79378 225992
rect 77390 214784 77446 214840
rect 73066 196560 73122 196616
rect 82956 241440 83012 241496
rect 84106 241440 84162 241496
rect 84750 239400 84806 239456
rect 84106 226208 84162 226264
rect 86866 204856 86922 204912
rect 85486 200912 85542 200968
rect 88982 220768 89038 220824
rect 88246 195200 88302 195256
rect 90914 228248 90970 228304
rect 89626 189624 89682 189680
rect 81346 188264 81402 188320
rect 92294 217232 92350 217288
rect 95238 212472 95294 212528
rect 95146 199280 95202 199336
rect 99286 213288 99342 213344
rect 101954 207712 102010 207768
rect 103334 231784 103390 231840
rect 103518 237224 103574 237280
rect 106922 239400 106978 239456
rect 107474 224712 107530 224768
rect 108302 230288 108358 230344
rect 107566 214648 107622 214704
rect 104898 213152 104954 213208
rect 104806 210976 104862 211032
rect 102046 200776 102102 200832
rect 112534 239400 112590 239456
rect 93766 186904 93822 186960
rect 79966 185544 80022 185600
rect 104806 183776 104862 183832
rect 101954 183640 102010 183696
rect 99470 182144 99526 182200
rect 101954 177520 102010 177576
rect 105450 179424 105506 179480
rect 104806 177520 104862 177576
rect 113178 232872 113234 232928
rect 114466 204040 114522 204096
rect 111706 188400 111762 188456
rect 117226 239808 117282 239864
rect 120078 235728 120134 235784
rect 118882 221992 118938 222048
rect 118606 202136 118662 202192
rect 124310 238312 124366 238368
rect 123482 228928 123538 228984
rect 126150 239944 126206 240000
rect 127070 237088 127126 237144
rect 126886 210840 126942 210896
rect 126794 209616 126850 209672
rect 125506 205400 125562 205456
rect 128358 236544 128414 236600
rect 129554 227296 129610 227352
rect 128266 206896 128322 206952
rect 129646 202272 129702 202328
rect 133694 198056 133750 198112
rect 135994 241984 136050 242040
rect 138202 241984 138258 242040
rect 150254 241984 150310 242040
rect 135994 234640 136050 234696
rect 135166 230152 135222 230208
rect 139214 233980 139270 234016
rect 139214 233960 139216 233980
rect 139216 233960 139268 233980
rect 139268 233960 139270 233980
rect 137282 223352 137338 223408
rect 140778 233008 140834 233064
rect 143446 231648 143502 231704
rect 142158 220496 142214 220552
rect 140686 207576 140742 207632
rect 146390 234232 146446 234288
rect 148138 241440 148194 241496
rect 148138 240488 148194 240544
rect 147678 237632 147734 237688
rect 150668 241440 150724 241496
rect 148138 238312 148194 238368
rect 145930 231512 145986 231568
rect 146206 231104 146262 231160
rect 146206 228792 146262 228848
rect 151082 228248 151138 228304
rect 139214 195880 139270 195936
rect 133786 193840 133842 193896
rect 152554 241848 152610 241904
rect 152462 237632 152518 237688
rect 151818 235592 151874 235648
rect 153014 234640 153070 234696
rect 153106 216280 153162 216336
rect 152462 214784 152518 214840
rect 154394 214784 154450 214840
rect 152462 206760 152518 206816
rect 155590 245792 155646 245848
rect 155498 241712 155554 241768
rect 155866 231376 155922 231432
rect 157246 326848 157302 326904
rect 156418 326440 156474 326496
rect 156142 310392 156198 310448
rect 157154 325372 157210 325408
rect 157154 325352 157156 325372
rect 157156 325352 157208 325372
rect 157208 325352 157210 325372
rect 156878 324264 156934 324320
rect 157246 322088 157302 322144
rect 157246 318844 157302 318880
rect 157246 318824 157248 318844
rect 157248 318824 157300 318844
rect 157300 318824 157302 318844
rect 156602 318688 156658 318744
rect 156602 317464 156658 317520
rect 156418 312568 156474 312624
rect 156234 308488 156290 308544
rect 157246 316920 157302 316976
rect 156786 315832 156842 315888
rect 157246 314744 157302 314800
rect 157246 311480 157302 311536
rect 157246 309576 157302 309632
rect 156694 308508 156750 308544
rect 156694 308488 156696 308508
rect 156696 308488 156748 308508
rect 156748 308488 156750 308508
rect 157246 306332 157302 306368
rect 157246 306312 157248 306332
rect 157248 306312 157300 306332
rect 157300 306312 157302 306332
rect 157246 305224 157302 305280
rect 157246 304136 157302 304192
rect 157246 303048 157302 303104
rect 157246 300056 157302 300112
rect 157246 298968 157302 299024
rect 156786 297880 156842 297936
rect 156602 296792 156658 296848
rect 157246 295704 157302 295760
rect 156418 294616 156474 294672
rect 157246 292712 157302 292768
rect 157246 291624 157302 291680
rect 157246 290536 157302 290592
rect 157246 289448 157302 289504
rect 156142 286184 156198 286240
rect 157246 285096 157302 285152
rect 156786 284280 156842 284336
rect 157154 283192 157210 283248
rect 157246 282104 157302 282160
rect 157246 281016 157302 281072
rect 157062 279928 157118 279984
rect 156970 278840 157026 278896
rect 156510 277752 156566 277808
rect 157246 275848 157302 275904
rect 157246 274760 157302 274816
rect 157246 273672 157302 273728
rect 157246 272584 157302 272640
rect 157246 271496 157302 271552
rect 156786 270408 156842 270464
rect 157246 269320 157302 269376
rect 156510 268232 156566 268288
rect 157246 267416 157302 267472
rect 157246 265240 157302 265296
rect 157246 263064 157302 263120
rect 156786 260888 156842 260944
rect 156694 259800 156750 259856
rect 156602 258984 156658 259040
rect 156050 254632 156106 254688
rect 156142 252456 156198 252512
rect 156602 245112 156658 245168
rect 156142 242972 156144 242992
rect 156144 242972 156196 242992
rect 156196 242972 156198 242992
rect 156142 242936 156198 242972
rect 155866 222264 155922 222320
rect 155866 217776 155922 217832
rect 157246 257932 157248 257952
rect 157248 257932 157300 257952
rect 157300 257932 157302 257952
rect 157246 257896 157302 257932
rect 157246 256808 157302 256864
rect 157246 255720 157302 255776
rect 157246 254632 157302 254688
rect 157246 253544 157302 253600
rect 156786 253136 156842 253192
rect 157246 251368 157302 251424
rect 157246 250552 157302 250608
rect 157154 249464 157210 249520
rect 157246 248376 157302 248432
rect 157246 247288 157302 247344
rect 157246 246200 157302 246256
rect 157246 244024 157302 244080
rect 156786 242120 156842 242176
rect 157430 329024 157486 329080
rect 157430 323176 157486 323232
rect 158074 337048 158130 337104
rect 158810 363568 158866 363624
rect 158810 319368 158866 319424
rect 159454 308352 159510 308408
rect 159362 297336 159418 297392
rect 159362 284280 159418 284336
rect 157338 235728 157394 235784
rect 156694 222808 156750 222864
rect 159454 243480 159510 243536
rect 158166 231512 158222 231568
rect 159730 243072 159786 243128
rect 159638 226072 159694 226128
rect 160190 357992 160246 358048
rect 160834 315288 160890 315344
rect 160926 303728 160982 303784
rect 160742 294480 160798 294536
rect 160098 237088 160154 237144
rect 159730 219136 159786 219192
rect 151726 190984 151782 191040
rect 160834 283464 160890 283520
rect 160926 275304 160982 275360
rect 162122 269048 162178 269104
rect 160834 234368 160890 234424
rect 162766 295996 162822 296032
rect 162766 295976 162768 295996
rect 162768 295976 162820 295996
rect 162820 295976 162822 295996
rect 162306 234232 162362 234288
rect 162398 228792 162454 228848
rect 164238 355408 164294 355464
rect 163778 332832 163834 332888
rect 163594 298152 163650 298208
rect 164974 289040 165030 289096
rect 164238 286320 164294 286376
rect 164238 269048 164294 269104
rect 163594 231648 163650 231704
rect 163502 227296 163558 227352
rect 165526 247016 165582 247072
rect 164974 241984 165030 242040
rect 166262 211792 166318 211848
rect 162122 200640 162178 200696
rect 172518 449948 172574 449984
rect 172518 449928 172520 449948
rect 172520 449928 172572 449948
rect 172572 449928 172574 449948
rect 168470 447344 168526 447400
rect 167826 325216 167882 325272
rect 167734 278024 167790 278080
rect 167642 237360 167698 237416
rect 166998 231784 167054 231840
rect 167642 230152 167698 230208
rect 167642 226072 167698 226128
rect 166538 225936 166594 225992
rect 167826 200912 167882 200968
rect 160742 187040 160798 187096
rect 107474 180920 107530 180976
rect 112258 179560 112314 179616
rect 106186 177520 106242 177576
rect 107474 177520 107530 177576
rect 116950 180784 117006 180840
rect 113730 177520 113786 177576
rect 112258 177112 112314 177168
rect 116950 177520 117006 177576
rect 119986 177520 120042 177576
rect 121366 177520 121422 177576
rect 118514 177112 118570 177168
rect 126058 177520 126114 177576
rect 129646 177520 129702 177576
rect 148966 177520 149022 177576
rect 99470 176704 99526 176760
rect 102046 176704 102102 176760
rect 103334 176704 103390 176760
rect 115846 176704 115902 176760
rect 124494 176704 124550 176760
rect 127622 176704 127678 176760
rect 132406 176704 132462 176760
rect 134430 176740 134432 176760
rect 134432 176740 134484 176760
rect 134484 176740 134486 176760
rect 134430 176704 134486 176740
rect 136086 176724 136142 176760
rect 158994 176740 158996 176760
rect 158996 176740 159048 176760
rect 159048 176740 159050 176760
rect 136086 176704 136088 176724
rect 136088 176704 136140 176724
rect 136140 176704 136142 176724
rect 130750 175752 130806 175808
rect 158994 176704 159050 176740
rect 123114 174936 123170 174992
rect 166354 176840 166410 176896
rect 166262 169632 166318 169688
rect 167734 180920 167790 180976
rect 67362 129240 67418 129296
rect 66166 126248 66222 126304
rect 66074 123528 66130 123584
rect 65982 120808 66038 120864
rect 67270 102312 67326 102368
rect 67270 95104 67326 95160
rect 67730 128016 67786 128072
rect 67454 125160 67510 125216
rect 67546 122576 67602 122632
rect 67454 81368 67510 81424
rect 64418 68312 64474 68368
rect 67638 100680 67694 100736
rect 67546 66136 67602 66192
rect 124034 94696 124090 94752
rect 86866 92384 86922 92440
rect 75826 91160 75882 91216
rect 86774 91160 86830 91216
rect 70214 76608 70270 76664
rect 67638 63416 67694 63472
rect 66166 60016 66222 60072
rect 64786 51720 64842 51776
rect 88154 91160 88210 91216
rect 79966 71032 80022 71088
rect 78586 61376 78642 61432
rect 73066 58520 73122 58576
rect 89074 92384 89130 92440
rect 98734 91432 98790 91488
rect 95054 91296 95110 91352
rect 91006 91160 91062 91216
rect 91926 91160 91982 91216
rect 93214 91160 93270 91216
rect 91926 88168 91982 88224
rect 93214 85448 93270 85504
rect 95146 91160 95202 91216
rect 96526 91160 96582 91216
rect 97906 91160 97962 91216
rect 99194 91160 99250 91216
rect 99286 80688 99342 80744
rect 99194 80008 99250 80064
rect 88246 75112 88302 75168
rect 82082 3576 82138 3632
rect 86774 17176 86830 17232
rect 95146 72528 95202 72584
rect 119710 93472 119766 93528
rect 121734 93472 121790 93528
rect 110142 93200 110198 93256
rect 105542 91704 105598 91760
rect 101862 91432 101918 91488
rect 100666 91160 100722 91216
rect 102046 91296 102102 91352
rect 101954 91160 102010 91216
rect 101862 86808 101918 86864
rect 100666 74296 100722 74352
rect 100666 58656 100722 58712
rect 102598 91160 102654 91216
rect 103426 91160 103482 91216
rect 104254 91160 104310 91216
rect 104806 91160 104862 91216
rect 104254 85176 104310 85232
rect 109958 92384 110014 92440
rect 107474 91704 107530 91760
rect 106186 85312 106242 85368
rect 105542 81232 105598 81288
rect 108854 91296 108910 91352
rect 107014 74432 107070 74488
rect 108946 91160 109002 91216
rect 158718 93064 158774 93120
rect 111614 92384 111670 92440
rect 114466 92384 114522 92440
rect 136086 92420 136088 92440
rect 136088 92420 136140 92440
rect 136140 92420 136142 92440
rect 136086 92384 136142 92420
rect 151358 92404 151414 92440
rect 151358 92384 151360 92404
rect 151360 92384 151412 92404
rect 151412 92384 151414 92404
rect 110326 91160 110382 91216
rect 111154 91160 111210 91216
rect 110142 89528 110198 89584
rect 112074 91160 112130 91216
rect 112994 91160 113050 91216
rect 113454 91160 113510 91216
rect 114282 91160 114338 91216
rect 126886 92248 126942 92304
rect 126610 91840 126666 91896
rect 114926 91704 114982 91760
rect 111154 88032 111210 88088
rect 112074 86672 112130 86728
rect 111062 82728 111118 82784
rect 117226 91568 117282 91624
rect 115754 91296 115810 91352
rect 118514 91296 118570 91352
rect 122838 91296 122894 91352
rect 125414 91296 125470 91352
rect 114926 89664 114982 89720
rect 115846 91160 115902 91216
rect 117226 91160 117282 91216
rect 115754 84088 115810 84144
rect 103426 57160 103482 57216
rect 111706 55800 111762 55856
rect 106922 54440 106978 54496
rect 108302 54440 108358 54496
rect 104162 28192 104218 28248
rect 105542 15816 105598 15872
rect 108302 3304 108358 3360
rect 116582 64232 116638 64288
rect 118606 91160 118662 91216
rect 119986 91160 120042 91216
rect 121366 91160 121422 91216
rect 122746 91160 122802 91216
rect 122102 82184 122158 82240
rect 124126 91160 124182 91216
rect 122746 83952 122802 84008
rect 125506 91160 125562 91216
rect 130750 91976 130806 92032
rect 126886 91568 126942 91624
rect 126702 91296 126758 91352
rect 126610 86536 126666 86592
rect 126794 91160 126850 91216
rect 127990 91160 128046 91216
rect 129646 91160 129702 91216
rect 151634 91296 151690 91352
rect 133786 91160 133842 91216
rect 134430 91160 134486 91216
rect 130750 90344 130806 90400
rect 151082 90344 151138 90400
rect 134430 87896 134486 87952
rect 151726 91160 151782 91216
rect 153106 91160 153162 91216
rect 151082 76744 151138 76800
rect 147034 66952 147090 67008
rect 126242 3576 126298 3632
rect 132958 10240 133014 10296
rect 121090 3440 121146 3496
rect 125874 3304 125930 3360
rect 163502 90344 163558 90400
rect 162214 88984 162270 89040
rect 151082 55936 151138 55992
rect 151082 40568 151138 40624
rect 165526 95104 165582 95160
rect 164974 92112 165030 92168
rect 166354 88168 166410 88224
rect 164882 86672 164938 86728
rect 167734 108976 167790 109032
rect 168286 111732 168288 111752
rect 168288 111732 168340 111752
rect 168340 111732 168342 111752
rect 168286 111696 168342 111732
rect 168010 111016 168066 111072
rect 167918 110372 167920 110392
rect 167920 110372 167972 110392
rect 167972 110372 167974 110392
rect 167918 110336 167974 110372
rect 167918 87896 167974 87952
rect 167826 85176 167882 85232
rect 164974 74296 165030 74352
rect 168470 237360 168526 237416
rect 169114 331472 169170 331528
rect 170402 298288 170458 298344
rect 170494 253136 170550 253192
rect 170954 247016 171010 247072
rect 170402 241440 170458 241496
rect 170954 233824 171010 233880
rect 170402 213288 170458 213344
rect 168470 174800 168526 174856
rect 169022 171264 169078 171320
rect 175922 343848 175978 343904
rect 171782 340992 171838 341048
rect 171138 247016 171194 247072
rect 172426 267824 172482 267880
rect 174634 339768 174690 339824
rect 174542 335960 174598 336016
rect 174542 300056 174598 300112
rect 173162 255448 173218 255504
rect 172518 241712 172574 241768
rect 172426 230288 172482 230344
rect 172426 228384 172482 228440
rect 173254 235728 173310 235784
rect 173714 227704 173770 227760
rect 171966 209480 172022 209536
rect 173162 187040 173218 187096
rect 171874 178200 171930 178256
rect 170494 117272 170550 117328
rect 169022 101360 169078 101416
rect 168654 93064 168710 93120
rect 169114 86808 169170 86864
rect 169022 81368 169078 81424
rect 170494 89528 170550 89584
rect 171782 88032 171838 88088
rect 172058 93608 172114 93664
rect 171966 74432 172022 74488
rect 136454 4800 136510 4856
rect 173714 223488 173770 223544
rect 173346 173848 173402 173904
rect 173254 86536 173310 86592
rect 177302 329976 177358 330032
rect 176014 319368 176070 319424
rect 176014 297472 176070 297528
rect 176014 284552 176070 284608
rect 176014 182144 176070 182200
rect 175922 160656 175978 160712
rect 175922 94016 175978 94072
rect 174726 85312 174782 85368
rect 178682 353504 178738 353560
rect 178682 293936 178738 293992
rect 178038 289040 178094 289096
rect 177394 236544 177450 236600
rect 177394 207712 177450 207768
rect 178958 236952 179014 237008
rect 202142 445984 202198 446040
rect 185582 371320 185638 371376
rect 181442 352008 181498 352064
rect 180062 346568 180118 346624
rect 180062 305632 180118 305688
rect 179418 235592 179474 235648
rect 178038 215328 178094 215384
rect 178682 214784 178738 214840
rect 177486 183776 177542 183832
rect 177394 111016 177450 111072
rect 177578 111016 177634 111072
rect 177394 108296 177450 108352
rect 177486 81232 177542 81288
rect 182822 338408 182878 338464
rect 182822 330384 182878 330440
rect 182822 315288 182878 315344
rect 183006 315288 183062 315344
rect 181626 291216 181682 291272
rect 181534 249056 181590 249112
rect 181534 217232 181590 217288
rect 181442 207712 181498 207768
rect 181442 175344 181498 175400
rect 182914 280880 182970 280936
rect 182822 231648 182878 231704
rect 182914 219272 182970 219328
rect 182086 187040 182142 187096
rect 180338 90344 180394 90400
rect 181534 82728 181590 82784
rect 182914 179560 182970 179616
rect 180062 12960 180118 13016
rect 177302 6160 177358 6216
rect 185582 281560 185638 281616
rect 184294 213968 184350 214024
rect 184294 198056 184350 198112
rect 185674 224168 185730 224224
rect 184386 97144 184442 97200
rect 184294 89664 184350 89720
rect 187054 347928 187110 347984
rect 187054 295432 187110 295488
rect 186962 247560 187018 247616
rect 187146 275984 187202 276040
rect 188342 271904 188398 271960
rect 188342 266328 188398 266384
rect 187146 234368 187202 234424
rect 187054 214648 187110 214704
rect 187238 214648 187294 214704
rect 186962 188400 187018 188456
rect 185766 175480 185822 175536
rect 195334 369824 195390 369880
rect 189814 305632 189870 305688
rect 189078 242936 189134 242992
rect 188986 228248 189042 228304
rect 188526 220632 188582 220688
rect 188434 196696 188490 196752
rect 189722 192480 189778 192536
rect 188434 183640 188490 183696
rect 188434 142160 188490 142216
rect 188526 80008 188582 80064
rect 193034 299784 193090 299840
rect 192574 287544 192630 287600
rect 189814 184320 189870 184376
rect 195242 345208 195298 345264
rect 195242 316648 195298 316704
rect 195242 313248 195298 313304
rect 193034 276936 193090 276992
rect 192942 248376 192998 248432
rect 192482 243072 192538 243128
rect 191838 219272 191894 219328
rect 192482 216688 192538 216744
rect 193034 213152 193090 213208
rect 193954 241440 194010 241496
rect 193862 221992 193918 222048
rect 194046 213152 194102 213208
rect 194506 241440 194562 241496
rect 194506 240488 194562 240544
rect 195058 225528 195114 225584
rect 194690 221720 194746 221776
rect 194690 213832 194746 213888
rect 193034 183096 193090 183152
rect 191746 179968 191802 180024
rect 191194 177248 191250 177304
rect 193862 202136 193918 202192
rect 193126 176568 193182 176624
rect 173162 3984 173218 4040
rect 191286 85448 191342 85504
rect 193862 43424 193918 43480
rect 195334 283736 195390 283792
rect 195978 278024 196034 278080
rect 195334 241576 195390 241632
rect 195334 230288 195390 230344
rect 196714 314744 196770 314800
rect 197266 314744 197322 314800
rect 197174 308352 197230 308408
rect 198002 292440 198058 292496
rect 198002 290128 198058 290184
rect 197358 282376 197414 282432
rect 197358 280744 197414 280800
rect 197450 280200 197506 280256
rect 197358 279384 197414 279440
rect 197358 278568 197414 278624
rect 197174 249056 197230 249112
rect 196714 247288 196770 247344
rect 196714 243752 196770 243808
rect 195886 229880 195942 229936
rect 197082 231512 197138 231568
rect 197082 230560 197138 230616
rect 197082 228384 197138 228440
rect 196714 223352 196770 223408
rect 195794 219272 195850 219328
rect 195334 215328 195390 215384
rect 195334 203496 195390 203552
rect 195334 202272 195390 202328
rect 197358 276664 197414 276720
rect 198278 288496 198334 288552
rect 198186 282920 198242 282976
rect 198094 278024 198150 278080
rect 198738 285776 198794 285832
rect 197450 275032 197506 275088
rect 197358 274488 197414 274544
rect 197358 273672 197414 273728
rect 197358 272856 197414 272912
rect 197358 271496 197414 271552
rect 197450 270952 197506 271008
rect 197358 270136 197414 270192
rect 197358 268776 197414 268832
rect 197358 266600 197414 266656
rect 197358 265784 197414 265840
rect 197358 264424 197414 264480
rect 197358 263628 197414 263664
rect 197358 263608 197360 263628
rect 197360 263608 197412 263628
rect 197412 263608 197414 263628
rect 197358 262284 197360 262304
rect 197360 262284 197412 262304
rect 197412 262284 197414 262304
rect 197358 262248 197414 262284
rect 197450 261432 197506 261488
rect 197358 260924 197360 260944
rect 197360 260924 197412 260944
rect 197412 260924 197414 260944
rect 197358 260888 197414 260924
rect 197358 260072 197414 260128
rect 197358 259256 197414 259312
rect 197450 258712 197506 258768
rect 197358 257896 197414 257952
rect 197358 256536 197414 256592
rect 198002 255176 198058 255232
rect 197358 254360 197414 254416
rect 197450 253544 197506 253600
rect 197450 252184 197506 252240
rect 197358 251640 197414 251696
rect 197450 250824 197506 250880
rect 197358 250008 197414 250064
rect 197450 249464 197506 249520
rect 197358 247832 197414 247888
rect 197358 246472 197414 246528
rect 197450 245928 197506 245984
rect 197450 245112 197506 245168
rect 197358 244316 197414 244352
rect 197358 244296 197360 244316
rect 197360 244296 197412 244316
rect 197412 244296 197414 244316
rect 197910 242120 197966 242176
rect 198002 241440 198058 241496
rect 199474 302096 199530 302152
rect 200946 302096 201002 302152
rect 200946 301008 201002 301064
rect 201314 301008 201370 301064
rect 200394 292440 200450 292496
rect 201130 292440 201186 292496
rect 201130 291760 201186 291816
rect 200578 290400 200634 290456
rect 582654 471416 582710 471472
rect 582470 458088 582526 458144
rect 582378 431568 582434 431624
rect 221462 367104 221518 367160
rect 206282 353640 206338 353696
rect 204902 352552 204958 352608
rect 202142 327120 202198 327176
rect 201682 303592 201738 303648
rect 204258 342352 204314 342408
rect 203522 292712 203578 292768
rect 202142 289856 202198 289912
rect 204166 292712 204222 292768
rect 210422 348336 210478 348392
rect 209042 334192 209098 334248
rect 207754 331200 207810 331256
rect 206374 309032 206430 309088
rect 206926 309032 206982 309088
rect 206926 307808 206982 307864
rect 206282 302232 206338 302288
rect 206650 302232 206706 302288
rect 204258 285640 204314 285696
rect 205178 285640 205234 285696
rect 204258 284552 204314 284608
rect 201958 284008 202014 284064
rect 206098 284280 206154 284336
rect 209134 332560 209190 332616
rect 209962 309304 210018 309360
rect 209042 309168 209098 309224
rect 209410 309168 209466 309224
rect 211158 331336 211214 331392
rect 210514 309304 210570 309360
rect 210422 304952 210478 305008
rect 210882 289992 210938 290048
rect 205362 283872 205418 283928
rect 211802 329160 211858 329216
rect 211986 293936 212042 293992
rect 211986 292848 212042 292904
rect 211802 284824 211858 284880
rect 212354 284824 212410 284880
rect 215942 363024 215998 363080
rect 213458 289040 213514 289096
rect 215390 336776 215446 336832
rect 214746 304952 214802 305008
rect 220082 338272 220138 338328
rect 215942 313928 215998 313984
rect 218702 336912 218758 336968
rect 216678 293936 216734 293992
rect 217690 293936 217746 293992
rect 216678 284824 216734 284880
rect 218610 292576 218666 292632
rect 218242 286320 218298 286376
rect 218702 285776 218758 285832
rect 220082 284280 220138 284336
rect 220726 285640 220782 285696
rect 221554 334328 221610 334384
rect 221554 310528 221610 310584
rect 221462 285776 221518 285832
rect 222934 296792 222990 296848
rect 222842 291896 222898 291952
rect 222106 285640 222162 285696
rect 223946 285640 224002 285696
rect 226430 342488 226486 342544
rect 225418 327392 225474 327448
rect 224222 284280 224278 284336
rect 225602 299648 225658 299704
rect 225970 297472 226026 297528
rect 216034 284008 216090 284064
rect 211618 283872 211674 283928
rect 214470 283872 214526 283928
rect 215942 283872 215998 283928
rect 226982 332696 227038 332752
rect 227810 299648 227866 299704
rect 226982 284280 227038 284336
rect 228454 335416 228510 335472
rect 230386 330384 230442 330440
rect 230018 310664 230074 310720
rect 228362 298424 228418 298480
rect 229006 298424 229062 298480
rect 231122 290128 231178 290184
rect 230478 284416 230534 284472
rect 231306 287136 231362 287192
rect 233882 357448 233938 357504
rect 232594 323584 232650 323640
rect 232502 285776 232558 285832
rect 231674 284416 231730 284472
rect 232778 284688 232834 284744
rect 234618 353368 234674 353424
rect 233974 328616 234030 328672
rect 226798 283872 226854 283928
rect 238206 327256 238262 327312
rect 238022 312432 238078 312488
rect 236826 299784 236882 299840
rect 236642 299512 236698 299568
rect 236458 287272 236514 287328
rect 239402 302368 239458 302424
rect 236826 293120 236882 293176
rect 238574 290128 238630 290184
rect 238114 287544 238170 287600
rect 238114 284552 238170 284608
rect 239586 302368 239642 302424
rect 239494 288360 239550 288416
rect 239954 291216 240010 291272
rect 240046 284280 240102 284336
rect 327078 368464 327134 368520
rect 240782 313928 240838 313984
rect 241426 295432 241482 295488
rect 243082 326304 243138 326360
rect 242346 285912 242402 285968
rect 243818 288360 243874 288416
rect 243174 284144 243230 284200
rect 243634 284008 243690 284064
rect 236274 283872 236330 283928
rect 244278 283192 244334 283248
rect 199474 263064 199530 263120
rect 199658 257352 199714 257408
rect 199934 257352 199990 257408
rect 200026 253000 200082 253056
rect 244462 268776 244518 268832
rect 245382 283192 245438 283248
rect 245658 282376 245714 282432
rect 245658 281016 245714 281072
rect 244646 278840 244702 278896
rect 244554 260888 244610 260944
rect 244462 255992 244518 256048
rect 200026 248512 200082 248568
rect 199474 245792 199530 245848
rect 198002 216688 198058 216744
rect 197266 197920 197322 197976
rect 197174 188400 197230 188456
rect 199842 244568 199898 244624
rect 199934 240352 199990 240408
rect 199842 240080 199898 240136
rect 244370 250280 244426 250336
rect 244370 247288 244426 247344
rect 244002 241304 244058 241360
rect 200118 240216 200174 240272
rect 200210 238584 200266 238640
rect 200578 240080 200634 240136
rect 200302 237904 200358 237960
rect 200578 237360 200634 237416
rect 200118 228928 200174 228984
rect 200210 227704 200266 227760
rect 200854 227704 200910 227760
rect 200762 215872 200818 215928
rect 199474 202136 199530 202192
rect 200854 210296 200910 210352
rect 201406 237360 201462 237416
rect 202050 238584 202106 238640
rect 202234 238448 202290 238504
rect 202234 213288 202290 213344
rect 204442 237224 204498 237280
rect 203522 233824 203578 233880
rect 204994 226072 205050 226128
rect 205086 224168 205142 224224
rect 203522 219272 203578 219328
rect 204902 215328 204958 215384
rect 203154 212336 203210 212392
rect 202970 205536 203026 205592
rect 203614 205536 203670 205592
rect 202234 186904 202290 186960
rect 198094 172352 198150 172408
rect 195242 13096 195298 13152
rect 191102 3440 191158 3496
rect 196806 84768 196862 84824
rect 198094 91704 198150 91760
rect 199474 95784 199530 95840
rect 202326 112376 202382 112432
rect 202234 73752 202290 73808
rect 205638 222128 205694 222184
rect 205638 221584 205694 221640
rect 205362 216552 205418 216608
rect 205362 215328 205418 215384
rect 205086 213152 205142 213208
rect 206466 221584 206522 221640
rect 206374 220768 206430 220824
rect 207386 216688 207442 216744
rect 209042 237360 209098 237416
rect 208858 234368 208914 234424
rect 207754 216688 207810 216744
rect 209686 233824 209742 233880
rect 209226 232872 209282 232928
rect 208398 206760 208454 206816
rect 210330 235592 210386 235648
rect 209870 221720 209926 221776
rect 211250 237360 211306 237416
rect 211802 232872 211858 232928
rect 212630 232872 212686 232928
rect 210422 209480 210478 209536
rect 209042 186904 209098 186960
rect 206926 184184 206982 184240
rect 206282 182960 206338 183016
rect 204902 178608 204958 178664
rect 203522 104216 203578 104272
rect 203614 84088 203670 84144
rect 206282 132504 206338 132560
rect 206374 115912 206430 115968
rect 206282 92248 206338 92304
rect 209226 120672 209282 120728
rect 209134 104080 209190 104136
rect 211802 199960 211858 200016
rect 213642 238584 213698 238640
rect 213090 237360 213146 237416
rect 213734 202952 213790 203008
rect 214562 237224 214618 237280
rect 214654 207032 214710 207088
rect 216034 234504 216090 234560
rect 216678 233960 216734 234016
rect 217322 222264 217378 222320
rect 217230 217912 217286 217968
rect 217230 217232 217286 217288
rect 218058 238040 218114 238096
rect 217506 210976 217562 211032
rect 215942 204040 215998 204096
rect 214654 195336 214710 195392
rect 213826 193976 213882 194032
rect 216034 177928 216090 177984
rect 218702 227568 218758 227624
rect 218978 213968 219034 214024
rect 220818 239400 220874 239456
rect 222106 233844 222162 233880
rect 222106 233824 222108 233844
rect 222108 233824 222160 233844
rect 222160 233824 222162 233844
rect 223394 238584 223450 238640
rect 221462 217776 221518 217832
rect 224314 239808 224370 239864
rect 224314 239400 224370 239456
rect 224774 237904 224830 237960
rect 223394 232464 223450 232520
rect 224222 231648 224278 231704
rect 223026 210432 223082 210488
rect 222934 199416 222990 199472
rect 220082 198600 220138 198656
rect 218702 192480 218758 192536
rect 218426 190440 218482 190496
rect 220082 178064 220138 178120
rect 214562 73888 214618 73944
rect 218702 104216 218758 104272
rect 222842 141344 222898 141400
rect 225234 240080 225290 240136
rect 224866 231648 224922 231704
rect 224866 218048 224922 218104
rect 225786 218048 225842 218104
rect 224774 119312 224830 119368
rect 226982 215872 227038 215928
rect 228178 240080 228234 240136
rect 228730 239944 228786 240000
rect 227626 238584 227682 238640
rect 230570 238176 230626 238232
rect 230202 233960 230258 234016
rect 227258 210840 227314 210896
rect 226154 205400 226210 205456
rect 231950 240116 231952 240136
rect 231952 240116 232004 240136
rect 232004 240116 232006 240136
rect 231950 240080 232006 240116
rect 231490 233144 231546 233200
rect 232502 239536 232558 239592
rect 229742 206896 229798 206952
rect 228362 189896 228418 189952
rect 227718 183096 227774 183152
rect 226982 182824 227038 182880
rect 224222 74024 224278 74080
rect 226982 90344 227038 90400
rect 220082 11600 220138 11656
rect 218702 4800 218758 4856
rect 229742 93880 229798 93936
rect 229834 93064 229890 93120
rect 228454 24112 228510 24168
rect 231306 135496 231362 135552
rect 231214 88984 231270 89040
rect 232686 239944 232742 240000
rect 232594 238448 232650 238504
rect 232594 229880 232650 229936
rect 232962 231784 233018 231840
rect 232594 204992 232650 205048
rect 234066 233008 234122 233064
rect 233882 229880 233938 229936
rect 233514 202816 233570 202872
rect 232594 180104 232650 180160
rect 232594 87488 232650 87544
rect 236458 238584 236514 238640
rect 235354 238448 235410 238504
rect 234986 224848 235042 224904
rect 237930 240080 237986 240136
rect 237930 237360 237986 237416
rect 238022 221584 238078 221640
rect 235998 215328 236054 215384
rect 236734 215328 236790 215384
rect 234066 133048 234122 133104
rect 234066 98640 234122 98696
rect 239218 239944 239274 240000
rect 238666 237360 238722 237416
rect 240690 237088 240746 237144
rect 239770 226208 239826 226264
rect 238298 216280 238354 216336
rect 241794 238584 241850 238640
rect 242254 239400 242310 239456
rect 242162 238312 242218 238368
rect 240782 192616 240838 192672
rect 238114 180784 238170 180840
rect 238022 176976 238078 177032
rect 237378 176704 237434 176760
rect 238114 165960 238170 166016
rect 240138 160656 240194 160712
rect 236642 88984 236698 89040
rect 236642 87624 236698 87680
rect 235998 61512 236054 61568
rect 238206 91024 238262 91080
rect 238114 86128 238170 86184
rect 236642 32408 236698 32464
rect 238114 28192 238170 28248
rect 232502 3304 232558 3360
rect 242346 235184 242402 235240
rect 242346 225528 242402 225584
rect 244094 234504 244150 234560
rect 244002 209616 244058 209672
rect 244370 227296 244426 227352
rect 245934 294480 245990 294536
rect 246118 281560 246174 281616
rect 246118 280200 246174 280256
rect 246118 279384 246174 279440
rect 246118 277480 246174 277536
rect 246026 276684 246082 276720
rect 246026 276664 246028 276684
rect 246028 276664 246080 276684
rect 246080 276664 246082 276684
rect 245934 275848 245990 275904
rect 245934 274488 245990 274544
rect 245842 273672 245898 273728
rect 245934 273128 245990 273184
rect 245842 272312 245898 272368
rect 245750 271496 245806 271552
rect 245658 270952 245714 271008
rect 245658 270136 245714 270192
rect 246302 270952 246358 271008
rect 245934 269592 245990 269648
rect 245934 267960 245990 268016
rect 246026 267416 246082 267472
rect 245934 266600 245990 266656
rect 245842 265784 245898 265840
rect 245750 265240 245806 265296
rect 245842 264424 245898 264480
rect 245934 263880 245990 263936
rect 245750 263064 245806 263120
rect 244922 260908 244978 260944
rect 244922 260888 244924 260908
rect 244924 260888 244976 260908
rect 244976 260888 244978 260908
rect 245934 262268 245990 262304
rect 245934 262248 245936 262268
rect 245936 262248 245988 262268
rect 245988 262248 245990 262268
rect 245842 261704 245898 261760
rect 245934 259528 245990 259584
rect 245934 258732 245990 258768
rect 245934 258712 245936 258732
rect 245936 258712 245988 258732
rect 245988 258712 245990 258732
rect 245842 258168 245898 258224
rect 245658 256536 245714 256592
rect 244922 248648 244978 248704
rect 244646 235728 244702 235784
rect 245750 251640 245806 251696
rect 245750 250824 245806 250880
rect 246026 255176 246082 255232
rect 245934 253852 245936 253872
rect 245936 253852 245988 253872
rect 245988 253852 245990 253872
rect 245934 253816 245990 253852
rect 245934 253000 245990 253056
rect 245934 249500 245936 249520
rect 245936 249500 245988 249520
rect 245988 249500 245990 249520
rect 245934 249464 245990 249500
rect 245934 248104 245990 248160
rect 245842 245112 245898 245168
rect 245750 240760 245806 240816
rect 245934 244568 245990 244624
rect 246026 239536 246082 239592
rect 246946 252184 247002 252240
rect 247130 278024 247186 278080
rect 247222 257372 247278 257408
rect 247222 257352 247224 257372
rect 247224 257352 247276 257372
rect 247276 257352 247278 257372
rect 248510 288496 248566 288552
rect 248418 254360 248474 254416
rect 246394 245928 246450 245984
rect 246302 244840 246358 244896
rect 246394 243752 246450 243808
rect 246302 242392 246358 242448
rect 245658 228928 245714 228984
rect 245658 227704 245714 227760
rect 245934 235864 245990 235920
rect 246302 227704 246358 227760
rect 244462 219272 244518 219328
rect 241518 189760 241574 189816
rect 240874 133864 240930 133920
rect 240874 111016 240930 111072
rect 240230 6976 240286 7032
rect 240230 3984 240286 4040
rect 244278 184320 244334 184376
rect 243542 142704 243598 142760
rect 242898 6160 242954 6216
rect 243634 82320 243690 82376
rect 243634 40568 243690 40624
rect 245658 200776 245714 200832
rect 244922 176432 244978 176488
rect 245014 91432 245070 91488
rect 245014 80824 245070 80880
rect 249890 317464 249946 317520
rect 249982 298152 250038 298208
rect 249706 235184 249762 235240
rect 262218 364384 262274 364440
rect 252558 356088 252614 356144
rect 251362 347792 251418 347848
rect 251454 295568 251510 295624
rect 248326 210568 248382 210624
rect 247682 207712 247738 207768
rect 246394 119312 246450 119368
rect 246302 94968 246358 95024
rect 243542 3304 243598 3360
rect 250442 204856 250498 204912
rect 249062 179424 249118 179480
rect 248602 172896 248658 172952
rect 248602 171536 248658 171592
rect 247774 169632 247830 169688
rect 248418 166948 248420 166968
rect 248420 166948 248472 166968
rect 248472 166948 248474 166968
rect 248418 166912 248474 166948
rect 248510 166368 248566 166424
rect 248418 165008 248474 165064
rect 248418 163648 248474 163704
rect 248510 162968 248566 163024
rect 248418 162288 248474 162344
rect 248510 161744 248566 161800
rect 248418 161064 248474 161120
rect 248510 160384 248566 160440
rect 248418 159024 248474 159080
rect 248418 158344 248474 158400
rect 249706 176432 249762 176488
rect 249522 175616 249578 175672
rect 249706 174936 249762 174992
rect 249706 173576 249762 173632
rect 249338 172216 249394 172272
rect 249706 171012 249762 171048
rect 249706 170992 249708 171012
rect 249708 170992 249760 171012
rect 249760 170992 249762 171012
rect 249614 170312 249670 170368
rect 249706 169668 249708 169688
rect 249708 169668 249760 169688
rect 249760 169668 249762 169688
rect 249706 169632 249762 169668
rect 249246 168952 249302 169008
rect 249706 168292 249762 168328
rect 249706 168272 249708 168292
rect 249708 168272 249760 168292
rect 249760 168272 249762 168292
rect 249614 167592 249670 167648
rect 249154 159704 249210 159760
rect 249062 157664 249118 157720
rect 249154 154400 249210 154456
rect 248970 153040 249026 153096
rect 249338 152496 249394 152552
rect 249246 151136 249302 151192
rect 248970 149096 249026 149152
rect 249246 147872 249302 147928
rect 249154 147192 249210 147248
rect 249154 144472 249210 144528
rect 249154 140528 249210 140584
rect 248970 139848 249026 139904
rect 247774 132776 247830 132832
rect 249062 139168 249118 139224
rect 249154 137944 249210 138000
rect 249154 136584 249210 136640
rect 248970 124072 249026 124128
rect 248786 122032 248842 122088
rect 248786 119448 248842 119504
rect 248786 118088 248842 118144
rect 248786 116728 248842 116784
rect 247866 114960 247922 115016
rect 247774 112376 247830 112432
rect 248970 112104 249026 112160
rect 248970 110744 249026 110800
rect 248786 106120 248842 106176
rect 248510 103536 248566 103592
rect 248786 101496 248842 101552
rect 248510 101360 248566 101416
rect 249706 157120 249762 157176
rect 249614 156440 249670 156496
rect 249706 155760 249762 155816
rect 249614 155080 249670 155136
rect 249706 153720 249762 153776
rect 249706 151852 249708 151872
rect 249708 151852 249760 151872
rect 249760 151852 249762 151872
rect 249706 151816 249762 151852
rect 249706 150476 249762 150512
rect 249706 150456 249708 150476
rect 249708 150456 249760 150476
rect 249760 150456 249762 150476
rect 249614 149776 249670 149832
rect 249430 148416 249486 148472
rect 249706 146512 249762 146568
rect 249614 145832 249670 145888
rect 249706 145152 249762 145208
rect 249706 143792 249762 143848
rect 249706 142568 249762 142624
rect 249614 141888 249670 141944
rect 249706 141208 249762 141264
rect 249706 138624 249762 138680
rect 249706 137264 249762 137320
rect 249706 135904 249762 135960
rect 249706 134544 249762 134600
rect 249706 131960 249762 132016
rect 249246 131280 249302 131336
rect 249614 130600 249670 130656
rect 249706 129920 249762 129976
rect 249706 129240 249762 129296
rect 249614 128016 249670 128072
rect 249706 127336 249762 127392
rect 249614 126656 249670 126712
rect 249706 125976 249762 126032
rect 249614 125296 249670 125352
rect 249706 124616 249762 124672
rect 249522 123392 249578 123448
rect 249706 122712 249762 122768
rect 249614 121352 249670 121408
rect 249246 120672 249302 120728
rect 249706 120672 249762 120728
rect 249706 119992 249762 120048
rect 249614 118768 249670 118824
rect 249706 114824 249762 114880
rect 249614 114144 249670 114200
rect 249706 113464 249762 113520
rect 249246 112784 249302 112840
rect 249246 111424 249302 111480
rect 249614 110200 249670 110256
rect 249706 109520 249762 109576
rect 249706 108840 249762 108896
rect 249154 108296 249210 108352
rect 249522 108160 249578 108216
rect 249706 107480 249762 107536
rect 249522 106800 249578 106856
rect 249706 105576 249762 105632
rect 249614 104896 249670 104952
rect 249706 104216 249762 104272
rect 249614 104080 249670 104136
rect 249706 102856 249762 102912
rect 249246 102176 249302 102232
rect 249154 100952 249210 101008
rect 249706 100272 249762 100328
rect 249522 99592 249578 99648
rect 249062 89120 249118 89176
rect 248418 71168 248474 71224
rect 247682 6160 247738 6216
rect 249246 96872 249302 96928
rect 249154 66136 249210 66192
rect 249338 96328 249394 96384
rect 249614 98912 249670 98968
rect 249706 98232 249762 98288
rect 249706 97552 249762 97608
rect 249522 95784 249578 95840
rect 249798 75248 249854 75304
rect 249246 63416 249302 63472
rect 250534 178064 250590 178120
rect 251454 259800 251510 259856
rect 255318 355272 255374 355328
rect 252558 240080 252614 240136
rect 253938 290128 253994 290184
rect 252650 238312 252706 238368
rect 252650 237360 252706 237416
rect 253202 237360 253258 237416
rect 251822 232600 251878 232656
rect 251362 224712 251418 224768
rect 250718 190576 250774 190632
rect 250718 172352 250774 172408
rect 250626 128696 250682 128752
rect 250718 98640 250774 98696
rect 250626 93744 250682 93800
rect 254122 298288 254178 298344
rect 259458 350648 259514 350704
rect 258170 326848 258226 326904
rect 256790 312432 256846 312488
rect 255962 293936 256018 293992
rect 253938 220768 253994 220824
rect 254582 220768 254638 220824
rect 255318 212472 255374 212528
rect 258722 282104 258778 282160
rect 256054 212472 256110 212528
rect 256054 185816 256110 185872
rect 259458 238448 259514 238504
rect 259458 237904 259514 237960
rect 258722 222944 258778 223000
rect 260102 220088 260158 220144
rect 260102 217232 260158 217288
rect 258722 189760 258778 189816
rect 258814 184320 258870 184376
rect 258078 180784 258134 180840
rect 259366 178200 259422 178256
rect 259366 177928 259422 177984
rect 260102 177384 260158 177440
rect 259734 176568 259790 176624
rect 261574 287272 261630 287328
rect 317418 320728 317474 320784
rect 262218 264152 262274 264208
rect 262954 287680 263010 287736
rect 263966 287136 264022 287192
rect 261482 175888 261538 175944
rect 262218 175752 262274 175808
rect 251822 173848 251878 173904
rect 264150 177520 264206 177576
rect 264334 176840 264390 176896
rect 264886 177248 264942 177304
rect 264242 174664 264298 174720
rect 264150 174256 264206 174312
rect 264978 175208 265034 175264
rect 264426 171400 264482 171456
rect 264058 164464 264114 164520
rect 265162 175888 265218 175944
rect 265162 164736 265218 164792
rect 265070 160520 265126 160576
rect 265070 154400 265126 154456
rect 264886 153720 264942 153776
rect 264886 150456 264942 150512
rect 266450 232600 266506 232656
rect 266358 193160 266414 193216
rect 265622 176568 265678 176624
rect 266358 173748 266360 173768
rect 266360 173748 266412 173768
rect 266412 173748 266414 173768
rect 266358 173712 266414 173748
rect 266358 172388 266360 172408
rect 266360 172388 266412 172408
rect 266412 172388 266414 172408
rect 266358 172352 266414 172388
rect 266358 170448 266414 170504
rect 266358 169496 266414 169552
rect 266358 168988 266360 169008
rect 266360 168988 266412 169008
rect 266412 168988 266414 169008
rect 266358 168952 266414 168988
rect 266358 167592 266414 167648
rect 266358 166096 266414 166152
rect 265346 165552 265402 165608
rect 266358 165144 266414 165200
rect 266358 163376 266414 163432
rect 266358 161880 266414 161936
rect 266358 160928 266414 160984
rect 267002 220224 267058 220280
rect 266634 172760 266690 172816
rect 266634 171808 266690 171864
rect 266542 161472 266598 161528
rect 266542 160112 266598 160168
rect 266450 159976 266506 160032
rect 266358 158072 266414 158128
rect 266358 157120 266414 157176
rect 266726 169904 266782 169960
rect 267002 169088 267058 169144
rect 266726 167592 266782 167648
rect 266726 162832 266782 162888
rect 266818 159296 266874 159352
rect 266634 157664 266690 157720
rect 266542 156848 266598 156904
rect 266450 156712 266506 156768
rect 266358 155760 266414 155816
rect 266450 155216 266506 155272
rect 265346 152496 265402 152552
rect 265254 149096 265310 149152
rect 264150 146240 264206 146296
rect 264150 139712 264206 139768
rect 264334 145560 264390 145616
rect 265438 142024 265494 142080
rect 264334 141616 264390 141672
rect 265438 140800 265494 140856
rect 265438 137264 265494 137320
rect 265438 136720 265494 136776
rect 264150 127880 264206 127936
rect 264886 131416 264942 131472
rect 264058 105304 264114 105360
rect 264150 96600 264206 96656
rect 257894 95920 257950 95976
rect 261022 95920 261078 95976
rect 262862 95920 262918 95976
rect 257802 95784 257858 95840
rect 254582 90480 254638 90536
rect 255318 69672 255374 69728
rect 255410 63552 255466 63608
rect 255410 61512 255466 61568
rect 254674 6160 254730 6216
rect 253478 3440 253534 3496
rect 257342 64232 257398 64288
rect 256698 43424 256754 43480
rect 258814 91840 258870 91896
rect 262218 68312 262274 68368
rect 258814 39208 258870 39264
rect 258722 22616 258778 22672
rect 258262 3304 258318 3360
rect 263046 95784 263102 95840
rect 262954 94424 263010 94480
rect 262954 66952 263010 67008
rect 264334 97144 264390 97200
rect 266358 153856 266414 153912
rect 266358 153348 266360 153368
rect 266360 153348 266412 153368
rect 266412 153348 266414 153368
rect 266358 153312 266414 153348
rect 266726 152904 266782 152960
rect 266726 152360 266782 152416
rect 266174 148280 266230 148336
rect 265714 126384 265770 126440
rect 265714 123800 265770 123856
rect 265622 102312 265678 102368
rect 264886 99048 264942 99104
rect 261758 14456 261814 14512
rect 265898 120536 265954 120592
rect 265714 72528 265770 72584
rect 266358 151580 266360 151600
rect 266360 151580 266412 151600
rect 266412 151580 266414 151600
rect 266358 151544 266414 151580
rect 266450 151272 266506 151328
rect 266358 149640 266414 149696
rect 266818 151952 266874 152008
rect 266726 150048 266782 150104
rect 266542 149640 266598 149696
rect 266542 148688 266598 148744
rect 266450 148144 266506 148200
rect 266358 147192 266414 147248
rect 266358 143928 266414 143984
rect 267646 168000 267702 168056
rect 269118 213868 269120 213888
rect 269120 213868 269172 213888
rect 269172 213868 269174 213888
rect 269118 213832 269174 213868
rect 267922 182960 267978 183016
rect 267646 166640 267702 166696
rect 267738 160656 267794 160712
rect 267646 159568 267702 159624
rect 267002 143384 267058 143440
rect 266358 142976 266414 143032
rect 266358 138760 266414 138816
rect 266358 135904 266414 135960
rect 266358 135360 266414 135416
rect 266450 134952 266506 135008
rect 267002 134544 267058 134600
rect 266358 134408 266414 134464
rect 266358 133048 266414 133104
rect 266358 132504 266414 132560
rect 266358 131552 266414 131608
rect 266450 131144 266506 131200
rect 266358 131008 266414 131064
rect 266358 130192 266414 130248
rect 266450 129784 266506 129840
rect 266358 129240 266414 129296
rect 266542 128832 266598 128888
rect 266542 128152 266598 128208
rect 266358 127336 266414 127392
rect 266358 125976 266414 126032
rect 266358 125432 266414 125488
rect 266450 125024 266506 125080
rect 267094 134000 267150 134056
rect 267646 144880 267702 144936
rect 268014 176568 268070 176624
rect 268382 159024 268438 159080
rect 267738 144744 267794 144800
rect 267186 133456 267242 133512
rect 266542 124072 266598 124128
rect 266634 123392 266690 123448
rect 266358 123156 266360 123176
rect 266360 123156 266412 123176
rect 266412 123156 266414 123176
rect 266358 123120 266414 123156
rect 266358 122576 266414 122632
rect 266358 118904 266414 118960
rect 266358 118088 266414 118144
rect 266174 117952 266230 118008
rect 266174 114960 266230 115016
rect 266358 116456 266414 116512
rect 266358 116048 266414 116104
rect 266358 115504 266414 115560
rect 266266 114688 266322 114744
rect 266358 113636 266360 113656
rect 266360 113636 266412 113656
rect 266412 113636 266414 113656
rect 266358 113600 266414 113636
rect 266358 112648 266414 112704
rect 266542 122168 266598 122224
rect 266910 121624 266966 121680
rect 266634 120672 266690 120728
rect 266542 119312 266598 119368
rect 266542 117408 266598 117464
rect 266542 115096 266598 115152
rect 267094 120264 267150 120320
rect 276662 285776 276718 285832
rect 269762 173304 269818 173360
rect 270038 170312 270094 170368
rect 269210 158480 269266 158536
rect 269118 157392 269174 157448
rect 268382 118360 268438 118416
rect 267186 118088 267242 118144
rect 267094 116456 267150 116512
rect 267002 114552 267058 114608
rect 266542 113192 266598 113248
rect 266542 112240 266598 112296
rect 266542 111968 266598 112024
rect 266450 110744 266506 110800
rect 266450 109792 266506 109848
rect 266358 109384 266414 109440
rect 266358 108432 266414 108488
rect 266542 107888 266598 107944
rect 266358 107072 266414 107128
rect 266450 106528 266506 106584
rect 266358 105576 266414 105632
rect 266358 103672 266414 103728
rect 266358 103264 266414 103320
rect 266450 102720 266506 102776
rect 266450 102040 266506 102096
rect 266358 101768 266414 101824
rect 266634 101360 266690 101416
rect 266450 100816 266506 100872
rect 266358 100408 266414 100464
rect 266542 100000 266598 100056
rect 266450 99864 266506 99920
rect 266358 98640 266414 98696
rect 266634 99456 266690 99512
rect 266542 98504 266598 98560
rect 266450 97960 266506 98016
rect 266358 97552 266414 97608
rect 266910 97280 266966 97336
rect 266910 96600 266966 96656
rect 266450 96192 266506 96248
rect 268934 124752 268990 124808
rect 268658 122168 268714 122224
rect 268566 111832 268622 111888
rect 267186 111288 267242 111344
rect 267278 110200 267334 110256
rect 267094 101496 267150 101552
rect 268382 105168 268438 105224
rect 268290 102448 268346 102504
rect 267646 97008 267702 97064
rect 267738 93472 267794 93528
rect 266542 4800 266598 4856
rect 268934 110472 268990 110528
rect 268658 110200 268714 110256
rect 269026 102176 269082 102232
rect 268658 86128 268714 86184
rect 268382 13096 268438 13152
rect 270682 177384 270738 177440
rect 271970 197920 272026 197976
rect 271878 194112 271934 194168
rect 270682 165688 270738 165744
rect 270590 162696 270646 162752
rect 271142 155216 271198 155272
rect 269854 102176 269910 102232
rect 270222 109112 270278 109168
rect 270130 103808 270186 103864
rect 271970 165552 272026 165608
rect 272706 170040 272762 170096
rect 272154 168544 272210 168600
rect 272522 157528 272578 157584
rect 271970 144744 272026 144800
rect 271786 129920 271842 129976
rect 271418 115776 271474 115832
rect 271326 107616 271382 107672
rect 270222 102312 270278 102368
rect 271234 100952 271290 101008
rect 271418 100816 271474 100872
rect 273442 164192 273498 164248
rect 273442 155896 273498 155952
rect 272706 130600 272762 130656
rect 273994 164600 274050 164656
rect 276018 223524 276020 223544
rect 276020 223524 276072 223544
rect 276072 223524 276074 223544
rect 276018 223488 276074 223524
rect 274822 176840 274878 176896
rect 275282 162016 275338 162072
rect 274730 159296 274786 159352
rect 272614 126928 272670 126984
rect 272522 111016 272578 111072
rect 272062 100816 272118 100872
rect 271786 96464 271842 96520
rect 271510 90480 271566 90536
rect 274086 124616 274142 124672
rect 273258 117816 273314 117872
rect 273258 113736 273314 113792
rect 273994 109792 274050 109848
rect 273166 104760 273222 104816
rect 271326 3304 271382 3360
rect 274178 103944 274234 104000
rect 276202 170176 276258 170232
rect 275558 157936 275614 157992
rect 274546 121624 274602 121680
rect 274546 121488 274602 121544
rect 276846 166368 276902 166424
rect 276754 151136 276810 151192
rect 275650 131688 275706 131744
rect 277582 170312 277638 170368
rect 277490 166504 277546 166560
rect 278042 160384 278098 160440
rect 275650 121488 275706 121544
rect 276662 117408 276718 117464
rect 275558 110744 275614 110800
rect 275374 68176 275430 68232
rect 273902 30912 273958 30968
rect 274822 3304 274878 3360
rect 277306 125976 277362 126032
rect 278226 153856 278282 153912
rect 278134 152360 278190 152416
rect 278042 119992 278098 120048
rect 277306 117952 277362 118008
rect 277030 114960 277086 115016
rect 277030 113736 277086 113792
rect 276846 106256 276902 106312
rect 277030 98776 277086 98832
rect 276846 58520 276902 58576
rect 278870 187040 278926 187096
rect 278778 167320 278834 167376
rect 278778 157392 278834 157448
rect 279514 172760 279570 172816
rect 278870 156848 278926 156904
rect 278318 132368 278374 132424
rect 280802 301008 280858 301064
rect 280342 232464 280398 232520
rect 279422 115776 279478 115832
rect 278778 25472 278834 25528
rect 276110 19896 276166 19952
rect 278318 3984 278374 4040
rect 280066 147056 280122 147112
rect 279790 143792 279846 143848
rect 280066 143520 280122 143576
rect 281538 167592 281594 167648
rect 282182 168408 282238 168464
rect 279790 116456 279846 116512
rect 279698 84768 279754 84824
rect 279606 55800 279662 55856
rect 294602 314744 294658 314800
rect 283010 222264 283066 222320
rect 282918 166232 282974 166288
rect 282274 148688 282330 148744
rect 282182 128288 282238 128344
rect 282182 115912 282238 115968
rect 281446 113328 281502 113384
rect 280894 87488 280950 87544
rect 281446 106120 281502 106176
rect 281078 60016 281134 60072
rect 282274 103536 282330 103592
rect 282182 46144 282238 46200
rect 287702 302368 287758 302424
rect 283010 157936 283066 157992
rect 282550 142704 282606 142760
rect 282458 122168 282514 122224
rect 283562 117136 283618 117192
rect 282458 108976 282514 109032
rect 285218 174392 285274 174448
rect 284942 168544 284998 168600
rect 284298 160656 284354 160712
rect 285034 155896 285090 155952
rect 283838 138624 283894 138680
rect 283838 122032 283894 122088
rect 283654 110336 283710 110392
rect 282918 102448 282974 102504
rect 282458 98232 282514 98288
rect 282458 91840 282514 91896
rect 283930 113736 283986 113792
rect 284298 112648 284354 112704
rect 284298 109656 284354 109712
rect 284022 105440 284078 105496
rect 285770 184320 285826 184376
rect 285678 162696 285734 162752
rect 287702 238176 287758 238232
rect 287610 173576 287666 173632
rect 287242 172216 287298 172272
rect 286414 170040 286470 170096
rect 286322 162832 286378 162888
rect 285770 156712 285826 156768
rect 287426 164464 287482 164520
rect 287426 163376 287482 163432
rect 287150 161880 287206 161936
rect 286506 160248 286562 160304
rect 286414 131008 286470 131064
rect 286414 123256 286470 123312
rect 283930 98640 283986 98696
rect 284114 97960 284170 98016
rect 284298 94424 284354 94480
rect 284942 82048 284998 82104
rect 284298 66816 284354 66872
rect 283930 59880 283986 59936
rect 280802 10240 280858 10296
rect 280710 3304 280766 3360
rect 286322 108704 286378 108760
rect 285586 100952 285642 101008
rect 285126 71032 285182 71088
rect 285034 62736 285090 62792
rect 287518 161064 287574 161120
rect 287426 158888 287482 158944
rect 287978 175616 288034 175672
rect 287794 175208 287850 175264
rect 287886 174800 287942 174856
rect 288346 173984 288402 174040
rect 288346 172624 288402 172680
rect 288254 171808 288310 171864
rect 288346 171400 288402 171456
rect 288346 170992 288402 171048
rect 288162 169632 288218 169688
rect 288254 169224 288310 169280
rect 287978 167864 288034 167920
rect 288346 167068 288402 167104
rect 288346 167048 288348 167068
rect 288348 167048 288400 167068
rect 288400 167048 288402 167068
rect 288346 166640 288402 166696
rect 288254 166368 288310 166424
rect 288254 166232 288310 166288
rect 288070 165824 288126 165880
rect 287794 164872 287850 164928
rect 287886 163648 287942 163704
rect 287702 157392 287758 157448
rect 286598 154808 286654 154864
rect 287242 148552 287298 148608
rect 287794 154536 287850 154592
rect 287702 147056 287758 147112
rect 287426 146920 287482 146976
rect 287426 145696 287482 145752
rect 287426 145152 287482 145208
rect 287702 144336 287758 144392
rect 287426 141208 287482 141264
rect 287150 133592 287206 133648
rect 288162 164056 288218 164112
rect 288254 163240 288310 163296
rect 288070 162016 288126 162072
rect 288346 162288 288402 162344
rect 288346 159704 288402 159760
rect 288254 158480 288310 158536
rect 288162 157120 288218 157176
rect 288070 156712 288126 156768
rect 287978 155896 288034 155952
rect 288070 155216 288126 155272
rect 288346 158072 288402 158128
rect 290462 284416 290518 284472
rect 288438 156576 288494 156632
rect 288346 155080 288402 155136
rect 288254 152496 288310 152552
rect 288346 151952 288402 152008
rect 288346 151544 288402 151600
rect 287978 151136 288034 151192
rect 288254 150728 288310 150784
rect 288346 150320 288402 150376
rect 288254 149776 288310 149832
rect 288346 148960 288402 149016
rect 288530 148688 288586 148744
rect 288530 147872 288586 147928
rect 288346 147328 288402 147384
rect 288070 145968 288126 146024
rect 287978 142976 288034 143032
rect 287886 142568 287942 142624
rect 287794 139576 287850 139632
rect 287150 128288 287206 128344
rect 287150 124480 287206 124536
rect 286690 121624 286746 121680
rect 286598 114416 286654 114472
rect 286506 112104 286562 112160
rect 287702 123664 287758 123720
rect 287610 119312 287666 119368
rect 286966 118904 287022 118960
rect 286782 113192 286838 113248
rect 286690 111016 286746 111072
rect 287426 116320 287482 116376
rect 287610 113736 287666 113792
rect 286966 111968 287022 112024
rect 287610 101768 287666 101824
rect 286598 97552 286654 97608
rect 286414 80688 286470 80744
rect 288254 145560 288310 145616
rect 288162 144744 288218 144800
rect 291934 235184 291990 235240
rect 291842 189624 291898 189680
rect 301226 299648 301282 299704
rect 296074 214648 296130 214704
rect 297362 181464 297418 181520
rect 295982 179968 296038 180024
rect 297454 178064 297510 178120
rect 294602 177384 294658 177440
rect 291934 177248 291990 177304
rect 302882 291216 302938 291272
rect 300858 176704 300914 176760
rect 300858 176024 300914 176080
rect 298190 175888 298246 175944
rect 289174 167456 289230 167512
rect 288714 164600 288770 164656
rect 289082 153720 289138 153776
rect 288622 139984 288678 140040
rect 288254 139168 288310 139224
rect 288346 138216 288402 138272
rect 288346 137400 288402 137456
rect 288346 133048 288402 133104
rect 288346 132232 288402 132288
rect 288346 130464 288402 130520
rect 288070 129648 288126 129704
rect 287978 129240 288034 129296
rect 287978 127880 288034 127936
rect 288162 127472 288218 127528
rect 288070 124752 288126 124808
rect 287978 124072 288034 124128
rect 288254 126248 288310 126304
rect 288346 125840 288402 125896
rect 288346 125296 288402 125352
rect 288530 123800 288586 123856
rect 288530 122984 288586 123040
rect 288254 121508 288310 121544
rect 288254 121488 288256 121508
rect 288256 121488 288308 121508
rect 288308 121488 288310 121508
rect 288254 121080 288310 121136
rect 288254 117680 288310 117736
rect 288162 117136 288218 117192
rect 288070 115096 288126 115152
rect 287978 114144 288034 114200
rect 287886 113056 287942 113112
rect 287794 108976 287850 109032
rect 287978 111560 288034 111616
rect 287978 107344 288034 107400
rect 287978 105576 288034 105632
rect 288254 114572 288310 114608
rect 288254 114552 288256 114572
rect 288256 114552 288308 114572
rect 288308 114552 288310 114572
rect 301686 189760 301742 189816
rect 301686 176568 301742 176624
rect 301410 175208 301466 175264
rect 301410 174392 301466 174448
rect 301318 170584 301374 170640
rect 301318 160792 301374 160848
rect 301318 150592 301374 150648
rect 289358 138624 289414 138680
rect 289266 136176 289322 136232
rect 289174 131008 289230 131064
rect 288346 111968 288402 112024
rect 288254 111152 288310 111208
rect 288254 110336 288310 110392
rect 288346 109520 288402 109576
rect 288346 108568 288402 108624
rect 289082 108160 289138 108216
rect 288346 106936 288402 106992
rect 288346 105984 288402 106040
rect 288530 103944 288586 104000
rect 288530 103536 288586 103592
rect 288346 103400 288402 103456
rect 288254 102584 288310 102640
rect 287978 102448 288034 102504
rect 288346 101224 288402 101280
rect 288254 100408 288310 100464
rect 288346 99592 288402 99648
rect 288530 98776 288586 98832
rect 288530 98232 288586 98288
rect 287794 97960 287850 98016
rect 287702 82184 287758 82240
rect 287886 97416 287942 97472
rect 288346 97008 288402 97064
rect 287886 86128 287942 86184
rect 287794 77968 287850 78024
rect 286598 77832 286654 77888
rect 289450 136584 289506 136640
rect 289358 130328 289414 130384
rect 302882 188400 302938 188456
rect 302330 185680 302386 185736
rect 302514 178064 302570 178120
rect 302330 161744 302386 161800
rect 304354 213288 304410 213344
rect 304262 202272 304318 202328
rect 304262 182960 304318 183016
rect 303618 172488 303674 172544
rect 302514 168680 302570 168736
rect 302422 159432 302478 159488
rect 303618 157936 303674 157992
rect 303618 154944 303674 155000
rect 303618 154128 303674 154184
rect 304446 179968 304502 180024
rect 303894 171672 303950 171728
rect 304906 170856 304962 170912
rect 315946 310528 316002 310584
rect 315946 306584 316002 306640
rect 315946 306312 316002 306368
rect 315946 296792 316002 296848
rect 315946 296656 316002 296712
rect 313278 292848 313334 292904
rect 309138 289856 309194 289912
rect 307022 284008 307078 284064
rect 303894 169360 303950 169416
rect 303894 167048 303950 167104
rect 303894 166368 303950 166424
rect 303894 164872 303950 164928
rect 303894 164056 303950 164112
rect 303894 163276 303896 163296
rect 303896 163276 303948 163296
rect 303948 163276 303950 163296
rect 303894 163240 303950 163276
rect 303894 162560 303950 162616
rect 303894 161064 303950 161120
rect 303802 158752 303858 158808
rect 303802 157292 303804 157312
rect 303804 157292 303856 157312
rect 303856 157292 303858 157312
rect 303802 157256 303858 157292
rect 303894 156440 303950 156496
rect 303802 155624 303858 155680
rect 303802 153448 303858 153504
rect 303802 152632 303858 152688
rect 303894 151816 303950 151872
rect 303710 151136 303766 151192
rect 303802 149640 303858 149696
rect 303802 148824 303858 148880
rect 303710 147328 303766 147384
rect 303802 145832 303858 145888
rect 303710 145016 303766 145072
rect 303802 144200 303858 144256
rect 303986 142024 304042 142080
rect 303802 141208 303858 141264
rect 303618 139712 303674 139768
rect 304906 148008 304962 148064
rect 304262 138896 304318 138952
rect 303802 138216 303858 138272
rect 303802 137400 303858 137456
rect 303618 135904 303674 135960
rect 303710 134408 303766 134464
rect 303802 133592 303858 133648
rect 303894 132776 303950 132832
rect 303802 132096 303858 132152
rect 303894 131280 303950 131336
rect 303802 130600 303858 130656
rect 303802 128968 303858 129024
rect 303802 128308 303858 128344
rect 303802 128288 303804 128308
rect 303804 128288 303856 128308
rect 303856 128288 303858 128308
rect 303618 127472 303674 127528
rect 302238 125160 302294 125216
rect 303710 124480 303766 124536
rect 303802 123664 303858 123720
rect 303710 122984 303766 123040
rect 289450 122168 289506 122224
rect 303618 122168 303674 122224
rect 289266 121896 289322 121952
rect 289174 79328 289230 79384
rect 303802 121388 303804 121408
rect 303804 121388 303856 121408
rect 303856 121388 303858 121408
rect 303802 121352 303858 121388
rect 303802 119176 303858 119232
rect 303802 118396 303804 118416
rect 303804 118396 303856 118416
rect 303856 118396 303858 118416
rect 303802 118360 303858 118396
rect 303894 117544 303950 117600
rect 289726 116728 289782 116784
rect 303802 116048 303858 116104
rect 303618 115404 303620 115424
rect 303620 115404 303672 115424
rect 303672 115404 303674 115424
rect 303618 115368 303674 115404
rect 303802 114552 303858 114608
rect 303802 113736 303858 113792
rect 303802 113092 303804 113112
rect 303804 113092 303856 113112
rect 303856 113092 303858 113112
rect 303802 113056 303858 113092
rect 303710 112240 303766 112296
rect 303802 111560 303858 111616
rect 303710 110744 303766 110800
rect 305182 129784 305238 129840
rect 304722 125976 304778 126032
rect 304354 123392 304410 123448
rect 304262 108432 304318 108488
rect 303802 107752 303858 107808
rect 303802 106936 303858 106992
rect 303710 105440 303766 105496
rect 307942 202136 307998 202192
rect 307850 182824 307906 182880
rect 309230 285912 309286 285968
rect 309322 177248 309378 177304
rect 309322 143520 309378 143576
rect 309230 123392 309286 123448
rect 315946 287136 316002 287192
rect 315946 287000 316002 287056
rect 315946 277480 316002 277536
rect 315946 277344 316002 277400
rect 315946 267824 316002 267880
rect 315946 267688 316002 267744
rect 315946 248376 316002 248432
rect 315946 248240 316002 248296
rect 315946 238720 316002 238776
rect 315946 238584 316002 238640
rect 313462 134544 313518 134600
rect 316038 233824 316094 233880
rect 315946 229064 316002 229120
rect 315946 228928 316002 228984
rect 315946 219408 316002 219464
rect 315946 219272 316002 219328
rect 315946 209752 316002 209808
rect 315946 209616 316002 209672
rect 315946 200096 316002 200152
rect 315946 199960 316002 200016
rect 315946 190440 316002 190496
rect 315946 190304 316002 190360
rect 314934 182960 314990 183016
rect 315946 180784 316002 180840
rect 315946 180648 316002 180704
rect 315946 171128 316002 171184
rect 315946 170992 316002 171048
rect 315946 161472 316002 161528
rect 315946 161336 316002 161392
rect 315946 151816 316002 151872
rect 315946 151680 316002 151736
rect 315946 142160 316002 142216
rect 315946 142024 316002 142080
rect 315946 132504 316002 132560
rect 315946 132368 316002 132424
rect 315946 122848 316002 122904
rect 315946 122712 316002 122768
rect 315946 119312 316002 119368
rect 304354 104624 304410 104680
rect 303802 103944 303858 104000
rect 303618 103128 303674 103184
rect 303710 101632 303766 101688
rect 289818 94832 289874 94888
rect 291106 95648 291162 95704
rect 289818 76744 289874 76800
rect 289266 75112 289322 75168
rect 289818 72392 289874 72448
rect 285678 24112 285734 24168
rect 288990 11600 289046 11656
rect 299478 91704 299534 91760
rect 298742 88984 298798 89040
rect 292578 12960 292634 13016
rect 294878 3440 294934 3496
rect 296718 26832 296774 26888
rect 298098 11600 298154 11656
rect 301318 100544 301374 100600
rect 301502 99592 301558 99648
rect 301410 97280 301466 97336
rect 301318 96600 301374 96656
rect 301318 95104 301374 95160
rect 303618 99320 303674 99376
rect 302238 98504 302294 98560
rect 301410 94968 301466 95024
rect 302238 93608 302294 93664
rect 303894 96328 303950 96384
rect 304262 90344 304318 90400
rect 299570 73752 299626 73808
rect 311898 65456 311954 65512
rect 307758 33768 307814 33824
rect 310518 29552 310574 29608
rect 310242 8880 310298 8936
rect 307942 3440 307998 3496
rect 313830 6976 313886 7032
rect 317326 3984 317382 4040
rect 317602 213152 317658 213208
rect 318798 203496 318854 203552
rect 318982 220088 319038 220144
rect 320178 190984 320234 191040
rect 318522 1944 318578 2000
rect 320454 181464 320510 181520
rect 322202 195200 322258 195256
rect 324318 218592 324374 218648
rect 323030 204992 323086 205048
rect 323214 179968 323270 180024
rect 324962 300872 325018 300928
rect 324502 184184 324558 184240
rect 325790 230560 325846 230616
rect 324410 47504 324466 47560
rect 320914 3440 320970 3496
rect 322110 3440 322166 3496
rect 328458 267008 328514 267064
rect 327354 186904 327410 186960
rect 329838 200640 329894 200696
rect 329194 4800 329250 4856
rect 582378 365064 582434 365120
rect 580170 351872 580226 351928
rect 340878 350512 340934 350568
rect 338118 343712 338174 343768
rect 333978 324944 334034 325000
rect 332690 228248 332746 228304
rect 332598 207576 332654 207632
rect 335450 211792 335506 211848
rect 336738 215328 336794 215384
rect 339498 338136 339554 338192
rect 339590 309168 339646 309224
rect 582378 345616 582434 345672
rect 353298 222808 353354 222864
rect 342258 214512 342314 214568
rect 345018 206216 345074 206272
rect 351918 199280 351974 199336
rect 344558 3304 344614 3360
rect 351642 3576 351698 3632
rect 348054 3440 348110 3496
rect 356058 221448 356114 221504
rect 582378 334056 582434 334112
rect 358818 196560 358874 196616
rect 574742 299512 574798 299568
rect 580262 272176 580318 272232
rect 580170 245520 580226 245576
rect 580170 240080 580226 240136
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580906 125976 580962 126032
rect 583022 418240 583078 418296
rect 582838 378392 582894 378448
rect 582746 298696 582802 298752
rect 582930 302232 582986 302288
rect 582838 237904 582894 237960
rect 582746 237224 582802 237280
rect 582654 232328 582710 232384
rect 582562 72936 582618 72992
rect 582470 19760 582526 19816
rect 358818 3576 358874 3632
rect 357438 3440 357494 3496
rect 583390 404912 583446 404968
rect 583298 325216 583354 325272
rect 583114 312024 583170 312080
rect 583022 289040 583078 289096
rect 583022 284280 583078 284336
rect 583114 264152 583170 264208
rect 583022 258848 583078 258904
rect 582930 112784 582986 112840
rect 583482 304952 583538 305008
rect 583390 291760 583446 291816
rect 583298 229744 583354 229800
rect 583206 139304 583262 139360
rect 583114 99456 583170 99512
rect 583666 303592 583722 303648
rect 583482 219272 583538 219328
rect 583482 208936 583538 208992
rect 583390 152632 583446 152688
rect 583298 86128 583354 86184
rect 583022 59608 583078 59664
rect 582838 46280 582894 46336
rect 582746 33088 582802 33144
rect 582654 6568 582710 6624
rect 583574 202952 583630 203008
rect 356058 3304 356114 3360
rect 583758 206216 583814 206272
rect 583666 193024 583722 193080
<< metal3 >>
rect 69606 702476 69612 702540
rect 69676 702538 69682 702540
rect 154113 702538 154179 702541
rect 69676 702536 154179 702538
rect 69676 702480 154118 702536
rect 154174 702480 154179 702536
rect 69676 702478 154179 702480
rect 69676 702476 69682 702478
rect 154113 702475 154179 702478
rect 72969 699818 73035 699821
rect 76046 699818 76052 699820
rect 72969 699816 76052 699818
rect 72969 699760 72974 699816
rect 73030 699760 76052 699816
rect 72969 699758 76052 699760
rect 72969 699755 73035 699758
rect 76046 699756 76052 699758
rect 76116 699756 76122 699820
rect -960 697220 480 697460
rect 582373 697234 582439 697237
rect 583520 697234 584960 697324
rect 582373 697232 584960 697234
rect 582373 697176 582378 697232
rect 582434 697176 584960 697232
rect 582373 697174 584960 697176
rect 582373 697171 582439 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 582465 683906 582531 683909
rect 583520 683906 584960 683996
rect 582465 683904 584960 683906
rect 582465 683848 582470 683904
rect 582526 683848 584960 683904
rect 582465 683846 584960 683848
rect 582465 683843 582531 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580257 670714 580323 670717
rect 583520 670714 584960 670804
rect 580257 670712 584960 670714
rect 580257 670656 580262 670712
rect 580318 670656 584960 670712
rect 580257 670654 584960 670656
rect 580257 670651 580323 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 2773 658202 2839 658205
rect -960 658200 2839 658202
rect -960 658144 2778 658200
rect 2834 658144 2839 658200
rect -960 658142 2839 658144
rect -960 658052 480 658142
rect 2773 658139 2839 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 582557 644058 582623 644061
rect 583520 644058 584960 644148
rect 582557 644056 584960 644058
rect 582557 644000 582562 644056
rect 582618 644000 584960 644056
rect 582557 643998 584960 644000
rect 582557 643995 582623 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 582649 630866 582715 630869
rect 583520 630866 584960 630956
rect 582649 630864 584960 630866
rect 582649 630808 582654 630864
rect 582710 630808 584960 630864
rect 582649 630806 584960 630808
rect 582649 630803 582715 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 582741 617538 582807 617541
rect 583520 617538 584960 617628
rect 582741 617536 584960 617538
rect 582741 617480 582746 617536
rect 582802 617480 584960 617536
rect 582741 617478 584960 617480
rect 582741 617475 582807 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 83457 592106 83523 592109
rect 110413 592106 110479 592109
rect 83457 592104 110479 592106
rect 83457 592048 83462 592104
rect 83518 592048 110418 592104
rect 110474 592048 110479 592104
rect 83457 592046 110479 592048
rect 83457 592043 83523 592046
rect 110413 592043 110479 592046
rect 72417 591018 72483 591021
rect 83733 591018 83799 591021
rect 72417 591016 83799 591018
rect 72417 590960 72422 591016
rect 72478 590960 83738 591016
rect 83794 590960 83799 591016
rect 72417 590958 83799 590960
rect 72417 590955 72483 590958
rect 83733 590955 83799 590958
rect 86861 591018 86927 591021
rect 112437 591018 112503 591021
rect 86861 591016 112503 591018
rect 86861 590960 86866 591016
rect 86922 590960 112442 591016
rect 112498 590960 112503 591016
rect 86861 590958 112503 590960
rect 86861 590955 86927 590958
rect 112437 590955 112503 590958
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 61929 590882 61995 590885
rect 71037 590882 71103 590885
rect 61929 590880 71103 590882
rect 61929 590824 61934 590880
rect 61990 590824 71042 590880
rect 71098 590824 71103 590880
rect 61929 590822 71103 590824
rect 61929 590819 61995 590822
rect 71037 590819 71103 590822
rect 82537 590882 82603 590885
rect 107009 590882 107075 590885
rect 82537 590880 107075 590882
rect 82537 590824 82542 590880
rect 82598 590824 107014 590880
rect 107070 590824 107075 590880
rect 583520 590868 584960 590958
rect 82537 590822 107075 590824
rect 82537 590819 82603 590822
rect 107009 590819 107075 590822
rect 53649 590746 53715 590749
rect 73613 590746 73679 590749
rect 53649 590744 73679 590746
rect 53649 590688 53654 590744
rect 53710 590688 73618 590744
rect 73674 590688 73679 590744
rect 53649 590686 73679 590688
rect 53649 590683 53715 590686
rect 73613 590683 73679 590686
rect 77017 590746 77083 590749
rect 82629 590746 82695 590749
rect 77017 590744 82695 590746
rect 77017 590688 77022 590744
rect 77078 590688 82634 590744
rect 82690 590688 82695 590744
rect 77017 590686 82695 590688
rect 77017 590683 77083 590686
rect 82629 590683 82695 590686
rect 81341 590610 81407 590613
rect 88977 590610 89043 590613
rect 81341 590608 89043 590610
rect 81341 590552 81346 590608
rect 81402 590552 88982 590608
rect 89038 590552 89043 590608
rect 81341 590550 89043 590552
rect 81341 590547 81407 590550
rect 88977 590547 89043 590550
rect 67725 589930 67791 589933
rect 580165 589930 580231 589933
rect 67725 589928 580231 589930
rect 67725 589872 67730 589928
rect 67786 589872 580170 589928
rect 580226 589872 580231 589928
rect 67725 589870 580231 589872
rect 67725 589867 67791 589870
rect 580165 589867 580231 589870
rect 75637 588842 75703 588845
rect 86953 588842 87019 588845
rect 101397 588842 101463 588845
rect 75637 588840 80070 588842
rect 75637 588784 75642 588840
rect 75698 588784 80070 588840
rect 75637 588782 80070 588784
rect 75637 588779 75703 588782
rect 80010 588706 80070 588782
rect 86953 588840 101463 588842
rect 86953 588784 86958 588840
rect 87014 588784 101402 588840
rect 101458 588784 101463 588840
rect 86953 588782 101463 588784
rect 86953 588779 87019 588782
rect 101397 588779 101463 588782
rect 98637 588706 98703 588709
rect 80010 588704 98703 588706
rect 80010 588648 98642 588704
rect 98698 588648 98703 588704
rect 80010 588646 98703 588648
rect 98637 588643 98703 588646
rect 88057 588570 88123 588573
rect 88190 588570 88196 588572
rect 88057 588568 88196 588570
rect 88057 588512 88062 588568
rect 88118 588512 88196 588568
rect 88057 588510 88196 588512
rect 88057 588507 88123 588510
rect 88190 588508 88196 588510
rect 88260 588508 88266 588572
rect 66805 588298 66871 588301
rect 68878 588298 68938 588472
rect 66805 588296 68938 588298
rect 66805 588240 66810 588296
rect 66866 588240 68938 588296
rect 66805 588238 68938 588240
rect 66805 588235 66871 588238
rect 66253 586530 66319 586533
rect 66253 586528 66362 586530
rect 66253 586472 66258 586528
rect 66314 586472 66362 586528
rect 66253 586467 66362 586472
rect 66302 586394 66362 586467
rect 68878 586394 68938 587112
rect 88566 586938 88626 587656
rect 88566 586878 96630 586938
rect 66302 586334 68938 586394
rect 96570 586394 96630 586878
rect 159214 586468 159220 586532
rect 159284 586468 159290 586532
rect 159222 586394 159282 586468
rect 96570 586334 159282 586394
rect 67725 585850 67791 585853
rect 88566 585850 88626 586296
rect 89897 585850 89963 585853
rect 67725 585848 68938 585850
rect 67725 585792 67730 585848
rect 67786 585792 68938 585848
rect 67725 585790 68938 585792
rect 88566 585848 89963 585850
rect 88566 585792 89902 585848
rect 89958 585792 89963 585848
rect 88566 585790 89963 585792
rect 67725 585787 67791 585790
rect 68878 585752 68938 585790
rect 89897 585787 89963 585790
rect 88190 585652 88196 585716
rect 88260 585714 88266 585716
rect 118693 585714 118759 585717
rect 88260 585712 118759 585714
rect 88260 585656 118698 585712
rect 118754 585656 118759 585712
rect 88260 585654 118759 585656
rect 88260 585652 88266 585654
rect 118693 585651 118759 585654
rect 88566 584626 88626 584936
rect 91921 584626 91987 584629
rect 88566 584624 91987 584626
rect 88566 584568 91926 584624
rect 91982 584568 91987 584624
rect 88566 584566 91987 584568
rect 91921 584563 91987 584566
rect 67766 583748 67772 583812
rect 67836 583810 67842 583812
rect 68878 583810 68938 584392
rect 67836 583750 68938 583810
rect 67836 583748 67842 583750
rect 91829 583674 91895 583677
rect 88566 583672 91895 583674
rect 88566 583616 91834 583672
rect 91890 583616 91895 583672
rect 88566 583614 91895 583616
rect 88566 583576 88626 583614
rect 91829 583611 91895 583614
rect 66805 582450 66871 582453
rect 68878 582450 68938 583032
rect 88977 582994 89043 582997
rect 123477 582994 123543 582997
rect 88977 582992 123543 582994
rect 88977 582936 88982 582992
rect 89038 582936 123482 582992
rect 123538 582936 123543 582992
rect 88977 582934 123543 582936
rect 88977 582931 89043 582934
rect 123477 582931 123543 582934
rect 66805 582448 68938 582450
rect 66805 582392 66810 582448
rect 66866 582392 68938 582448
rect 66805 582390 68938 582392
rect 66805 582387 66871 582390
rect 69422 581844 69428 581908
rect 69492 581844 69498 581908
rect 69430 581702 69490 581844
rect 68908 581672 69490 581702
rect 68878 581642 69460 581672
rect 66069 581634 66135 581637
rect 68878 581634 68938 581642
rect 66069 581632 68938 581634
rect 66069 581576 66074 581632
rect 66130 581576 68938 581632
rect 66069 581574 68938 581576
rect 88566 581634 88626 582216
rect 91093 581634 91159 581637
rect 88566 581632 91159 581634
rect 88566 581576 91098 581632
rect 91154 581576 91159 581632
rect 88566 581574 91159 581576
rect 66069 581571 66135 581574
rect 91093 581571 91159 581574
rect 97901 580954 97967 580957
rect 88566 580952 97967 580954
rect 88566 580896 97906 580952
rect 97962 580896 97967 580952
rect 88566 580894 97967 580896
rect 88566 580856 88626 580894
rect 97901 580891 97967 580894
rect -960 580002 480 580092
rect 2773 580002 2839 580005
rect -960 580000 2839 580002
rect -960 579944 2778 580000
rect 2834 579944 2839 580000
rect -960 579942 2839 579944
rect -960 579852 480 579942
rect 2773 579939 2839 579942
rect 66805 579730 66871 579733
rect 68878 579730 68938 580312
rect 97901 580274 97967 580277
rect 119470 580274 119476 580276
rect 97901 580272 119476 580274
rect 97901 580216 97906 580272
rect 97962 580216 119476 580272
rect 97901 580214 119476 580216
rect 97901 580211 97967 580214
rect 119470 580212 119476 580214
rect 119540 580212 119546 580276
rect 66805 579728 68938 579730
rect 66805 579672 66810 579728
rect 66866 579672 68938 579728
rect 66805 579670 68938 579672
rect 66805 579667 66871 579670
rect 67725 578370 67791 578373
rect 68878 578370 68938 578952
rect 88566 578914 88626 579496
rect 91093 578914 91159 578917
rect 88566 578912 91159 578914
rect 88566 578856 91098 578912
rect 91154 578856 91159 578912
rect 88566 578854 91159 578856
rect 91093 578851 91159 578854
rect 67725 578368 68938 578370
rect 67725 578312 67730 578368
rect 67786 578312 68938 578368
rect 67725 578310 68938 578312
rect 67725 578307 67791 578310
rect 67817 577010 67883 577013
rect 68878 577010 68938 577592
rect 88566 577554 88626 578136
rect 580257 577690 580323 577693
rect 583520 577690 584960 577780
rect 580257 577688 584960 577690
rect 580257 577632 580262 577688
rect 580318 577632 584960 577688
rect 580257 577630 584960 577632
rect 580257 577627 580323 577630
rect 91093 577554 91159 577557
rect 88566 577552 91159 577554
rect 88566 577496 91098 577552
rect 91154 577496 91159 577552
rect 583520 577540 584960 577630
rect 88566 577494 91159 577496
rect 91093 577491 91159 577494
rect 67817 577008 68938 577010
rect 67817 576952 67822 577008
rect 67878 576952 68938 577008
rect 67817 576950 68938 576952
rect 67817 576947 67883 576950
rect 88566 576738 88626 576776
rect 91185 576738 91251 576741
rect 88566 576736 91251 576738
rect 88566 576680 91190 576736
rect 91246 576680 91251 576736
rect 88566 576678 91251 576680
rect 91185 576675 91251 576678
rect 66897 575650 66963 575653
rect 68878 575650 68938 576232
rect 66897 575648 68938 575650
rect 66897 575592 66902 575648
rect 66958 575592 68938 575648
rect 66897 575590 68938 575592
rect 66897 575587 66963 575590
rect 67449 575378 67515 575381
rect 67449 575376 68938 575378
rect 67449 575320 67454 575376
rect 67510 575320 68938 575376
rect 67449 575318 68938 575320
rect 67449 575315 67515 575318
rect 68878 574872 68938 575318
rect 88566 575106 88626 575416
rect 91093 575106 91159 575109
rect 88566 575104 91159 575106
rect 88566 575048 91098 575104
rect 91154 575048 91159 575104
rect 88566 575046 91159 575048
rect 91093 575043 91159 575046
rect 65977 572930 66043 572933
rect 68878 572930 68938 573512
rect 88566 573474 88626 574056
rect 91093 573474 91159 573477
rect 88566 573472 91159 573474
rect 88566 573416 91098 573472
rect 91154 573416 91159 573472
rect 88566 573414 91159 573416
rect 91093 573411 91159 573414
rect 65977 572928 68938 572930
rect 65977 572872 65982 572928
rect 66038 572872 68938 572928
rect 65977 572870 68938 572872
rect 65977 572867 66043 572870
rect 66437 571842 66503 571845
rect 68878 571842 68938 572152
rect 88566 572114 88626 572696
rect 91185 572114 91251 572117
rect 88566 572112 91251 572114
rect 88566 572056 91190 572112
rect 91246 572056 91251 572112
rect 88566 572054 91251 572056
rect 91185 572051 91251 572054
rect 66437 571840 68938 571842
rect 66437 571784 66442 571840
rect 66498 571784 68938 571840
rect 66437 571782 68938 571784
rect 66437 571779 66503 571782
rect 91093 571434 91159 571437
rect 88566 571432 91159 571434
rect 88566 571376 91098 571432
rect 91154 571376 91159 571432
rect 88566 571374 91159 571376
rect 88566 571336 88626 571374
rect 91093 571371 91159 571374
rect 67357 570210 67423 570213
rect 68878 570210 68938 570792
rect 67357 570208 68938 570210
rect 67357 570152 67362 570208
rect 67418 570152 68938 570208
rect 67357 570150 68938 570152
rect 67357 570147 67423 570150
rect 91093 570074 91159 570077
rect 88566 570072 91159 570074
rect 88566 570016 91098 570072
rect 91154 570016 91159 570072
rect 88566 570014 91159 570016
rect 88566 569976 88626 570014
rect 91093 570011 91159 570014
rect 66897 568850 66963 568853
rect 68878 568850 68938 569432
rect 66897 568848 68938 568850
rect 66897 568792 66902 568848
rect 66958 568792 68938 568848
rect 66897 568790 68938 568792
rect 66897 568787 66963 568790
rect 92197 568714 92263 568717
rect 88566 568712 92263 568714
rect 88566 568656 92202 568712
rect 92258 568656 92263 568712
rect 88566 568654 92263 568656
rect 88566 568616 88626 568654
rect 92197 568651 92263 568654
rect 66897 567490 66963 567493
rect 68878 567490 68938 568072
rect 66897 567488 68938 567490
rect 66897 567432 66902 567488
rect 66958 567432 68938 567488
rect 66897 567430 68938 567432
rect 66897 567427 66963 567430
rect 88885 567286 88951 567289
rect 88596 567284 88951 567286
rect 88596 567228 88890 567284
rect 88946 567228 88951 567284
rect 88596 567226 88951 567228
rect 88885 567223 88951 567226
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 67541 566810 67607 566813
rect 67541 566808 68938 566810
rect 67541 566752 67546 566808
rect 67602 566752 68938 566808
rect 67541 566750 68938 566752
rect 67541 566747 67607 566750
rect 68878 566712 68938 566750
rect 88566 565858 88626 565896
rect 91093 565858 91159 565861
rect 88566 565856 91159 565858
rect 88566 565800 91098 565856
rect 91154 565800 91159 565856
rect 88566 565798 91159 565800
rect 91093 565795 91159 565798
rect 65517 564498 65583 564501
rect 68878 564498 68938 565080
rect 65517 564496 68938 564498
rect 65517 564440 65522 564496
rect 65578 564440 68938 564496
rect 65517 564438 68938 564440
rect 88566 564498 88626 564536
rect 91737 564498 91803 564501
rect 88566 564496 91803 564498
rect 88566 564440 91742 564496
rect 91798 564440 91803 564496
rect 88566 564438 91803 564440
rect 65517 564435 65583 564438
rect 91737 564435 91803 564438
rect 66805 564362 66871 564365
rect 582741 564362 582807 564365
rect 583520 564362 584960 564452
rect 66805 564360 68938 564362
rect 66805 564304 66810 564360
rect 66866 564304 68938 564360
rect 66805 564302 68938 564304
rect 66805 564299 66871 564302
rect 68878 563720 68938 564302
rect 582741 564360 584960 564362
rect 582741 564304 582746 564360
rect 582802 564304 584960 564360
rect 582741 564302 584960 564304
rect 582741 564299 582807 564302
rect 583520 564212 584960 564302
rect 88566 563138 88626 563176
rect 91093 563138 91159 563141
rect 88566 563136 91159 563138
rect 88566 563080 91098 563136
rect 91154 563080 91159 563136
rect 88566 563078 91159 563080
rect 91093 563075 91159 563078
rect 66805 561778 66871 561781
rect 68878 561778 68938 562360
rect 66805 561776 68938 561778
rect 66805 561720 66810 561776
rect 66866 561720 68938 561776
rect 66805 561718 68938 561720
rect 66805 561715 66871 561718
rect 66529 560554 66595 560557
rect 68878 560554 68938 561000
rect 88566 560962 88626 561544
rect 91093 560962 91159 560965
rect 88566 560960 91159 560962
rect 88566 560904 91098 560960
rect 91154 560904 91159 560960
rect 88566 560902 91159 560904
rect 91093 560899 91159 560902
rect 66529 560552 68938 560554
rect 66529 560496 66534 560552
rect 66590 560496 68938 560552
rect 66529 560494 68938 560496
rect 66529 560491 66595 560494
rect 88566 560146 88626 560184
rect 89805 560146 89871 560149
rect 91829 560146 91895 560149
rect 88566 560144 91895 560146
rect 88566 560088 89810 560144
rect 89866 560088 91834 560144
rect 91890 560088 91895 560144
rect 88566 560086 91895 560088
rect 89805 560083 89871 560086
rect 91829 560083 91895 560086
rect 66529 559194 66595 559197
rect 68878 559194 68938 559640
rect 66529 559192 68938 559194
rect 66529 559136 66534 559192
rect 66590 559136 68938 559192
rect 66529 559134 68938 559136
rect 66529 559131 66595 559134
rect 67633 558922 67699 558925
rect 67633 558920 68938 558922
rect 67633 558864 67638 558920
rect 67694 558864 68938 558920
rect 67633 558862 68938 558864
rect 67633 558859 67699 558862
rect 68878 558280 68938 558862
rect 88566 558242 88626 558824
rect 91185 558242 91251 558245
rect 88566 558240 91251 558242
rect 88566 558184 91190 558240
rect 91246 558184 91251 558240
rect 88566 558182 91251 558184
rect 91185 558179 91251 558182
rect 66897 556338 66963 556341
rect 68878 556338 68938 556920
rect 88566 556882 88626 557464
rect 91185 556882 91251 556885
rect 88566 556880 91251 556882
rect 88566 556824 91190 556880
rect 91246 556824 91251 556880
rect 88566 556822 91251 556824
rect 91185 556819 91251 556822
rect 66897 556336 68938 556338
rect 66897 556280 66902 556336
rect 66958 556280 68938 556336
rect 66897 556278 68938 556280
rect 66897 556275 66963 556278
rect 66621 554978 66687 554981
rect 68878 554978 68938 555560
rect 88566 555522 88626 556104
rect 91185 555522 91251 555525
rect 88566 555520 91251 555522
rect 88566 555464 91190 555520
rect 91246 555464 91251 555520
rect 88566 555462 91251 555464
rect 91185 555459 91251 555462
rect 66621 554976 68938 554978
rect 66621 554920 66626 554976
rect 66682 554920 68938 554976
rect 66621 554918 68938 554920
rect 66621 554915 66687 554918
rect -960 553890 480 553980
rect 3509 553890 3575 553893
rect -960 553888 3575 553890
rect -960 553832 3514 553888
rect 3570 553832 3575 553888
rect -960 553830 3575 553832
rect -960 553740 480 553830
rect 3509 553827 3575 553830
rect 66529 553754 66595 553757
rect 68878 553754 68938 554200
rect 88566 554026 88626 554744
rect 88566 553966 93870 554026
rect 66529 553752 68938 553754
rect 66529 553696 66534 553752
rect 66590 553696 68938 553752
rect 66529 553694 68938 553696
rect 66529 553691 66595 553694
rect 93810 553482 93870 553966
rect 111006 553482 111012 553484
rect 93810 553422 111012 553482
rect 111006 553420 111012 553422
rect 111076 553420 111082 553484
rect 88566 552938 88626 553384
rect 91185 552938 91251 552941
rect 88566 552936 91251 552938
rect 88566 552880 91190 552936
rect 91246 552880 91251 552936
rect 88566 552878 91251 552880
rect 91185 552875 91251 552878
rect 67449 552258 67515 552261
rect 68878 552258 68938 552840
rect 67449 552256 68938 552258
rect 67449 552200 67454 552256
rect 67510 552200 68938 552256
rect 67449 552198 68938 552200
rect 67449 552195 67515 552198
rect 91185 552122 91251 552125
rect 88566 552120 91251 552122
rect 88566 552064 91190 552120
rect 91246 552064 91251 552120
rect 88566 552062 91251 552064
rect 88566 552024 88626 552062
rect 91185 552059 91251 552062
rect 66662 550836 66668 550900
rect 66732 550898 66738 550900
rect 68878 550898 68938 551480
rect 583520 551020 584960 551260
rect 66732 550838 68938 550898
rect 66732 550836 66738 550838
rect 99966 550762 99972 550764
rect 88566 550702 99972 550762
rect 88566 550664 88626 550702
rect 99966 550700 99972 550702
rect 100036 550700 100042 550764
rect 66437 549674 66503 549677
rect 68878 549674 68938 550120
rect 66437 549672 68938 549674
rect 66437 549616 66442 549672
rect 66498 549616 68938 549672
rect 66437 549614 68938 549616
rect 66437 549611 66503 549614
rect 91185 549402 91251 549405
rect 88566 549400 91251 549402
rect 88566 549344 91190 549400
rect 91246 549344 91251 549400
rect 88566 549342 91251 549344
rect 88566 549304 88626 549342
rect 91185 549339 91251 549342
rect 66529 548314 66595 548317
rect 68878 548314 68938 548760
rect 66529 548312 68938 548314
rect 66529 548256 66534 548312
rect 66590 548256 68938 548312
rect 66529 548254 68938 548256
rect 66529 548251 66595 548254
rect 88566 547906 88626 547944
rect 91277 547906 91343 547909
rect 88566 547904 91343 547906
rect 88566 547848 91282 547904
rect 91338 547848 91343 547904
rect 88566 547846 91343 547848
rect 91277 547843 91343 547846
rect 66621 547634 66687 547637
rect 66621 547632 68938 547634
rect 66621 547576 66626 547632
rect 66682 547576 68938 547632
rect 66621 547574 68938 547576
rect 66621 547571 66687 547574
rect 68878 547400 68938 547574
rect 88566 546546 88626 546584
rect 91369 546546 91435 546549
rect 109350 546546 109356 546548
rect 88566 546544 109356 546546
rect 88566 546488 91374 546544
rect 91430 546488 109356 546544
rect 88566 546486 109356 546488
rect 91369 546483 91435 546486
rect 109350 546484 109356 546486
rect 109420 546484 109426 546548
rect 66161 546410 66227 546413
rect 66161 546408 68938 546410
rect 66161 546352 66166 546408
rect 66222 546352 68938 546408
rect 66161 546350 68938 546352
rect 66161 546347 66227 546350
rect 68878 546040 68938 546350
rect 89989 545322 90055 545325
rect 88566 545320 90055 545322
rect 88566 545264 89994 545320
rect 90050 545264 90055 545320
rect 88566 545262 90055 545264
rect 88566 545224 88626 545262
rect 89989 545259 90055 545262
rect 66805 544098 66871 544101
rect 68878 544098 68938 544680
rect 91185 544098 91251 544101
rect 66805 544096 68938 544098
rect 66805 544040 66810 544096
rect 66866 544040 68938 544096
rect 66805 544038 68938 544040
rect 88566 544096 91251 544098
rect 88566 544040 91190 544096
rect 91246 544040 91251 544096
rect 88566 544038 91251 544040
rect 66805 544035 66871 544038
rect 88566 543864 88626 544038
rect 91185 544035 91251 544038
rect 66805 542738 66871 542741
rect 68878 542738 68938 543320
rect 66805 542736 68938 542738
rect 66805 542680 66810 542736
rect 66866 542680 68938 542736
rect 66805 542678 68938 542680
rect 66805 542675 66871 542678
rect 88566 542466 88626 542504
rect 91185 542466 91251 542469
rect 88566 542464 91251 542466
rect 88566 542408 91190 542464
rect 91246 542408 91251 542464
rect 88566 542406 91251 542408
rect 91185 542403 91251 542406
rect 67081 541786 67147 541789
rect 68878 541786 68938 541960
rect 67081 541784 68938 541786
rect 67081 541728 67086 541784
rect 67142 541728 68938 541784
rect 67081 541726 68938 541728
rect 67081 541723 67147 541726
rect 91185 541378 91251 541381
rect 88566 541376 91251 541378
rect 88566 541320 91190 541376
rect 91246 541320 91251 541376
rect 88566 541318 91251 541320
rect 88566 541144 88626 541318
rect 91185 541315 91251 541318
rect -960 540684 480 540924
rect 68645 540834 68711 540837
rect 68645 540832 68938 540834
rect 68645 540776 68650 540832
rect 68706 540776 68938 540832
rect 68645 540774 68938 540776
rect 68645 540771 68711 540774
rect 68878 540600 68938 540774
rect 88566 539746 88626 539784
rect 91185 539746 91251 539749
rect 88566 539744 91251 539746
rect 88566 539688 91190 539744
rect 91246 539688 91251 539744
rect 88566 539686 91251 539688
rect 91185 539683 91251 539686
rect 76046 538052 76052 538116
rect 76116 538114 76122 538116
rect 76741 538114 76807 538117
rect 76116 538112 76807 538114
rect 76116 538056 76746 538112
rect 76802 538056 76807 538112
rect 76116 538054 76807 538056
rect 76116 538052 76122 538054
rect 76741 538051 76807 538054
rect 579797 537842 579863 537845
rect 583520 537842 584960 537932
rect 579797 537840 584960 537842
rect 579797 537784 579802 537840
rect 579858 537784 584960 537840
rect 579797 537782 584960 537784
rect 579797 537779 579863 537782
rect 583520 537692 584960 537782
rect 76465 536754 76531 536757
rect 124857 536754 124923 536757
rect 76465 536752 124923 536754
rect 76465 536696 76470 536752
rect 76526 536696 124862 536752
rect 124918 536696 124923 536752
rect 76465 536694 124923 536696
rect 76465 536691 76531 536694
rect 124857 536691 124923 536694
rect 84745 536074 84811 536077
rect 128997 536074 129063 536077
rect 582373 536074 582439 536077
rect 84745 536072 582439 536074
rect 84745 536016 84750 536072
rect 84806 536016 129002 536072
rect 129058 536016 582378 536072
rect 582434 536016 582439 536072
rect 84745 536014 582439 536016
rect 84745 536011 84811 536014
rect 128997 536011 129063 536014
rect 582373 536011 582439 536014
rect 69657 535532 69723 535533
rect 69606 535468 69612 535532
rect 69676 535530 69723 535532
rect 70669 535530 70735 535533
rect 71814 535530 71820 535532
rect 69676 535528 69768 535530
rect 69718 535472 69768 535528
rect 69676 535470 69768 535472
rect 70669 535528 71820 535530
rect 70669 535472 70674 535528
rect 70730 535472 71820 535528
rect 70669 535470 71820 535472
rect 69676 535468 69723 535470
rect 69657 535467 69723 535468
rect 70669 535467 70735 535470
rect 71814 535468 71820 535470
rect 71884 535468 71890 535532
rect 75913 535530 75979 535533
rect 76741 535530 76807 535533
rect 75913 535528 76807 535530
rect 75913 535472 75918 535528
rect 75974 535472 76746 535528
rect 76802 535472 76807 535528
rect 75913 535470 76807 535472
rect 75913 535467 75979 535470
rect 76741 535467 76807 535470
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 582465 524514 582531 524517
rect 583520 524514 584960 524604
rect 582465 524512 584960 524514
rect 582465 524456 582470 524512
rect 582526 524456 584960 524512
rect 582465 524454 584960 524456
rect 582465 524451 582531 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 2773 501802 2839 501805
rect -960 501800 2839 501802
rect -960 501744 2778 501800
rect 2834 501744 2839 501800
rect -960 501742 2839 501744
rect -960 501652 480 501742
rect 2773 501739 2839 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 582373 484666 582439 484669
rect 583520 484666 584960 484756
rect 582373 484664 584960 484666
rect 582373 484608 582378 484664
rect 582434 484608 584960 484664
rect 582373 484606 584960 484608
rect 582373 484603 582439 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 582649 471474 582715 471477
rect 583520 471474 584960 471564
rect 582649 471472 584960 471474
rect 582649 471416 582654 471472
rect 582710 471416 584960 471472
rect 582649 471414 584960 471416
rect 582649 471411 582715 471414
rect 583520 471324 584960 471414
rect 93761 469842 93827 469845
rect 122598 469842 122604 469844
rect 93761 469840 122604 469842
rect 93761 469784 93766 469840
rect 93822 469784 122604 469840
rect 93761 469782 122604 469784
rect 93761 469779 93827 469782
rect 122598 469780 122604 469782
rect 122668 469780 122674 469844
rect 95141 467122 95207 467125
rect 106406 467122 106412 467124
rect 95141 467120 106412 467122
rect 95141 467064 95146 467120
rect 95202 467064 106412 467120
rect 95141 467062 106412 467064
rect 95141 467059 95207 467062
rect 106406 467060 106412 467062
rect 106476 467060 106482 467124
rect 86861 462906 86927 462909
rect 96838 462906 96844 462908
rect 86861 462904 96844 462906
rect 86861 462848 86866 462904
rect 86922 462848 96844 462904
rect 86861 462846 96844 462848
rect 86861 462843 86927 462846
rect 96838 462844 96844 462846
rect 96908 462844 96914 462908
rect 100661 462906 100727 462909
rect 120206 462906 120212 462908
rect 100661 462904 120212 462906
rect 100661 462848 100666 462904
rect 100722 462848 120212 462904
rect 100661 462846 120212 462848
rect 100661 462843 100727 462846
rect 120206 462844 120212 462846
rect 120276 462844 120282 462908
rect -960 462634 480 462724
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 81433 461546 81499 461549
rect 89662 461546 89668 461548
rect 81433 461544 89668 461546
rect 81433 461488 81438 461544
rect 81494 461488 89668 461544
rect 81433 461486 89668 461488
rect 81433 461483 81499 461486
rect 89662 461484 89668 461486
rect 89732 461484 89738 461548
rect 98729 461546 98795 461549
rect 111742 461546 111748 461548
rect 98729 461544 111748 461546
rect 98729 461488 98734 461544
rect 98790 461488 111748 461544
rect 98729 461486 111748 461488
rect 98729 461483 98795 461486
rect 111742 461484 111748 461486
rect 111812 461484 111818 461548
rect 84101 460186 84167 460189
rect 92606 460186 92612 460188
rect 84101 460184 92612 460186
rect 84101 460128 84106 460184
rect 84162 460128 92612 460184
rect 84101 460126 92612 460128
rect 84101 460123 84167 460126
rect 92606 460124 92612 460126
rect 92676 460124 92682 460188
rect 93117 460186 93183 460189
rect 102726 460186 102732 460188
rect 93117 460184 102732 460186
rect 93117 460128 93122 460184
rect 93178 460128 102732 460184
rect 93117 460126 102732 460128
rect 93117 460123 93183 460126
rect 102726 460124 102732 460126
rect 102796 460124 102802 460188
rect 104249 459642 104315 459645
rect 104934 459642 104940 459644
rect 104249 459640 104940 459642
rect 104249 459584 104254 459640
rect 104310 459584 104940 459640
rect 104249 459582 104940 459584
rect 104249 459579 104315 459582
rect 104934 459580 104940 459582
rect 105004 459580 105010 459644
rect 91001 458826 91067 458829
rect 107694 458826 107700 458828
rect 91001 458824 107700 458826
rect 91001 458768 91006 458824
rect 91062 458768 107700 458824
rect 91001 458766 107700 458768
rect 91001 458763 91067 458766
rect 107694 458764 107700 458766
rect 107764 458764 107770 458828
rect 582465 458146 582531 458149
rect 583520 458146 584960 458236
rect 582465 458144 584960 458146
rect 582465 458088 582470 458144
rect 582526 458088 584960 458144
rect 582465 458086 584960 458088
rect 582465 458083 582531 458086
rect 583520 457996 584960 458086
rect 67766 457404 67772 457468
rect 67836 457466 67842 457468
rect 82077 457466 82143 457469
rect 67836 457464 82143 457466
rect 67836 457408 82082 457464
rect 82138 457408 82143 457464
rect 67836 457406 82143 457408
rect 67836 457404 67842 457406
rect 82077 457403 82143 457406
rect 87045 457466 87111 457469
rect 98126 457466 98132 457468
rect 87045 457464 98132 457466
rect 87045 457408 87050 457464
rect 87106 457408 98132 457464
rect 87045 457406 98132 457408
rect 87045 457403 87111 457406
rect 98126 457404 98132 457406
rect 98196 457404 98202 457468
rect 82721 456242 82787 456245
rect 91134 456242 91140 456244
rect 82721 456240 91140 456242
rect 82721 456184 82726 456240
rect 82782 456184 91140 456240
rect 82721 456182 91140 456184
rect 82721 456179 82787 456182
rect 91134 456180 91140 456182
rect 91204 456180 91210 456244
rect 89621 456106 89687 456109
rect 100702 456106 100708 456108
rect 89621 456104 100708 456106
rect 89621 456048 89626 456104
rect 89682 456048 100708 456104
rect 89621 456046 100708 456048
rect 89621 456043 89687 456046
rect 100702 456044 100708 456046
rect 100772 456044 100778 456108
rect 106917 456106 106983 456109
rect 115974 456106 115980 456108
rect 106917 456104 115980 456106
rect 106917 456048 106922 456104
rect 106978 456048 115980 456104
rect 106917 456046 115980 456048
rect 106917 456043 106983 456046
rect 115974 456044 115980 456046
rect 116044 456044 116050 456108
rect 95877 455562 95943 455565
rect 148174 455562 148180 455564
rect 95877 455560 148180 455562
rect 95877 455504 95882 455560
rect 95938 455504 148180 455560
rect 95877 455502 148180 455504
rect 95877 455499 95943 455502
rect 148174 455500 148180 455502
rect 148244 455500 148250 455564
rect 91737 451890 91803 451893
rect 121678 451890 121684 451892
rect 91737 451888 121684 451890
rect 91737 451832 91742 451888
rect 91798 451832 121684 451888
rect 91737 451830 121684 451832
rect 91737 451827 91803 451830
rect 121678 451828 121684 451830
rect 121748 451828 121754 451892
rect 104157 450530 104223 450533
rect 123109 450530 123175 450533
rect 104157 450528 123175 450530
rect 104157 450472 104162 450528
rect 104218 450472 123114 450528
rect 123170 450472 123175 450528
rect 104157 450470 123175 450472
rect 104157 450467 104223 450470
rect 123109 450467 123175 450470
rect 172513 449988 172579 449989
rect 172462 449986 172468 449988
rect 172422 449926 172468 449986
rect 172532 449984 172579 449988
rect 172574 449928 172579 449984
rect 172462 449924 172468 449926
rect 172532 449924 172579 449928
rect 172513 449923 172579 449924
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 86217 449170 86283 449173
rect 95182 449170 95188 449172
rect 86217 449168 95188 449170
rect 86217 449112 86222 449168
rect 86278 449112 95188 449168
rect 86217 449110 95188 449112
rect 86217 449107 86283 449110
rect 95182 449108 95188 449110
rect 95252 449108 95258 449172
rect 65977 448626 66043 448629
rect 72417 448626 72483 448629
rect 65977 448624 72483 448626
rect 65977 448568 65982 448624
rect 66038 448568 72422 448624
rect 72478 448568 72483 448624
rect 65977 448566 72483 448568
rect 65977 448563 66043 448566
rect 72417 448563 72483 448566
rect 91553 448626 91619 448629
rect 160686 448626 160692 448628
rect 91553 448624 160692 448626
rect 91553 448568 91558 448624
rect 91614 448568 160692 448624
rect 91553 448566 160692 448568
rect 91553 448563 91619 448566
rect 160686 448564 160692 448566
rect 160756 448564 160762 448628
rect 108389 447810 108455 447813
rect 123017 447810 123083 447813
rect 108389 447808 123083 447810
rect 108389 447752 108394 447808
rect 108450 447752 123022 447808
rect 123078 447752 123083 447808
rect 108389 447750 123083 447752
rect 108389 447747 108455 447750
rect 123017 447747 123083 447750
rect 123334 447612 123340 447676
rect 123404 447674 123410 447676
rect 123477 447674 123543 447677
rect 123404 447672 132510 447674
rect 123404 447616 123482 447672
rect 123538 447616 132510 447672
rect 123404 447614 132510 447616
rect 123404 447612 123410 447614
rect 123477 447611 123543 447614
rect 132450 447402 132510 447614
rect 168465 447402 168531 447405
rect 132450 447400 168531 447402
rect 132450 447344 168470 447400
rect 168526 447344 168531 447400
rect 132450 447342 168531 447344
rect 168465 447339 168531 447342
rect 71773 447266 71839 447269
rect 130469 447266 130535 447269
rect 71773 447264 130535 447266
rect 71773 447208 71778 447264
rect 71834 447208 130474 447264
rect 130530 447208 130535 447264
rect 71773 447206 130535 447208
rect 71773 447203 71839 447206
rect 130469 447203 130535 447206
rect 95233 446450 95299 446453
rect 96470 446450 96476 446452
rect 95233 446448 96476 446450
rect 95233 446392 95238 446448
rect 95294 446392 96476 446448
rect 95233 446390 96476 446392
rect 95233 446387 95299 446390
rect 96470 446388 96476 446390
rect 96540 446388 96546 446452
rect 128261 446314 128327 446317
rect 128537 446314 128603 446317
rect 128261 446312 128603 446314
rect 128261 446256 128266 446312
rect 128322 446256 128542 446312
rect 128598 446256 128603 446312
rect 128261 446254 128603 446256
rect 128261 446251 128327 446254
rect 128537 446251 128603 446254
rect 53649 446042 53715 446045
rect 85573 446042 85639 446045
rect 53649 446040 85639 446042
rect 53649 445984 53654 446040
rect 53710 445984 85578 446040
rect 85634 445984 85639 446040
rect 53649 445982 85639 445984
rect 53649 445979 53715 445982
rect 85573 445979 85639 445982
rect 105537 446042 105603 446045
rect 202137 446042 202203 446045
rect 105537 446040 202203 446042
rect 105537 445984 105542 446040
rect 105598 445984 202142 446040
rect 202198 445984 202203 446040
rect 105537 445982 202203 445984
rect 105537 445979 105603 445982
rect 202137 445979 202203 445982
rect 55029 445906 55095 445909
rect 78673 445906 78739 445909
rect 55029 445904 78739 445906
rect 55029 445848 55034 445904
rect 55090 445848 78678 445904
rect 78734 445848 78739 445904
rect 55029 445846 78739 445848
rect 55029 445843 55095 445846
rect 78673 445843 78739 445846
rect 82077 445906 82143 445909
rect 90214 445906 90220 445908
rect 82077 445904 90220 445906
rect 82077 445848 82082 445904
rect 82138 445848 90220 445904
rect 82077 445846 90220 445848
rect 82077 445843 82143 445846
rect 90214 445844 90220 445846
rect 90284 445844 90290 445908
rect 116393 445906 116459 445909
rect 128261 445906 128327 445909
rect 116393 445904 128327 445906
rect 116393 445848 116398 445904
rect 116454 445848 128266 445904
rect 128322 445848 128327 445904
rect 116393 445846 128327 445848
rect 116393 445843 116459 445846
rect 128261 445843 128327 445846
rect 67817 445770 67883 445773
rect 68461 445770 68527 445773
rect 67817 445768 68527 445770
rect 67817 445712 67822 445768
rect 67878 445712 68466 445768
rect 68522 445712 68527 445768
rect 67817 445710 68527 445712
rect 67817 445707 67883 445710
rect 68461 445707 68527 445710
rect 93853 445770 93919 445773
rect 94497 445770 94563 445773
rect 96613 445772 96679 445773
rect 94998 445770 95004 445772
rect 93853 445768 95004 445770
rect 93853 445712 93858 445768
rect 93914 445712 94502 445768
rect 94558 445712 95004 445768
rect 93853 445710 95004 445712
rect 93853 445707 93919 445710
rect 94497 445707 94563 445710
rect 94998 445708 95004 445710
rect 95068 445708 95074 445772
rect 96613 445770 96660 445772
rect 96532 445768 96660 445770
rect 96724 445770 96730 445772
rect 97349 445770 97415 445773
rect 96724 445768 97415 445770
rect 96532 445712 96618 445768
rect 96724 445712 97354 445768
rect 97410 445712 97415 445768
rect 96532 445710 96660 445712
rect 96613 445708 96660 445710
rect 96724 445710 97415 445712
rect 96724 445708 96730 445710
rect 96613 445707 96679 445708
rect 97349 445707 97415 445710
rect 99046 445708 99052 445772
rect 99116 445770 99122 445772
rect 102133 445770 102199 445773
rect 99116 445768 102199 445770
rect 99116 445712 102138 445768
rect 102194 445712 102199 445768
rect 99116 445710 102199 445712
rect 99116 445708 99122 445710
rect 102133 445707 102199 445710
rect 110413 445770 110479 445773
rect 110638 445770 110644 445772
rect 110413 445768 110644 445770
rect 110413 445712 110418 445768
rect 110474 445712 110644 445768
rect 110413 445710 110644 445712
rect 110413 445707 110479 445710
rect 110638 445708 110644 445710
rect 110708 445770 110714 445772
rect 111149 445770 111215 445773
rect 110708 445768 111215 445770
rect 110708 445712 111154 445768
rect 111210 445712 111215 445768
rect 110708 445710 111215 445712
rect 110708 445708 110714 445710
rect 111149 445707 111215 445710
rect 113173 445770 113239 445773
rect 114093 445770 114159 445773
rect 114318 445770 114324 445772
rect 113173 445768 114324 445770
rect 113173 445712 113178 445768
rect 113234 445712 114098 445768
rect 114154 445712 114324 445768
rect 113173 445710 114324 445712
rect 113173 445707 113239 445710
rect 114093 445707 114159 445710
rect 114318 445708 114324 445710
rect 114388 445708 114394 445772
rect 117313 445770 117379 445773
rect 118550 445770 118556 445772
rect 117313 445768 118556 445770
rect 117313 445712 117318 445768
rect 117374 445712 118556 445768
rect 117313 445710 118556 445712
rect 117313 445707 117379 445710
rect 118550 445708 118556 445710
rect 118620 445708 118626 445772
rect 109033 444682 109099 444685
rect 109166 444682 109172 444684
rect 109033 444680 109172 444682
rect 109033 444624 109038 444680
rect 109094 444624 109172 444680
rect 109033 444622 109172 444624
rect 109033 444619 109099 444622
rect 109166 444620 109172 444622
rect 109236 444620 109242 444684
rect 119015 444682 119081 444685
rect 119838 444682 119844 444684
rect 119015 444680 119844 444682
rect 119015 444624 119020 444680
rect 119076 444624 119844 444680
rect 119015 444622 119844 444624
rect 119015 444619 119081 444622
rect 119838 444620 119844 444622
rect 119908 444620 119914 444684
rect 583520 444668 584960 444908
rect 90127 444546 90193 444549
rect 137277 444546 137343 444549
rect 90127 444544 137343 444546
rect 90127 444488 90132 444544
rect 90188 444488 137282 444544
rect 137338 444488 137343 444544
rect 90127 444486 137343 444488
rect 90127 444483 90193 444486
rect 137277 444483 137343 444486
rect 68645 444274 68711 444277
rect 68870 444274 68876 444276
rect 68645 444272 68876 444274
rect 68645 444216 68650 444272
rect 68706 444216 68876 444272
rect 68645 444214 68876 444216
rect 68645 444211 68711 444214
rect 68870 444212 68876 444214
rect 68940 444212 68946 444276
rect 123334 444274 123340 444276
rect 120612 444214 123340 444274
rect 123334 444212 123340 444214
rect 123404 444212 123410 444276
rect 120022 442716 120028 442780
rect 120092 442778 120098 442780
rect 120092 442718 122850 442778
rect 120092 442716 120098 442718
rect 122790 442370 122850 442718
rect 143574 442370 143580 442372
rect 122790 442310 143580 442370
rect 143574 442308 143580 442310
rect 143644 442308 143650 442372
rect 67725 442098 67791 442101
rect 67725 442096 68908 442098
rect 67725 442040 67730 442096
rect 67786 442040 68908 442096
rect 67725 442038 68908 442040
rect 67725 442035 67791 442038
rect 120582 441690 120642 442068
rect 165654 441690 165660 441692
rect 120582 441630 165660 441690
rect 165654 441628 165660 441630
rect 165724 441628 165730 441692
rect 66989 439922 67055 439925
rect 124121 439922 124187 439925
rect 66989 439920 68908 439922
rect 66989 439864 66994 439920
rect 67050 439864 68908 439920
rect 66989 439862 68908 439864
rect 120612 439920 124187 439922
rect 120612 439864 124126 439920
rect 124182 439864 124187 439920
rect 120612 439862 124187 439864
rect 66989 439859 67055 439862
rect 124121 439859 124187 439862
rect 66529 437746 66595 437749
rect 123661 437746 123727 437749
rect 66529 437744 68908 437746
rect 66529 437688 66534 437744
rect 66590 437688 68908 437744
rect 66529 437686 68908 437688
rect 120612 437744 123727 437746
rect 120612 437688 123666 437744
rect 123722 437688 123727 437744
rect 120612 437686 123727 437688
rect 66529 437683 66595 437686
rect 123661 437683 123727 437686
rect -960 436508 480 436748
rect 66805 435298 66871 435301
rect 122782 435298 122788 435300
rect 66805 435296 68908 435298
rect 66805 435240 66810 435296
rect 66866 435240 68908 435296
rect 120428 435268 122788 435298
rect 66805 435238 68908 435240
rect 120398 435238 122788 435268
rect 66805 435235 66871 435238
rect 120398 434756 120458 435238
rect 122782 435236 122788 435238
rect 122852 435236 122858 435300
rect 120390 434692 120396 434756
rect 120460 434692 120466 434756
rect 66437 433122 66503 433125
rect 123109 433122 123175 433125
rect 123845 433122 123911 433125
rect 66437 433120 68908 433122
rect 66437 433064 66442 433120
rect 66498 433064 68908 433120
rect 66437 433062 68908 433064
rect 120612 433120 123911 433122
rect 120612 433064 123114 433120
rect 123170 433064 123850 433120
rect 123906 433064 123911 433120
rect 120612 433062 123911 433064
rect 66437 433059 66503 433062
rect 123109 433059 123175 433062
rect 123845 433059 123911 433062
rect 582373 431626 582439 431629
rect 583520 431626 584960 431716
rect 582373 431624 584960 431626
rect 582373 431568 582378 431624
rect 582434 431568 584960 431624
rect 582373 431566 584960 431568
rect 582373 431563 582439 431566
rect 120206 431428 120212 431492
rect 120276 431428 120282 431492
rect 583520 431476 584960 431566
rect 66805 430946 66871 430949
rect 120214 430946 120274 431428
rect 122741 430946 122807 430949
rect 66805 430944 68908 430946
rect 66805 430888 66810 430944
rect 66866 430888 68908 430944
rect 120214 430944 122807 430946
rect 120214 430916 122746 430944
rect 66805 430886 68908 430888
rect 120244 430888 122746 430916
rect 122802 430888 122807 430944
rect 120244 430886 122807 430888
rect 66805 430883 66871 430886
rect 122741 430883 122807 430886
rect 66805 428498 66871 428501
rect 121637 428498 121703 428501
rect 123109 428498 123175 428501
rect 66805 428496 68908 428498
rect 66805 428440 66810 428496
rect 66866 428440 68908 428496
rect 66805 428438 68908 428440
rect 120612 428496 123175 428498
rect 120612 428440 121642 428496
rect 121698 428440 123114 428496
rect 123170 428440 123175 428496
rect 120612 428438 123175 428440
rect 66805 428435 66871 428438
rect 121637 428435 121703 428438
rect 123109 428435 123175 428438
rect 66805 426322 66871 426325
rect 66805 426320 68908 426322
rect 66805 426264 66810 426320
rect 66866 426264 68908 426320
rect 66805 426262 68908 426264
rect 66805 426259 66871 426262
rect 120582 425642 120642 426292
rect 122598 425642 122604 425644
rect 120582 425582 122604 425642
rect 122598 425580 122604 425582
rect 122668 425642 122674 425644
rect 142153 425642 142219 425645
rect 122668 425640 142219 425642
rect 122668 425584 142158 425640
rect 142214 425584 142219 425640
rect 122668 425582 142219 425584
rect 122668 425580 122674 425582
rect 142153 425579 142219 425582
rect 66805 424146 66871 424149
rect 122925 424146 122991 424149
rect 66805 424144 68908 424146
rect 66805 424088 66810 424144
rect 66866 424088 68908 424144
rect 66805 424086 68908 424088
rect 120612 424144 122991 424146
rect 120612 424088 122930 424144
rect 122986 424088 122991 424144
rect 120612 424086 122991 424088
rect 66805 424083 66871 424086
rect 122925 424083 122991 424086
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 66805 421970 66871 421973
rect 123201 421970 123267 421973
rect 66805 421968 68908 421970
rect 66805 421912 66810 421968
rect 66866 421912 68908 421968
rect 66805 421910 68908 421912
rect 120612 421968 123267 421970
rect 120612 421912 123206 421968
rect 123262 421912 123267 421968
rect 120612 421910 123267 421912
rect 66805 421907 66871 421910
rect 123201 421907 123267 421910
rect 66897 419522 66963 419525
rect 120809 419522 120875 419525
rect 66897 419520 68908 419522
rect 66897 419464 66902 419520
rect 66958 419464 68908 419520
rect 120612 419520 120875 419522
rect 120612 419492 120814 419520
rect 66897 419462 68908 419464
rect 120582 419464 120814 419492
rect 120870 419464 120875 419520
rect 120582 419462 120875 419464
rect 66897 419459 66963 419462
rect 120582 419389 120642 419462
rect 120809 419459 120875 419462
rect 120582 419384 120691 419389
rect 120582 419328 120630 419384
rect 120686 419328 120691 419384
rect 120582 419326 120691 419328
rect 120625 419323 120691 419326
rect 583017 418298 583083 418301
rect 583520 418298 584960 418388
rect 583017 418296 584960 418298
rect 583017 418240 583022 418296
rect 583078 418240 584960 418296
rect 583017 418238 584960 418240
rect 583017 418235 583083 418238
rect 583520 418148 584960 418238
rect 66437 417346 66503 417349
rect 123017 417346 123083 417349
rect 66437 417344 68908 417346
rect 66437 417288 66442 417344
rect 66498 417288 68908 417344
rect 120612 417344 123083 417346
rect 120612 417316 123022 417344
rect 66437 417286 68908 417288
rect 120582 417288 123022 417316
rect 123078 417288 123083 417344
rect 120582 417286 123083 417288
rect 66437 417283 66503 417286
rect 120582 416805 120642 417286
rect 123017 417283 123083 417286
rect 120582 416800 120691 416805
rect 120582 416744 120630 416800
rect 120686 416744 120691 416800
rect 120582 416742 120691 416744
rect 120625 416739 120691 416742
rect 66805 415170 66871 415173
rect 124121 415170 124187 415173
rect 66805 415168 68908 415170
rect 66805 415112 66810 415168
rect 66866 415112 68908 415168
rect 66805 415110 68908 415112
rect 120612 415168 124187 415170
rect 120612 415112 124126 415168
rect 124182 415112 124187 415168
rect 120612 415110 124187 415112
rect 66805 415107 66871 415110
rect 124121 415107 124187 415110
rect 67449 412722 67515 412725
rect 123017 412722 123083 412725
rect 67449 412720 68908 412722
rect 67449 412664 67454 412720
rect 67510 412664 68908 412720
rect 67449 412662 68908 412664
rect 120612 412720 123083 412722
rect 120612 412664 123022 412720
rect 123078 412664 123083 412720
rect 120612 412662 123083 412664
rect 67449 412659 67515 412662
rect 123017 412659 123083 412662
rect 120717 411090 120783 411093
rect 120582 411088 120783 411090
rect 120582 411032 120722 411088
rect 120778 411032 120783 411088
rect 120582 411030 120783 411032
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 66662 410484 66668 410548
rect 66732 410546 66738 410548
rect 67817 410546 67883 410549
rect 120582 410546 120642 411030
rect 120717 411027 120783 411030
rect 121177 410546 121243 410549
rect 66732 410544 68908 410546
rect 66732 410488 67822 410544
rect 67878 410488 68908 410544
rect 120582 410544 121243 410546
rect 120582 410516 121182 410544
rect 66732 410486 68908 410488
rect 120612 410488 121182 410516
rect 121238 410488 121243 410544
rect 120612 410486 121243 410488
rect 66732 410484 66738 410486
rect 67817 410483 67883 410486
rect 121177 410483 121243 410486
rect 68369 408370 68435 408373
rect 124121 408370 124187 408373
rect 68369 408368 69276 408370
rect 68369 408312 68374 408368
rect 68430 408340 69276 408368
rect 120612 408368 124187 408370
rect 68430 408312 69306 408340
rect 68369 408310 69306 408312
rect 120612 408312 124126 408368
rect 124182 408312 124187 408368
rect 120612 408310 124187 408312
rect 68369 408307 68435 408310
rect 69246 408236 69306 408310
rect 124121 408307 124187 408310
rect 69238 408172 69244 408236
rect 69308 408172 69314 408236
rect 66253 406194 66319 406197
rect 124121 406194 124187 406197
rect 66253 406192 68908 406194
rect 66253 406136 66258 406192
rect 66314 406136 68908 406192
rect 66253 406134 68908 406136
rect 120612 406192 124187 406194
rect 120612 406136 124126 406192
rect 124182 406136 124187 406192
rect 120612 406134 124187 406136
rect 66253 406131 66319 406134
rect 124121 406131 124187 406134
rect 583385 404970 583451 404973
rect 583520 404970 584960 405060
rect 583385 404968 584960 404970
rect 583385 404912 583390 404968
rect 583446 404912 584960 404968
rect 583385 404910 584960 404912
rect 583385 404907 583451 404910
rect 583520 404820 584960 404910
rect 66253 403746 66319 403749
rect 121678 403746 121684 403748
rect 66253 403744 68908 403746
rect 66253 403688 66258 403744
rect 66314 403688 68908 403744
rect 66253 403686 68908 403688
rect 120612 403686 121684 403746
rect 66253 403683 66319 403686
rect 121678 403684 121684 403686
rect 121748 403746 121754 403748
rect 124029 403746 124095 403749
rect 121748 403744 124095 403746
rect 121748 403688 124034 403744
rect 124090 403688 124095 403744
rect 121748 403686 124095 403688
rect 121748 403684 121754 403686
rect 124029 403683 124095 403686
rect 133781 401706 133847 401709
rect 140814 401706 140820 401708
rect 133781 401704 140820 401706
rect 133781 401648 133786 401704
rect 133842 401648 140820 401704
rect 133781 401646 140820 401648
rect 133781 401643 133847 401646
rect 140814 401644 140820 401646
rect 140884 401644 140890 401708
rect 66253 401570 66319 401573
rect 124121 401570 124187 401573
rect 66253 401568 68908 401570
rect 66253 401512 66258 401568
rect 66314 401512 68908 401568
rect 66253 401510 68908 401512
rect 120612 401568 124187 401570
rect 120612 401512 124126 401568
rect 124182 401512 124187 401568
rect 120612 401510 124187 401512
rect 66253 401507 66319 401510
rect 124121 401507 124187 401510
rect 66437 399394 66503 399397
rect 123661 399394 123727 399397
rect 66437 399392 68908 399394
rect 66437 399336 66442 399392
rect 66498 399336 68908 399392
rect 66437 399334 68908 399336
rect 120612 399392 123727 399394
rect 120612 399336 123666 399392
rect 123722 399336 123727 399392
rect 120612 399334 123727 399336
rect 66437 399331 66503 399334
rect 123661 399331 123727 399334
rect -960 397490 480 397580
rect 2773 397490 2839 397493
rect -960 397488 2839 397490
rect -960 397432 2778 397488
rect 2834 397432 2839 397488
rect -960 397430 2839 397432
rect -960 397340 480 397430
rect 2773 397427 2839 397430
rect 66989 396946 67055 396949
rect 121545 396946 121611 396949
rect 66989 396944 68908 396946
rect 66989 396888 66994 396944
rect 67050 396888 68908 396944
rect 66989 396886 68908 396888
rect 120612 396944 121611 396946
rect 120612 396888 121550 396944
rect 121606 396888 121611 396944
rect 120612 396886 121611 396888
rect 66989 396883 67055 396886
rect 121545 396883 121611 396886
rect 67541 394770 67607 394773
rect 122925 394770 122991 394773
rect 123661 394770 123727 394773
rect 67541 394768 68908 394770
rect 67541 394712 67546 394768
rect 67602 394712 68908 394768
rect 67541 394710 68908 394712
rect 120612 394768 123727 394770
rect 120612 394712 122930 394768
rect 122986 394712 123666 394768
rect 123722 394712 123727 394768
rect 120612 394710 123727 394712
rect 67541 394707 67607 394710
rect 122925 394707 122991 394710
rect 123661 394707 123727 394710
rect 61929 393276 61995 393277
rect 61878 393274 61884 393276
rect 61838 393214 61884 393274
rect 61948 393272 61995 393276
rect 61990 393216 61995 393272
rect 61878 393212 61884 393214
rect 61948 393212 61995 393216
rect 61929 393211 61995 393212
rect 66805 392594 66871 392597
rect 121453 392594 121519 392597
rect 66805 392592 68908 392594
rect 66805 392536 66810 392592
rect 66866 392536 68908 392592
rect 120060 392592 121519 392594
rect 120060 392564 121458 392592
rect 66805 392534 68908 392536
rect 120030 392536 121458 392564
rect 121514 392536 121519 392592
rect 120030 392534 121519 392536
rect 66805 392531 66871 392534
rect 113030 391988 113036 392052
rect 113100 392050 113106 392052
rect 120030 392050 120090 392534
rect 121453 392531 121519 392534
rect 113100 391990 120090 392050
rect 113100 391988 113106 391990
rect 583520 391628 584960 391868
rect 17217 391234 17283 391237
rect 17217 391232 103530 391234
rect 17217 391176 17222 391232
rect 17278 391176 103530 391232
rect 17217 391174 103530 391176
rect 17217 391171 17283 391174
rect 92606 390900 92612 390964
rect 92676 390962 92682 390964
rect 92749 390962 92815 390965
rect 92676 390960 92815 390962
rect 92676 390904 92754 390960
rect 92810 390904 92815 390960
rect 92676 390902 92815 390904
rect 92676 390900 92682 390902
rect 92749 390899 92815 390902
rect 102593 390962 102659 390965
rect 102726 390962 102732 390964
rect 102593 390960 102732 390962
rect 102593 390904 102598 390960
rect 102654 390904 102732 390960
rect 102593 390902 102732 390904
rect 102593 390899 102659 390902
rect 102726 390900 102732 390902
rect 102796 390900 102802 390964
rect 103470 390962 103530 391174
rect 110413 390962 110479 390965
rect 111149 390962 111215 390965
rect 103470 390960 111215 390962
rect 103470 390904 110418 390960
rect 110474 390904 111154 390960
rect 111210 390904 111215 390960
rect 103470 390902 111215 390904
rect 110413 390899 110479 390902
rect 111149 390899 111215 390902
rect 100661 390556 100727 390557
rect 100661 390552 100708 390556
rect 100772 390554 100778 390556
rect 100661 390496 100666 390552
rect 100661 390492 100708 390496
rect 100772 390494 100818 390554
rect 100772 390492 100778 390494
rect 100661 390491 100727 390492
rect 69606 390356 69612 390420
rect 69676 390418 69682 390420
rect 69933 390418 69999 390421
rect 71865 390420 71931 390421
rect 71814 390418 71820 390420
rect 69676 390416 69999 390418
rect 69676 390360 69938 390416
rect 69994 390360 69999 390416
rect 69676 390358 69999 390360
rect 71774 390358 71820 390418
rect 71884 390416 71931 390420
rect 71926 390360 71931 390416
rect 69676 390356 69682 390358
rect 69933 390355 69999 390358
rect 71814 390356 71820 390358
rect 71884 390356 71931 390360
rect 89662 390356 89668 390420
rect 89732 390418 89738 390420
rect 89805 390418 89871 390421
rect 89732 390416 89871 390418
rect 89732 390360 89810 390416
rect 89866 390360 89871 390416
rect 89732 390358 89871 390360
rect 89732 390356 89738 390358
rect 71865 390355 71931 390356
rect 89805 390355 89871 390358
rect 91134 390356 91140 390420
rect 91204 390418 91210 390420
rect 91277 390418 91343 390421
rect 91204 390416 91343 390418
rect 91204 390360 91282 390416
rect 91338 390360 91343 390416
rect 91204 390358 91343 390360
rect 91204 390356 91210 390358
rect 91277 390355 91343 390358
rect 96838 390356 96844 390420
rect 96908 390418 96914 390420
rect 97349 390418 97415 390421
rect 96908 390416 97415 390418
rect 96908 390360 97354 390416
rect 97410 390360 97415 390416
rect 96908 390358 97415 390360
rect 96908 390356 96914 390358
rect 97349 390355 97415 390358
rect 98126 390356 98132 390420
rect 98196 390418 98202 390420
rect 98821 390418 98887 390421
rect 98196 390416 98887 390418
rect 98196 390360 98826 390416
rect 98882 390360 98887 390416
rect 98196 390358 98887 390360
rect 98196 390356 98202 390358
rect 98821 390355 98887 390358
rect 104934 390356 104940 390420
rect 105004 390418 105010 390420
rect 105077 390418 105143 390421
rect 105004 390416 105143 390418
rect 105004 390360 105082 390416
rect 105138 390360 105143 390416
rect 105004 390358 105143 390360
rect 105004 390356 105010 390358
rect 105077 390355 105143 390358
rect 106406 390356 106412 390420
rect 106476 390418 106482 390420
rect 106549 390418 106615 390421
rect 106476 390416 106615 390418
rect 106476 390360 106554 390416
rect 106610 390360 106615 390416
rect 106476 390358 106615 390360
rect 106476 390356 106482 390358
rect 106549 390355 106615 390358
rect 107694 390356 107700 390420
rect 107764 390418 107770 390420
rect 108021 390418 108087 390421
rect 107764 390416 108087 390418
rect 107764 390360 108026 390416
rect 108082 390360 108087 390416
rect 107764 390358 108087 390360
rect 107764 390356 107770 390358
rect 108021 390355 108087 390358
rect 109350 390356 109356 390420
rect 109420 390418 109426 390420
rect 109493 390418 109559 390421
rect 109420 390416 109559 390418
rect 109420 390360 109498 390416
rect 109554 390360 109559 390416
rect 109420 390358 109559 390360
rect 109420 390356 109426 390358
rect 109493 390355 109559 390358
rect 115933 390420 115999 390421
rect 120257 390420 120323 390421
rect 115933 390416 115980 390420
rect 116044 390418 116050 390420
rect 120206 390418 120212 390420
rect 115933 390360 115938 390416
rect 115933 390356 115980 390360
rect 116044 390358 116090 390418
rect 120166 390358 120212 390418
rect 120276 390416 120323 390420
rect 120318 390360 120323 390416
rect 116044 390356 116050 390358
rect 120206 390356 120212 390358
rect 120276 390356 120323 390360
rect 115933 390355 115999 390356
rect 120257 390355 120323 390356
rect 67817 389874 67883 389877
rect 100109 389874 100175 389877
rect 67817 389872 100175 389874
rect 67817 389816 67822 389872
rect 67878 389816 100114 389872
rect 100170 389816 100175 389872
rect 67817 389814 100175 389816
rect 67817 389811 67883 389814
rect 100109 389811 100175 389814
rect 111006 389404 111012 389468
rect 111076 389466 111082 389468
rect 118693 389466 118759 389469
rect 111076 389464 118759 389466
rect 111076 389408 118698 389464
rect 118754 389408 118759 389464
rect 111076 389406 118759 389408
rect 111076 389404 111082 389406
rect 118693 389403 118759 389406
rect 108297 389330 108363 389333
rect 114093 389330 114159 389333
rect 108297 389328 114159 389330
rect 108297 389272 108302 389328
rect 108358 389272 114098 389328
rect 114154 389272 114159 389328
rect 108297 389270 114159 389272
rect 108297 389267 108363 389270
rect 114093 389267 114159 389270
rect 96470 389132 96476 389196
rect 96540 389194 96546 389196
rect 117773 389194 117839 389197
rect 96540 389192 117839 389194
rect 96540 389136 117778 389192
rect 117834 389136 117839 389192
rect 96540 389134 117839 389136
rect 96540 389132 96546 389134
rect 117773 389131 117839 389134
rect 72049 389058 72115 389061
rect 73061 389058 73127 389061
rect 72049 389056 73127 389058
rect 72049 389000 72054 389056
rect 72110 389000 73066 389056
rect 73122 389000 73127 389056
rect 72049 388998 73127 389000
rect 72049 388995 72115 388998
rect 73061 388995 73127 388998
rect 85481 389058 85547 389061
rect 90357 389058 90423 389061
rect 85481 389056 90423 389058
rect 85481 389000 85486 389056
rect 85542 389000 90362 389056
rect 90418 389000 90423 389056
rect 85481 388998 90423 389000
rect 85481 388995 85547 388998
rect 90357 388995 90423 388998
rect 95182 388996 95188 389060
rect 95252 389058 95258 389060
rect 95877 389058 95943 389061
rect 95252 389056 95943 389058
rect 95252 389000 95882 389056
rect 95938 389000 95943 389056
rect 95252 388998 95943 389000
rect 95252 388996 95258 388998
rect 95877 388995 95943 388998
rect 102593 389058 102659 389061
rect 105537 389058 105603 389061
rect 111793 389060 111859 389061
rect 111742 389058 111748 389060
rect 102593 389056 105603 389058
rect 102593 389000 102598 389056
rect 102654 389000 105542 389056
rect 105598 389000 105603 389056
rect 102593 388998 105603 389000
rect 111666 388998 111748 389058
rect 111812 389058 111859 389060
rect 112621 389058 112687 389061
rect 111812 389056 112687 389058
rect 111854 389000 112626 389056
rect 112682 389000 112687 389056
rect 102593 388995 102659 388998
rect 105537 388995 105603 388998
rect 111742 388996 111748 388998
rect 111812 388998 112687 389000
rect 111812 388996 111859 388998
rect 111793 388995 111859 388996
rect 112621 388995 112687 388998
rect 65977 388922 66043 388925
rect 74533 388922 74599 388925
rect 65977 388920 74599 388922
rect 65977 388864 65982 388920
rect 66038 388864 74538 388920
rect 74594 388864 74599 388920
rect 65977 388862 74599 388864
rect 65977 388859 66043 388862
rect 74533 388859 74599 388862
rect 136633 388786 136699 388789
rect 137134 388786 137140 388788
rect 136633 388784 137140 388786
rect 136633 388728 136638 388784
rect 136694 388728 137140 388784
rect 136633 388726 137140 388728
rect 136633 388723 136699 388726
rect 137134 388724 137140 388726
rect 137204 388724 137210 388788
rect 66161 388378 66227 388381
rect 79961 388378 80027 388381
rect 66161 388376 80027 388378
rect 66161 388320 66166 388376
rect 66222 388320 79966 388376
rect 80022 388320 80027 388376
rect 66161 388318 80027 388320
rect 66161 388315 66227 388318
rect 79961 388315 80027 388318
rect 93761 388378 93827 388381
rect 99966 388378 99972 388380
rect 93761 388376 99972 388378
rect 93761 388320 93766 388376
rect 93822 388320 99972 388376
rect 93761 388318 99972 388320
rect 93761 388315 93827 388318
rect 99966 388316 99972 388318
rect 100036 388378 100042 388380
rect 108297 388378 108363 388381
rect 100036 388376 108363 388378
rect 100036 388320 108302 388376
rect 108358 388320 108363 388376
rect 100036 388318 108363 388320
rect 100036 388316 100042 388318
rect 108297 388315 108363 388318
rect 76557 387154 76623 387157
rect 122598 387154 122604 387156
rect 76557 387152 122604 387154
rect 76557 387096 76562 387152
rect 76618 387096 122604 387152
rect 76557 387094 122604 387096
rect 76557 387091 76623 387094
rect 122598 387092 122604 387094
rect 122668 387092 122674 387156
rect 33777 387018 33843 387021
rect 105629 387018 105695 387021
rect 33777 387016 105695 387018
rect 33777 386960 33782 387016
rect 33838 386960 105634 387016
rect 105690 386960 105695 387016
rect 33777 386958 105695 386960
rect 33777 386955 33843 386958
rect 105629 386955 105695 386958
rect 114318 386276 114324 386340
rect 114388 386338 114394 386340
rect 119337 386338 119403 386341
rect 114388 386336 119403 386338
rect 114388 386280 119342 386336
rect 119398 386280 119403 386336
rect 114388 386278 119403 386280
rect 114388 386276 114394 386278
rect 119337 386275 119403 386278
rect 64597 385658 64663 385661
rect 108297 385658 108363 385661
rect 64597 385656 108363 385658
rect 64597 385600 64602 385656
rect 64658 385600 108302 385656
rect 108358 385600 108363 385656
rect 64597 385598 108363 385600
rect 64597 385595 64663 385598
rect 108297 385595 108363 385598
rect -960 384284 480 384524
rect 84009 383074 84075 383077
rect 109166 383074 109172 383076
rect 84009 383072 109172 383074
rect 84009 383016 84014 383072
rect 84070 383016 109172 383072
rect 84009 383014 109172 383016
rect 84009 383011 84075 383014
rect 109166 383012 109172 383014
rect 109236 383012 109242 383076
rect 7557 382938 7623 382941
rect 95182 382938 95188 382940
rect 7557 382936 95188 382938
rect 7557 382880 7562 382936
rect 7618 382880 95188 382936
rect 7557 382878 95188 382880
rect 7557 382875 7623 382878
rect 95182 382876 95188 382878
rect 95252 382876 95258 382940
rect 68686 378660 68692 378724
rect 68756 378722 68762 378724
rect 122833 378722 122899 378725
rect 68756 378720 122899 378722
rect 68756 378664 122838 378720
rect 122894 378664 122899 378720
rect 68756 378662 122899 378664
rect 68756 378660 68762 378662
rect 122833 378659 122899 378662
rect 582833 378450 582899 378453
rect 583520 378450 584960 378540
rect 582833 378448 584960 378450
rect 582833 378392 582838 378448
rect 582894 378392 584960 378448
rect 582833 378390 584960 378392
rect 582833 378387 582899 378390
rect 583520 378300 584960 378390
rect 68870 377300 68876 377364
rect 68940 377362 68946 377364
rect 145557 377362 145623 377365
rect 68940 377360 145623 377362
rect 68940 377304 145562 377360
rect 145618 377304 145623 377360
rect 68940 377302 145623 377304
rect 68940 377300 68946 377302
rect 145557 377299 145623 377302
rect 84101 374642 84167 374645
rect 119429 374642 119495 374645
rect 84101 374640 119495 374642
rect 84101 374584 84106 374640
rect 84162 374584 119434 374640
rect 119490 374584 119495 374640
rect 84101 374582 119495 374584
rect 84101 374579 84167 374582
rect 119429 374579 119495 374582
rect -960 371378 480 371468
rect 3141 371378 3207 371381
rect -960 371376 3207 371378
rect -960 371320 3146 371376
rect 3202 371320 3207 371376
rect -960 371318 3207 371320
rect -960 371228 480 371318
rect 3141 371315 3207 371318
rect 90214 371316 90220 371380
rect 90284 371378 90290 371380
rect 91001 371378 91067 371381
rect 185577 371378 185643 371381
rect 90284 371376 185643 371378
rect 90284 371320 91006 371376
rect 91062 371320 185582 371376
rect 185638 371320 185643 371376
rect 90284 371318 185643 371320
rect 90284 371316 90290 371318
rect 91001 371315 91067 371318
rect 185577 371315 185643 371318
rect 94497 369882 94563 369885
rect 94998 369882 95004 369884
rect 94497 369880 95004 369882
rect 94497 369824 94502 369880
rect 94558 369824 95004 369880
rect 94497 369822 95004 369824
rect 94497 369819 94563 369822
rect 94998 369820 95004 369822
rect 95068 369882 95074 369884
rect 195329 369882 195395 369885
rect 95068 369880 195395 369882
rect 95068 369824 195334 369880
rect 195390 369824 195395 369880
rect 95068 369822 195395 369824
rect 95068 369820 95074 369822
rect 195329 369819 195395 369822
rect 81341 369066 81407 369069
rect 96654 369066 96660 369068
rect 81341 369064 96660 369066
rect 81341 369008 81346 369064
rect 81402 369008 96660 369064
rect 81341 369006 96660 369008
rect 81341 369003 81407 369006
rect 96654 369004 96660 369006
rect 96724 369004 96730 369068
rect 137921 368522 137987 368525
rect 327073 368522 327139 368525
rect 137921 368520 327139 368522
rect 137921 368464 137926 368520
rect 137982 368464 327078 368520
rect 327134 368464 327139 368520
rect 137921 368462 327139 368464
rect 137921 368459 137987 368462
rect 327073 368459 327139 368462
rect 98637 368386 98703 368389
rect 99046 368386 99052 368388
rect 98637 368384 99052 368386
rect 98637 368328 98642 368384
rect 98698 368328 99052 368384
rect 98637 368326 99052 368328
rect 98637 368323 98703 368326
rect 99046 368324 99052 368326
rect 99116 368324 99122 368388
rect 79961 367706 80027 367709
rect 110638 367706 110644 367708
rect 79961 367704 110644 367706
rect 79961 367648 79966 367704
rect 80022 367648 110644 367704
rect 79961 367646 110644 367648
rect 79961 367643 80027 367646
rect 110638 367644 110644 367646
rect 110708 367644 110714 367708
rect 98637 367162 98703 367165
rect 221457 367162 221523 367165
rect 98637 367160 221523 367162
rect 98637 367104 98642 367160
rect 98698 367104 221462 367160
rect 221518 367104 221523 367160
rect 98637 367102 221523 367104
rect 98637 367099 98703 367102
rect 221457 367099 221523 367102
rect 76649 366346 76715 366349
rect 138054 366346 138060 366348
rect 76649 366344 138060 366346
rect 76649 366288 76654 366344
rect 76710 366288 138060 366344
rect 76649 366286 138060 366288
rect 76649 366283 76715 366286
rect 138054 366284 138060 366286
rect 138124 366284 138130 366348
rect 130469 365802 130535 365805
rect 207974 365802 207980 365804
rect 130469 365800 207980 365802
rect 130469 365744 130474 365800
rect 130530 365744 207980 365800
rect 130469 365742 207980 365744
rect 130469 365739 130535 365742
rect 207974 365740 207980 365742
rect 208044 365740 208050 365804
rect 117313 365666 117379 365669
rect 118550 365666 118556 365668
rect 117313 365664 118556 365666
rect 117313 365608 117318 365664
rect 117374 365608 118556 365664
rect 117313 365606 118556 365608
rect 117313 365603 117379 365606
rect 118550 365604 118556 365606
rect 118620 365604 118626 365668
rect 582373 365122 582439 365125
rect 583520 365122 584960 365212
rect 582373 365120 584960 365122
rect 582373 365064 582378 365120
rect 582434 365064 584960 365120
rect 582373 365062 584960 365064
rect 582373 365059 582439 365062
rect 583520 364972 584960 365062
rect 121361 364578 121427 364581
rect 184054 364578 184060 364580
rect 121361 364576 184060 364578
rect 121361 364520 121366 364576
rect 121422 364520 184060 364576
rect 121361 364518 184060 364520
rect 121361 364515 121427 364518
rect 184054 364516 184060 364518
rect 184124 364516 184130 364580
rect 117313 364442 117379 364445
rect 262213 364442 262279 364445
rect 117313 364440 262279 364442
rect 117313 364384 117318 364440
rect 117374 364384 262218 364440
rect 262274 364384 262279 364440
rect 117313 364382 262279 364384
rect 117313 364379 117379 364382
rect 262213 364379 262279 364382
rect 128261 363626 128327 363629
rect 158805 363626 158871 363629
rect 128261 363624 158871 363626
rect 128261 363568 128266 363624
rect 128322 363568 158810 363624
rect 158866 363568 158871 363624
rect 128261 363566 158871 363568
rect 128261 363563 128327 363566
rect 158805 363563 158871 363566
rect 107837 363082 107903 363085
rect 215937 363082 216003 363085
rect 107837 363080 216003 363082
rect 107837 363024 107842 363080
rect 107898 363024 215942 363080
rect 215998 363024 216003 363080
rect 107837 363022 216003 363024
rect 107837 363019 107903 363022
rect 215937 363019 216003 363022
rect 63217 362266 63283 362269
rect 126973 362266 127039 362269
rect 63217 362264 132510 362266
rect 63217 362208 63222 362264
rect 63278 362208 126978 362264
rect 127034 362208 132510 362264
rect 63217 362206 132510 362208
rect 63217 362203 63283 362206
rect 126973 362203 127039 362206
rect 132450 361722 132510 362206
rect 233734 361722 233740 361724
rect 132450 361662 233740 361722
rect 233734 361660 233740 361662
rect 233804 361660 233810 361724
rect 66069 360906 66135 360909
rect 156454 360906 156460 360908
rect 66069 360904 156460 360906
rect 66069 360848 66074 360904
rect 66130 360848 156460 360904
rect 66069 360846 156460 360848
rect 66069 360843 66135 360846
rect 156454 360844 156460 360846
rect 156524 360844 156530 360908
rect 120022 360300 120028 360364
rect 120092 360362 120098 360364
rect 120717 360362 120783 360365
rect 248454 360362 248460 360364
rect 120092 360360 248460 360362
rect 120092 360304 120722 360360
rect 120778 360304 248460 360360
rect 120092 360302 248460 360304
rect 120092 360300 120098 360302
rect 120717 360299 120783 360302
rect 248454 360300 248460 360302
rect 248524 360300 248530 360364
rect 102041 360226 102107 360229
rect 322974 360226 322980 360228
rect 102041 360224 322980 360226
rect 102041 360168 102046 360224
rect 102102 360168 322980 360224
rect 102041 360166 322980 360168
rect 102041 360163 102107 360166
rect 322974 360164 322980 360166
rect 323044 360164 323050 360228
rect 89621 358866 89687 358869
rect 317454 358866 317460 358868
rect 89621 358864 317460 358866
rect 89621 358808 89626 358864
rect 89682 358808 317460 358864
rect 89621 358806 317460 358808
rect 89621 358803 89687 358806
rect 317454 358804 317460 358806
rect 317524 358804 317530 358868
rect -960 358458 480 358548
rect 3417 358458 3483 358461
rect -960 358456 3483 358458
rect -960 358400 3422 358456
rect 3478 358400 3483 358456
rect -960 358398 3483 358400
rect -960 358308 480 358398
rect 3417 358395 3483 358398
rect 58985 358050 59051 358053
rect 160185 358050 160251 358053
rect 58985 358048 160251 358050
rect 58985 357992 58990 358048
rect 59046 357992 160190 358048
rect 160246 357992 160251 358048
rect 58985 357990 160251 357992
rect 58985 357987 59051 357990
rect 160185 357987 160251 357990
rect 119429 357506 119495 357509
rect 233877 357506 233943 357509
rect 119429 357504 233943 357506
rect 119429 357448 119434 357504
rect 119490 357448 233882 357504
rect 233938 357448 233943 357504
rect 119429 357446 233943 357448
rect 119429 357443 119495 357446
rect 233877 357443 233943 357446
rect 125685 357370 125751 357373
rect 126881 357370 126947 357373
rect 125685 357368 126947 357370
rect 125685 357312 125690 357368
rect 125746 357312 126886 357368
rect 126942 357312 126947 357368
rect 125685 357310 126947 357312
rect 125685 357307 125751 357310
rect 126881 357307 126947 357310
rect 112437 356690 112503 356693
rect 151169 356690 151235 356693
rect 155861 356690 155927 356693
rect 112437 356688 155927 356690
rect 112437 356632 112442 356688
rect 112498 356632 151174 356688
rect 151230 356632 155866 356688
rect 155922 356632 155927 356688
rect 112437 356630 155927 356632
rect 112437 356627 112503 356630
rect 151169 356627 151235 356630
rect 155861 356627 155927 356630
rect 125685 356146 125751 356149
rect 252553 356146 252619 356149
rect 125685 356144 252619 356146
rect 125685 356088 125690 356144
rect 125746 356088 252558 356144
rect 252614 356088 252619 356144
rect 125685 356086 252619 356088
rect 125685 356083 125751 356086
rect 252553 356083 252619 356086
rect 135897 355602 135963 355605
rect 151854 355602 151860 355604
rect 135897 355600 151860 355602
rect 135897 355544 135902 355600
rect 135958 355544 151860 355600
rect 135897 355542 151860 355544
rect 135897 355539 135963 355542
rect 151854 355540 151860 355542
rect 151924 355540 151930 355604
rect 77937 355466 78003 355469
rect 136030 355466 136036 355468
rect 77937 355464 136036 355466
rect 77937 355408 77942 355464
rect 77998 355408 136036 355464
rect 77937 355406 136036 355408
rect 77937 355403 78003 355406
rect 136030 355404 136036 355406
rect 136100 355404 136106 355468
rect 152457 355466 152523 355469
rect 164233 355466 164299 355469
rect 152457 355464 164299 355466
rect 152457 355408 152462 355464
rect 152518 355408 164238 355464
rect 164294 355408 164299 355464
rect 152457 355406 164299 355408
rect 152457 355403 152523 355406
rect 164233 355403 164299 355406
rect 116577 355330 116643 355333
rect 131113 355330 131179 355333
rect 255313 355330 255379 355333
rect 116577 355328 255379 355330
rect 116577 355272 116582 355328
rect 116638 355272 131118 355328
rect 131174 355272 255318 355328
rect 255374 355272 255379 355328
rect 116577 355270 255379 355272
rect 116577 355267 116643 355270
rect 131113 355267 131179 355270
rect 255313 355267 255379 355270
rect 144913 353834 144979 353837
rect 145557 353834 145623 353837
rect 144913 353832 151830 353834
rect 144913 353776 144918 353832
rect 144974 353776 145562 353832
rect 145618 353776 151830 353832
rect 144913 353774 151830 353776
rect 144913 353771 144979 353774
rect 145557 353771 145623 353774
rect 112437 353698 112503 353701
rect 113030 353698 113036 353700
rect 112437 353696 113036 353698
rect 112437 353640 112442 353696
rect 112498 353640 113036 353696
rect 112437 353638 113036 353640
rect 112437 353635 112503 353638
rect 113030 353636 113036 353638
rect 113100 353698 113106 353700
rect 144821 353698 144887 353701
rect 113100 353696 144887 353698
rect 113100 353640 144826 353696
rect 144882 353640 144887 353696
rect 113100 353638 144887 353640
rect 151770 353698 151830 353774
rect 206277 353698 206343 353701
rect 151770 353696 206343 353698
rect 151770 353640 206282 353696
rect 206338 353640 206343 353696
rect 151770 353638 206343 353640
rect 113100 353636 113106 353638
rect 144821 353635 144887 353638
rect 206277 353635 206343 353638
rect 83457 353562 83523 353565
rect 84009 353562 84075 353565
rect 178677 353562 178743 353565
rect 83457 353560 178743 353562
rect 83457 353504 83462 353560
rect 83518 353504 84014 353560
rect 84070 353504 178682 353560
rect 178738 353504 178743 353560
rect 83457 353502 178743 353504
rect 83457 353499 83523 353502
rect 84009 353499 84075 353502
rect 178677 353499 178743 353502
rect 121453 353426 121519 353429
rect 122741 353426 122807 353429
rect 234613 353426 234679 353429
rect 121453 353424 234679 353426
rect 121453 353368 121458 353424
rect 121514 353368 122746 353424
rect 122802 353368 234618 353424
rect 234674 353368 234679 353424
rect 121453 353366 234679 353368
rect 121453 353363 121519 353366
rect 122741 353363 122807 353366
rect 234613 353363 234679 353366
rect 69790 352548 69796 352612
rect 69860 352610 69866 352612
rect 85757 352610 85823 352613
rect 69860 352608 85823 352610
rect 69860 352552 85762 352608
rect 85818 352552 85823 352608
rect 69860 352550 85823 352552
rect 69860 352548 69866 352550
rect 85757 352547 85823 352550
rect 88977 352610 89043 352613
rect 129825 352610 129891 352613
rect 88977 352608 129891 352610
rect 88977 352552 88982 352608
rect 89038 352552 129830 352608
rect 129886 352552 129891 352608
rect 88977 352550 129891 352552
rect 88977 352547 89043 352550
rect 129825 352547 129891 352550
rect 144821 352610 144887 352613
rect 204897 352610 204963 352613
rect 144821 352608 204963 352610
rect 144821 352552 144826 352608
rect 144882 352552 204902 352608
rect 204958 352552 204963 352608
rect 144821 352550 204963 352552
rect 144821 352547 144887 352550
rect 204897 352547 204963 352550
rect 106917 352066 106983 352069
rect 181437 352066 181503 352069
rect 106917 352064 181503 352066
rect 106917 352008 106922 352064
rect 106978 352008 181442 352064
rect 181498 352008 181503 352064
rect 106917 352006 181503 352008
rect 106917 352003 106983 352006
rect 181437 352003 181503 352006
rect 129825 351930 129891 351933
rect 231894 351930 231900 351932
rect 129825 351928 231900 351930
rect 129825 351872 129830 351928
rect 129886 351872 231900 351928
rect 129825 351870 231900 351872
rect 129825 351867 129891 351870
rect 231894 351868 231900 351870
rect 231964 351868 231970 351932
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 70158 351052 70164 351116
rect 70228 351114 70234 351116
rect 85573 351114 85639 351117
rect 70228 351112 85639 351114
rect 70228 351056 85578 351112
rect 85634 351056 85639 351112
rect 70228 351054 85639 351056
rect 70228 351052 70234 351054
rect 85573 351051 85639 351054
rect 64781 350842 64847 350845
rect 229686 350842 229692 350844
rect 64781 350840 229692 350842
rect 64781 350784 64786 350840
rect 64842 350784 229692 350840
rect 64781 350782 229692 350784
rect 64781 350779 64847 350782
rect 229686 350780 229692 350782
rect 229756 350780 229762 350844
rect 93209 350706 93275 350709
rect 93761 350706 93827 350709
rect 259453 350706 259519 350709
rect 93209 350704 259519 350706
rect 93209 350648 93214 350704
rect 93270 350648 93766 350704
rect 93822 350648 259458 350704
rect 259514 350648 259519 350704
rect 93209 350646 259519 350648
rect 93209 350643 93275 350646
rect 93761 350643 93827 350646
rect 259453 350643 259519 350646
rect 136541 350570 136607 350573
rect 340873 350570 340939 350573
rect 136541 350568 340939 350570
rect 136541 350512 136546 350568
rect 136602 350512 340878 350568
rect 340934 350512 340939 350568
rect 136541 350510 340939 350512
rect 136541 350507 136607 350510
rect 340873 350507 340939 350510
rect 130377 349890 130443 349893
rect 139710 349890 139716 349892
rect 130377 349888 139716 349890
rect 130377 349832 130382 349888
rect 130438 349832 139716 349888
rect 130377 349830 139716 349832
rect 130377 349827 130443 349830
rect 139710 349828 139716 349830
rect 139780 349828 139786 349892
rect 67766 349692 67772 349756
rect 67836 349754 67842 349756
rect 115933 349754 115999 349757
rect 67836 349752 115999 349754
rect 67836 349696 115938 349752
rect 115994 349696 115999 349752
rect 67836 349694 115999 349696
rect 67836 349692 67842 349694
rect 115933 349691 115999 349694
rect 134517 349754 134583 349757
rect 156137 349754 156203 349757
rect 134517 349752 156203 349754
rect 134517 349696 134522 349752
rect 134578 349696 156142 349752
rect 156198 349696 156203 349752
rect 134517 349694 156203 349696
rect 134517 349691 134583 349694
rect 156137 349691 156203 349694
rect 113081 349210 113147 349213
rect 188286 349210 188292 349212
rect 113081 349208 188292 349210
rect 113081 349152 113086 349208
rect 113142 349152 188292 349208
rect 113081 349150 188292 349152
rect 113081 349147 113147 349150
rect 188286 349148 188292 349150
rect 188356 349148 188362 349212
rect 128445 348394 128511 348397
rect 210417 348394 210483 348397
rect 128445 348392 210483 348394
rect 128445 348336 128450 348392
rect 128506 348336 210422 348392
rect 210478 348336 210483 348392
rect 128445 348334 210483 348336
rect 128445 348331 128511 348334
rect 210417 348331 210483 348334
rect 70301 347986 70367 347989
rect 187049 347986 187115 347989
rect 70301 347984 187115 347986
rect 70301 347928 70306 347984
rect 70362 347928 187054 347984
rect 187110 347928 187115 347984
rect 70301 347926 187115 347928
rect 70301 347923 70367 347926
rect 187049 347923 187115 347926
rect 110413 347850 110479 347853
rect 111701 347850 111767 347853
rect 251357 347850 251423 347853
rect 110413 347848 251423 347850
rect 110413 347792 110418 347848
rect 110474 347792 111706 347848
rect 111762 347792 251362 347848
rect 251418 347792 251423 347848
rect 110413 347790 251423 347792
rect 110413 347787 110479 347790
rect 111701 347787 111767 347790
rect 251357 347787 251423 347790
rect 105537 347034 105603 347037
rect 153837 347034 153903 347037
rect 105537 347032 153903 347034
rect 105537 346976 105542 347032
rect 105598 346976 153842 347032
rect 153898 346976 153903 347032
rect 105537 346974 153903 346976
rect 105537 346971 105603 346974
rect 153837 346971 153903 346974
rect 115289 346626 115355 346629
rect 180057 346626 180123 346629
rect 115289 346624 180123 346626
rect 115289 346568 115294 346624
rect 115350 346568 180062 346624
rect 180118 346568 180123 346624
rect 115289 346566 180123 346568
rect 115289 346563 115355 346566
rect 180057 346563 180123 346566
rect 101397 346490 101463 346493
rect 277158 346490 277164 346492
rect 101397 346488 277164 346490
rect 101397 346432 101402 346488
rect 101458 346432 277164 346488
rect 101397 346430 277164 346432
rect 101397 346427 101463 346430
rect 277158 346428 277164 346430
rect 277228 346428 277234 346492
rect 124857 345674 124923 345677
rect 155953 345674 156019 345677
rect 124857 345672 156019 345674
rect 124857 345616 124862 345672
rect 124918 345616 155958 345672
rect 156014 345616 156019 345672
rect 124857 345614 156019 345616
rect 124857 345611 124923 345614
rect 155953 345611 156019 345614
rect 203006 345612 203012 345676
rect 203076 345674 203082 345676
rect 582373 345674 582439 345677
rect 203076 345672 582439 345674
rect 203076 345616 582378 345672
rect 582434 345616 582439 345672
rect 203076 345614 582439 345616
rect 203076 345612 203082 345614
rect 582373 345611 582439 345614
rect -960 345402 480 345492
rect 3141 345402 3207 345405
rect -960 345400 3207 345402
rect -960 345344 3146 345400
rect 3202 345344 3207 345400
rect -960 345342 3207 345344
rect -960 345252 480 345342
rect 3141 345339 3207 345342
rect 133086 345204 133092 345268
rect 133156 345266 133162 345268
rect 195237 345266 195303 345269
rect 133156 345264 195303 345266
rect 133156 345208 195242 345264
rect 195298 345208 195303 345264
rect 133156 345206 195303 345208
rect 133156 345204 133162 345206
rect 195237 345203 195303 345206
rect 85757 345130 85823 345133
rect 203006 345130 203012 345132
rect 85757 345128 203012 345130
rect 85757 345072 85762 345128
rect 85818 345072 203012 345128
rect 85757 345070 203012 345072
rect 85757 345067 85823 345070
rect 203006 345068 203012 345070
rect 203076 345068 203082 345132
rect 114461 343906 114527 343909
rect 175917 343906 175983 343909
rect 114461 343904 175983 343906
rect 114461 343848 114466 343904
rect 114522 343848 175922 343904
rect 175978 343848 175983 343904
rect 114461 343846 175983 343848
rect 114461 343843 114527 343846
rect 175917 343843 175983 343846
rect 111701 343770 111767 343773
rect 338113 343770 338179 343773
rect 111701 343768 338179 343770
rect 111701 343712 111706 343768
rect 111762 343712 338118 343768
rect 338174 343712 338179 343768
rect 111701 343710 338179 343712
rect 111701 343707 111767 343710
rect 338113 343707 338179 343710
rect 106181 342546 106247 342549
rect 226425 342546 226491 342549
rect 106181 342544 226491 342546
rect 106181 342488 106186 342544
rect 106242 342488 226430 342544
rect 226486 342488 226491 342544
rect 106181 342486 226491 342488
rect 106181 342483 106247 342486
rect 226425 342483 226491 342486
rect 77201 342410 77267 342413
rect 204253 342410 204319 342413
rect 77201 342408 204319 342410
rect 77201 342352 77206 342408
rect 77262 342352 204258 342408
rect 204314 342352 204319 342408
rect 77201 342350 204319 342352
rect 77201 342347 77267 342350
rect 204253 342347 204319 342350
rect 102777 342274 102843 342277
rect 240726 342274 240732 342276
rect 102777 342272 240732 342274
rect 102777 342216 102782 342272
rect 102838 342216 240732 342272
rect 102777 342214 240732 342216
rect 102777 342211 102843 342214
rect 240726 342212 240732 342214
rect 240796 342212 240802 342276
rect 74993 341458 75059 341461
rect 100753 341458 100819 341461
rect 74993 341456 100819 341458
rect 74993 341400 74998 341456
rect 75054 341400 100758 341456
rect 100814 341400 100819 341456
rect 74993 341398 100819 341400
rect 74993 341395 75059 341398
rect 100753 341395 100819 341398
rect 144821 341186 144887 341189
rect 155166 341186 155172 341188
rect 144821 341184 155172 341186
rect 144821 341128 144826 341184
rect 144882 341128 155172 341184
rect 144821 341126 155172 341128
rect 144821 341123 144887 341126
rect 155166 341124 155172 341126
rect 155236 341124 155242 341188
rect 95141 341050 95207 341053
rect 171777 341050 171843 341053
rect 95141 341048 171843 341050
rect 95141 340992 95146 341048
rect 95202 340992 171782 341048
rect 171838 340992 171843 341048
rect 95141 340990 171843 340992
rect 95141 340987 95207 340990
rect 171777 340987 171843 340990
rect 118601 340914 118667 340917
rect 146201 340914 146267 340917
rect 118601 340912 146267 340914
rect 118601 340856 118606 340912
rect 118662 340856 146206 340912
rect 146262 340856 146267 340912
rect 118601 340854 146267 340856
rect 118601 340851 118667 340854
rect 146201 340851 146267 340854
rect 150341 340914 150407 340917
rect 244222 340914 244228 340916
rect 150341 340912 244228 340914
rect 150341 340856 150346 340912
rect 150402 340856 244228 340912
rect 150341 340854 244228 340856
rect 150341 340851 150407 340854
rect 244222 340852 244228 340854
rect 244292 340852 244298 340916
rect 97901 339826 97967 339829
rect 174629 339826 174695 339829
rect 97901 339824 174695 339826
rect 97901 339768 97906 339824
rect 97962 339768 174634 339824
rect 174690 339768 174695 339824
rect 97901 339766 174695 339768
rect 97901 339763 97967 339766
rect 174629 339763 174695 339766
rect 111793 339690 111859 339693
rect 212574 339690 212580 339692
rect 111793 339688 212580 339690
rect 111793 339632 111798 339688
rect 111854 339632 212580 339688
rect 111793 339630 212580 339632
rect 111793 339627 111859 339630
rect 212574 339628 212580 339630
rect 212644 339628 212650 339692
rect 80697 339554 80763 339557
rect 230974 339554 230980 339556
rect 80697 339552 230980 339554
rect 80697 339496 80702 339552
rect 80758 339496 230980 339552
rect 80697 339494 230980 339496
rect 80697 339491 80763 339494
rect 230974 339492 230980 339494
rect 231044 339492 231050 339556
rect 67357 338466 67423 338469
rect 182817 338466 182883 338469
rect 67357 338464 182883 338466
rect 67357 338408 67362 338464
rect 67418 338408 182822 338464
rect 182878 338408 182883 338464
rect 583520 338452 584960 338692
rect 67357 338406 182883 338408
rect 67357 338403 67423 338406
rect 182817 338403 182883 338406
rect 89437 338330 89503 338333
rect 220077 338330 220143 338333
rect 89437 338328 220143 338330
rect 89437 338272 89442 338328
rect 89498 338272 220082 338328
rect 220138 338272 220143 338328
rect 89437 338270 220143 338272
rect 89437 338267 89503 338270
rect 220077 338267 220143 338270
rect 125501 338194 125567 338197
rect 339493 338194 339559 338197
rect 125501 338192 339559 338194
rect 125501 338136 125506 338192
rect 125562 338136 339498 338192
rect 339554 338136 339559 338192
rect 125501 338134 339559 338136
rect 125501 338131 125567 338134
rect 339493 338131 339559 338134
rect 64597 337378 64663 337381
rect 133137 337378 133203 337381
rect 64597 337376 133203 337378
rect 64597 337320 64602 337376
rect 64658 337320 133142 337376
rect 133198 337320 133203 337376
rect 64597 337318 133203 337320
rect 64597 337315 64663 337318
rect 133137 337315 133203 337318
rect 139393 337106 139459 337109
rect 158069 337106 158135 337109
rect 139393 337104 158135 337106
rect 139393 337048 139398 337104
rect 139454 337048 158074 337104
rect 158130 337048 158135 337104
rect 139393 337046 158135 337048
rect 139393 337043 139459 337046
rect 158069 337043 158135 337046
rect 132585 336970 132651 336973
rect 218697 336970 218763 336973
rect 132585 336968 218763 336970
rect 132585 336912 132590 336968
rect 132646 336912 218702 336968
rect 218758 336912 218763 336968
rect 132585 336910 218763 336912
rect 132585 336907 132651 336910
rect 218697 336907 218763 336910
rect 87137 336834 87203 336837
rect 215385 336834 215451 336837
rect 87137 336832 215451 336834
rect 87137 336776 87142 336832
rect 87198 336776 215390 336832
rect 215446 336776 215451 336832
rect 87137 336774 215451 336776
rect 87137 336771 87203 336774
rect 215385 336771 215451 336774
rect 66662 335956 66668 336020
rect 66732 336018 66738 336020
rect 112437 336018 112503 336021
rect 66732 336016 112503 336018
rect 66732 335960 112442 336016
rect 112498 335960 112503 336016
rect 66732 335958 112503 335960
rect 66732 335956 66738 335958
rect 112437 335955 112503 335958
rect 145373 336018 145439 336021
rect 174537 336018 174603 336021
rect 145373 336016 174603 336018
rect 145373 335960 145378 336016
rect 145434 335960 174542 336016
rect 174598 335960 174603 336016
rect 145373 335958 174603 335960
rect 145373 335955 145439 335958
rect 174537 335955 174603 335958
rect 64689 335610 64755 335613
rect 153929 335610 153995 335613
rect 64689 335608 153995 335610
rect 64689 335552 64694 335608
rect 64750 335552 153934 335608
rect 153990 335552 153995 335608
rect 64689 335550 153995 335552
rect 64689 335547 64755 335550
rect 153929 335547 153995 335550
rect 107745 335474 107811 335477
rect 228449 335474 228515 335477
rect 107745 335472 228515 335474
rect 107745 335416 107750 335472
rect 107806 335416 228454 335472
rect 228510 335416 228515 335472
rect 107745 335414 228515 335416
rect 107745 335411 107811 335414
rect 228449 335411 228515 335414
rect 92749 334386 92815 334389
rect 221549 334386 221615 334389
rect 92749 334384 221615 334386
rect 92749 334328 92754 334384
rect 92810 334328 221554 334384
rect 221610 334328 221615 334384
rect 92749 334326 221615 334328
rect 92749 334323 92815 334326
rect 221549 334323 221615 334326
rect 72969 334250 73035 334253
rect 209037 334250 209103 334253
rect 72969 334248 209103 334250
rect 72969 334192 72974 334248
rect 73030 334192 209042 334248
rect 209098 334192 209103 334248
rect 72969 334190 209103 334192
rect 72969 334187 73035 334190
rect 209037 334187 209103 334190
rect 108757 334114 108823 334117
rect 582373 334114 582439 334117
rect 108757 334112 582439 334114
rect 108757 334056 108762 334112
rect 108818 334056 582378 334112
rect 582434 334056 582439 334112
rect 108757 334054 582439 334056
rect 108757 334051 108823 334054
rect 582373 334051 582439 334054
rect 86309 333298 86375 333301
rect 98637 333298 98703 333301
rect 86309 333296 98703 333298
rect 86309 333240 86314 333296
rect 86370 333240 98642 333296
rect 98698 333240 98703 333296
rect 86309 333238 98703 333240
rect 86309 333235 86375 333238
rect 98637 333235 98703 333238
rect 143441 332890 143507 332893
rect 163773 332890 163839 332893
rect 143441 332888 163839 332890
rect 143441 332832 143446 332888
rect 143502 332832 163778 332888
rect 163834 332832 163839 332888
rect 143441 332830 163839 332832
rect 143441 332827 143507 332830
rect 163773 332827 163839 332830
rect 98545 332754 98611 332757
rect 226977 332754 227043 332757
rect 98545 332752 227043 332754
rect 98545 332696 98550 332752
rect 98606 332696 226982 332752
rect 227038 332696 227043 332752
rect 98545 332694 227043 332696
rect 98545 332691 98611 332694
rect 226977 332691 227043 332694
rect 70669 332618 70735 332621
rect 209129 332618 209195 332621
rect 70669 332616 209195 332618
rect 70669 332560 70674 332616
rect 70730 332560 209134 332616
rect 209190 332560 209195 332616
rect 70669 332558 209195 332560
rect 70669 332555 70735 332558
rect 209129 332555 209195 332558
rect -960 332196 480 332436
rect 132033 331530 132099 331533
rect 169109 331530 169175 331533
rect 132033 331528 169175 331530
rect 132033 331472 132038 331528
rect 132094 331472 169114 331528
rect 169170 331472 169175 331528
rect 132033 331470 169175 331472
rect 132033 331467 132099 331470
rect 169109 331467 169175 331470
rect 90817 331394 90883 331397
rect 211153 331394 211219 331397
rect 90817 331392 211219 331394
rect 90817 331336 90822 331392
rect 90878 331336 211158 331392
rect 211214 331336 211219 331392
rect 90817 331334 211219 331336
rect 90817 331331 90883 331334
rect 211153 331331 211219 331334
rect 69381 331258 69447 331261
rect 207749 331258 207815 331261
rect 69381 331256 207815 331258
rect 69381 331200 69386 331256
rect 69442 331200 207754 331256
rect 207810 331200 207815 331256
rect 69381 331198 207815 331200
rect 69381 331195 69447 331198
rect 207749 331195 207815 331198
rect 109953 331122 110019 331125
rect 115289 331122 115355 331125
rect 109953 331120 115355 331122
rect 109953 331064 109958 331120
rect 110014 331064 115294 331120
rect 115350 331064 115355 331120
rect 109953 331062 115355 331064
rect 109953 331059 110019 331062
rect 115289 331059 115355 331062
rect 84101 330578 84167 330581
rect 84694 330578 84700 330580
rect 84101 330576 84700 330578
rect 84101 330520 84106 330576
rect 84162 330520 84700 330576
rect 84101 330518 84700 330520
rect 84101 330515 84167 330518
rect 84694 330516 84700 330518
rect 84764 330516 84770 330580
rect 99281 330442 99347 330445
rect 106917 330442 106983 330445
rect 99281 330440 106983 330442
rect 99281 330384 99286 330440
rect 99342 330384 106922 330440
rect 106978 330384 106983 330440
rect 99281 330382 106983 330384
rect 99281 330379 99347 330382
rect 106917 330379 106983 330382
rect 182817 330442 182883 330445
rect 230381 330442 230447 330445
rect 182817 330440 230447 330442
rect 182817 330384 182822 330440
rect 182878 330384 230386 330440
rect 230442 330384 230447 330440
rect 182817 330382 230447 330384
rect 182817 330379 182883 330382
rect 230381 330379 230447 330382
rect 134149 330306 134215 330309
rect 196566 330306 196572 330308
rect 134149 330304 196572 330306
rect 134149 330248 134154 330304
rect 134210 330248 196572 330304
rect 134149 330246 196572 330248
rect 134149 330243 134215 330246
rect 196566 330244 196572 330246
rect 196636 330244 196642 330308
rect 132677 330170 132743 330173
rect 154062 330170 154068 330172
rect 132677 330168 154068 330170
rect 132677 330112 132682 330168
rect 132738 330112 154068 330168
rect 132677 330110 154068 330112
rect 132677 330107 132743 330110
rect 154062 330108 154068 330110
rect 154132 330108 154138 330172
rect 69606 329972 69612 330036
rect 69676 330034 69682 330036
rect 70158 330034 70164 330036
rect 69676 329974 70164 330034
rect 69676 329972 69682 329974
rect 70158 329972 70164 329974
rect 70228 330034 70234 330036
rect 133321 330034 133387 330037
rect 70228 330032 133387 330034
rect 70228 329976 133326 330032
rect 133382 329976 133387 330032
rect 70228 329974 133387 329976
rect 70228 329972 70234 329974
rect 133321 329971 133387 329974
rect 147581 330034 147647 330037
rect 177297 330034 177363 330037
rect 147581 330032 177363 330034
rect 147581 329976 147586 330032
rect 147642 329976 177302 330032
rect 177358 329976 177363 330032
rect 147581 329974 177363 329976
rect 147581 329971 147647 329974
rect 177297 329971 177363 329974
rect 131481 329898 131547 329901
rect 133086 329898 133092 329900
rect 131481 329896 133092 329898
rect 131481 329840 131486 329896
rect 131542 329840 133092 329896
rect 131481 329838 133092 329840
rect 131481 329835 131547 329838
rect 133086 329836 133092 329838
rect 133156 329836 133162 329900
rect 129733 329218 129799 329221
rect 211797 329218 211863 329221
rect 129733 329216 211863 329218
rect 129733 329160 129738 329216
rect 129794 329160 211802 329216
rect 211858 329160 211863 329216
rect 129733 329158 211863 329160
rect 129733 329155 129799 329158
rect 211797 329155 211863 329158
rect 68277 329082 68343 329085
rect 149053 329082 149119 329085
rect 68277 329080 149119 329082
rect 68277 329024 68282 329080
rect 68338 329024 149058 329080
rect 149114 329024 149119 329080
rect 68277 329022 149119 329024
rect 68277 329019 68343 329022
rect 149053 329019 149119 329022
rect 151077 329082 151143 329085
rect 157425 329082 157491 329085
rect 151077 329080 157491 329082
rect 151077 329024 151082 329080
rect 151138 329024 157430 329080
rect 157486 329024 157491 329080
rect 151077 329022 157491 329024
rect 151077 329019 151143 329022
rect 157425 329019 157491 329022
rect 153653 328674 153719 328677
rect 233969 328674 234035 328677
rect 153653 328672 234035 328674
rect 153653 328616 153658 328672
rect 153714 328616 233974 328672
rect 234030 328616 234035 328672
rect 153653 328614 234035 328616
rect 153653 328611 153719 328614
rect 233969 328611 234035 328614
rect 17217 328538 17283 328541
rect 115013 328538 115079 328541
rect 17217 328536 115079 328538
rect 17217 328480 17222 328536
rect 17278 328480 115018 328536
rect 115074 328480 115079 328536
rect 17217 328478 115079 328480
rect 17217 328475 17283 328478
rect 115013 328475 115079 328478
rect 122097 328538 122163 328541
rect 133086 328538 133092 328540
rect 122097 328536 133092 328538
rect 122097 328480 122102 328536
rect 122158 328480 133092 328536
rect 122097 328478 133092 328480
rect 122097 328475 122163 328478
rect 133086 328476 133092 328478
rect 133156 328476 133162 328540
rect 146201 328538 146267 328541
rect 151721 328538 151787 328541
rect 146201 328536 151787 328538
rect 146201 328480 146206 328536
rect 146262 328480 151726 328536
rect 151782 328480 151787 328536
rect 146201 328478 151787 328480
rect 146201 328475 146267 328478
rect 151721 328475 151787 328478
rect 67582 328340 67588 328404
rect 67652 328402 67658 328404
rect 68686 328402 68692 328404
rect 67652 328342 68692 328402
rect 67652 328340 67658 328342
rect 68686 328340 68692 328342
rect 68756 328340 68762 328404
rect 83641 327722 83707 327725
rect 84694 327722 84700 327724
rect 83641 327720 84700 327722
rect 83641 327664 83646 327720
rect 83702 327664 84700 327720
rect 83641 327662 84700 327664
rect 83641 327659 83707 327662
rect 84694 327660 84700 327662
rect 84764 327660 84770 327724
rect 148271 327722 148337 327725
rect 154246 327722 154252 327724
rect 148271 327720 154252 327722
rect 148271 327664 148276 327720
rect 148332 327664 154252 327720
rect 148271 327662 154252 327664
rect 148271 327659 148337 327662
rect 154246 327660 154252 327662
rect 154316 327660 154322 327724
rect 150382 327524 150388 327588
rect 150452 327586 150458 327588
rect 150709 327586 150775 327589
rect 150452 327584 150775 327586
rect 150452 327528 150714 327584
rect 150770 327528 150775 327584
rect 150452 327526 150775 327528
rect 150452 327524 150458 327526
rect 150709 327523 150775 327526
rect 152825 327586 152891 327589
rect 155718 327586 155724 327588
rect 152825 327584 155724 327586
rect 152825 327528 152830 327584
rect 152886 327528 155724 327584
rect 152825 327526 155724 327528
rect 152825 327523 152891 327526
rect 155718 327524 155724 327526
rect 155788 327524 155794 327588
rect 68686 327388 68692 327452
rect 68756 327450 68762 327452
rect 225413 327450 225479 327453
rect 68756 327448 225479 327450
rect 68756 327392 225418 327448
rect 225474 327392 225479 327448
rect 68756 327390 225479 327392
rect 68756 327388 68762 327390
rect 225413 327387 225479 327390
rect 7557 327314 7623 327317
rect 93853 327314 93919 327317
rect 7557 327312 93919 327314
rect 7557 327256 7562 327312
rect 7618 327256 93858 327312
rect 93914 327256 93919 327312
rect 7557 327254 93919 327256
rect 7557 327251 7623 327254
rect 93853 327251 93919 327254
rect 154389 327314 154455 327317
rect 238201 327314 238267 327317
rect 154389 327312 238267 327314
rect 154389 327256 154394 327312
rect 154450 327256 238206 327312
rect 238262 327256 238267 327312
rect 154389 327254 238267 327256
rect 154389 327251 154455 327254
rect 238201 327251 238267 327254
rect 66110 327116 66116 327180
rect 66180 327178 66186 327180
rect 68645 327178 68711 327181
rect 66180 327176 68711 327178
rect 66180 327120 68650 327176
rect 68706 327120 68711 327176
rect 66180 327118 68711 327120
rect 66180 327116 66186 327118
rect 68645 327115 68711 327118
rect 75729 327178 75795 327181
rect 75729 327176 77034 327178
rect 75729 327120 75734 327176
rect 75790 327120 77034 327176
rect 75729 327118 77034 327120
rect 75729 327115 75795 327118
rect 67214 326980 67220 327044
rect 67284 327042 67290 327044
rect 67357 327042 67423 327045
rect 70025 327042 70091 327045
rect 67284 327040 67423 327042
rect 67284 326984 67362 327040
rect 67418 326984 67423 327040
rect 67284 326982 67423 326984
rect 67284 326980 67290 326982
rect 67357 326979 67423 326982
rect 69430 327040 70091 327042
rect 69430 326984 70030 327040
rect 70086 326984 70091 327040
rect 69430 326982 70091 326984
rect 76974 327042 77034 327118
rect 77150 327116 77156 327180
rect 77220 327178 77226 327180
rect 77293 327178 77359 327181
rect 83917 327180 83983 327181
rect 77220 327176 77359 327178
rect 77220 327120 77298 327176
rect 77354 327120 77359 327176
rect 77220 327118 77359 327120
rect 77220 327116 77226 327118
rect 77293 327115 77359 327118
rect 77526 327118 83842 327178
rect 77526 327042 77586 327118
rect 76974 326982 77586 327042
rect 83782 327042 83842 327118
rect 83917 327176 83964 327180
rect 84028 327178 84034 327180
rect 202137 327178 202203 327181
rect 83917 327120 83922 327176
rect 83917 327116 83964 327120
rect 84028 327118 84074 327178
rect 84150 327176 202203 327178
rect 84150 327120 202142 327176
rect 202198 327120 202203 327176
rect 84150 327118 202203 327120
rect 84028 327116 84034 327118
rect 83917 327115 83983 327116
rect 84150 327042 84210 327118
rect 202137 327115 202203 327118
rect 83782 326982 84210 327042
rect 142889 327042 142955 327045
rect 143390 327042 143396 327044
rect 142889 327040 143396 327042
rect 142889 326984 142894 327040
rect 142950 326984 143396 327040
rect 142889 326982 143396 326984
rect 67173 326770 67239 326773
rect 69430 326770 69490 326982
rect 70025 326979 70091 326982
rect 142889 326979 142955 326982
rect 143390 326980 143396 326982
rect 143460 326980 143466 327044
rect 153101 327042 153167 327045
rect 154389 327042 154455 327045
rect 153101 327040 154314 327042
rect 153101 326984 153106 327040
rect 153162 326984 154314 327040
rect 153101 326982 154314 326984
rect 153101 326979 153167 326982
rect 67173 326768 69490 326770
rect 67173 326712 67178 326768
rect 67234 326740 69490 326768
rect 154254 326770 154314 326982
rect 154389 327040 161490 327042
rect 154389 326984 154394 327040
rect 154450 326984 161490 327040
rect 154389 326982 161490 326984
rect 154389 326979 154455 326982
rect 154849 326906 154915 326909
rect 157241 326906 157307 326909
rect 154849 326904 157307 326906
rect 154849 326848 154854 326904
rect 154910 326848 157246 326904
rect 157302 326848 157307 326904
rect 154849 326846 157307 326848
rect 161430 326906 161490 326982
rect 258165 326906 258231 326909
rect 161430 326904 258231 326906
rect 161430 326848 258170 326904
rect 258226 326848 258231 326904
rect 161430 326846 258231 326848
rect 154849 326843 154915 326846
rect 157241 326843 157307 326846
rect 258165 326843 258231 326846
rect 67234 326712 69460 326740
rect 67173 326710 69460 326712
rect 154254 326710 161490 326770
rect 67173 326707 67239 326710
rect 68553 326498 68619 326501
rect 156413 326498 156479 326501
rect 68553 326496 68938 326498
rect 68553 326440 68558 326496
rect 68614 326440 68938 326496
rect 68553 326438 68938 326440
rect 154652 326496 156479 326498
rect 154652 326440 156418 326496
rect 156474 326440 156479 326496
rect 154652 326438 156479 326440
rect 68553 326435 68619 326438
rect 21357 326226 21423 326229
rect 68645 326226 68711 326229
rect 21357 326224 68711 326226
rect 21357 326168 21362 326224
rect 21418 326168 68650 326224
rect 68706 326168 68711 326224
rect 21357 326166 68711 326168
rect 21357 326163 21423 326166
rect 68645 326163 68711 326166
rect 68878 325924 68938 326438
rect 156413 326435 156479 326438
rect 161430 326362 161490 326710
rect 243077 326362 243143 326365
rect 161430 326360 243143 326362
rect 161430 326304 243082 326360
rect 243138 326304 243143 326360
rect 161430 326302 243143 326304
rect 243077 326299 243143 326302
rect 157149 325410 157215 325413
rect 154652 325408 157215 325410
rect 154652 325352 157154 325408
rect 157210 325352 157215 325408
rect 154652 325350 157215 325352
rect 157149 325347 157215 325350
rect 154246 325212 154252 325276
rect 154316 325274 154322 325276
rect 167821 325274 167887 325277
rect 154316 325272 167887 325274
rect 154316 325216 167826 325272
rect 167882 325216 167887 325272
rect 154316 325214 167887 325216
rect 154316 325212 154322 325214
rect 167821 325211 167887 325214
rect 583293 325274 583359 325277
rect 583520 325274 584960 325364
rect 583293 325272 584960 325274
rect 583293 325216 583298 325272
rect 583354 325216 584960 325272
rect 583293 325214 584960 325216
rect 583293 325211 583359 325214
rect 583520 325124 584960 325214
rect 155718 324940 155724 325004
rect 155788 325002 155794 325004
rect 333973 325002 334039 325005
rect 155788 325000 334039 325002
rect 155788 324944 333978 325000
rect 334034 324944 334039 325000
rect 155788 324942 334039 324944
rect 155788 324940 155794 324942
rect 333973 324939 334039 324942
rect 66897 324866 66963 324869
rect 66897 324864 68908 324866
rect 66897 324808 66902 324864
rect 66958 324808 68908 324864
rect 66897 324806 68908 324808
rect 66897 324803 66963 324806
rect 156873 324322 156939 324325
rect 154652 324320 156939 324322
rect 154652 324264 156878 324320
rect 156934 324264 156939 324320
rect 154652 324262 156939 324264
rect 156873 324259 156939 324262
rect 66805 323778 66871 323781
rect 66805 323776 68908 323778
rect 66805 323720 66810 323776
rect 66866 323720 68908 323776
rect 66805 323718 68908 323720
rect 66805 323715 66871 323718
rect 154246 323580 154252 323644
rect 154316 323642 154322 323644
rect 232589 323642 232655 323645
rect 154316 323640 232655 323642
rect 154316 323584 232594 323640
rect 232650 323584 232655 323640
rect 154316 323582 232655 323584
rect 154316 323580 154322 323582
rect 232589 323579 232655 323582
rect 157425 323234 157491 323237
rect 161974 323234 161980 323236
rect 154652 323232 161980 323234
rect 154652 323176 157430 323232
rect 157486 323176 161980 323232
rect 154652 323174 161980 323176
rect 157425 323171 157491 323174
rect 161974 323172 161980 323174
rect 162044 323172 162050 323236
rect 67633 322690 67699 322693
rect 67633 322688 68908 322690
rect 67633 322632 67638 322688
rect 67694 322632 68908 322688
rect 67633 322630 68908 322632
rect 67633 322627 67699 322630
rect 157241 322146 157307 322149
rect 154652 322144 157307 322146
rect 154652 322088 157246 322144
rect 157302 322088 157307 322144
rect 154652 322086 157307 322088
rect 157241 322083 157307 322086
rect 67357 321602 67423 321605
rect 67357 321600 68908 321602
rect 67357 321544 67362 321600
rect 67418 321544 68908 321600
rect 67357 321542 68908 321544
rect 67357 321539 67423 321542
rect 66437 320514 66503 320517
rect 66437 320512 68908 320514
rect 66437 320456 66442 320512
rect 66498 320456 68908 320512
rect 66437 320454 68908 320456
rect 66437 320451 66503 320454
rect 154622 320378 154682 321028
rect 155166 320724 155172 320788
rect 155236 320786 155242 320788
rect 317413 320786 317479 320789
rect 155236 320784 317479 320786
rect 155236 320728 317418 320784
rect 317474 320728 317479 320784
rect 155236 320726 317479 320728
rect 155236 320724 155242 320726
rect 317413 320723 317479 320726
rect 170254 320378 170260 320380
rect 154622 320318 170260 320378
rect 170254 320316 170260 320318
rect 170324 320316 170330 320380
rect 66805 319426 66871 319429
rect 154622 319426 154682 319940
rect 158805 319426 158871 319429
rect 176009 319426 176075 319429
rect 66805 319424 68908 319426
rect -960 319290 480 319380
rect 66805 319368 66810 319424
rect 66866 319368 68908 319424
rect 66805 319366 68908 319368
rect 154622 319424 176075 319426
rect 154622 319368 158810 319424
rect 158866 319368 176014 319424
rect 176070 319368 176075 319424
rect 154622 319366 176075 319368
rect 66805 319363 66871 319366
rect 158805 319363 158871 319366
rect 176009 319363 176075 319366
rect 4061 319290 4127 319293
rect -960 319288 4127 319290
rect -960 319232 4066 319288
rect 4122 319232 4127 319288
rect -960 319230 4127 319232
rect -960 319140 480 319230
rect 4061 319227 4127 319230
rect 157241 318882 157307 318885
rect 154652 318880 157307 318882
rect 154652 318824 157246 318880
rect 157302 318824 157307 318880
rect 154652 318822 157307 318824
rect 157241 318819 157307 318822
rect 156454 318684 156460 318748
rect 156524 318746 156530 318748
rect 156597 318746 156663 318749
rect 156524 318744 156663 318746
rect 156524 318688 156602 318744
rect 156658 318688 156663 318744
rect 156524 318686 156663 318688
rect 156524 318684 156530 318686
rect 156597 318683 156663 318686
rect 66897 318338 66963 318341
rect 66897 318336 68908 318338
rect 66897 318280 66902 318336
rect 66958 318280 68908 318336
rect 66897 318278 68908 318280
rect 66897 318275 66963 318278
rect 155953 318066 156019 318069
rect 154652 318064 156019 318066
rect 154652 318008 155958 318064
rect 156014 318008 156019 318064
rect 154652 318006 156019 318008
rect 155953 318003 156019 318006
rect 66805 317522 66871 317525
rect 156597 317522 156663 317525
rect 249885 317522 249951 317525
rect 66805 317520 68908 317522
rect 66805 317464 66810 317520
rect 66866 317464 68908 317520
rect 66805 317462 68908 317464
rect 156597 317520 249951 317522
rect 156597 317464 156602 317520
rect 156658 317464 249890 317520
rect 249946 317464 249951 317520
rect 156597 317462 249951 317464
rect 66805 317459 66871 317462
rect 156597 317459 156663 317462
rect 249885 317459 249951 317462
rect 157241 316978 157307 316981
rect 154652 316976 157307 316978
rect 154652 316920 157246 316976
rect 157302 316920 157307 316976
rect 154652 316918 157307 316920
rect 157241 316915 157307 316918
rect 195237 316706 195303 316709
rect 320214 316706 320220 316708
rect 195237 316704 320220 316706
rect 195237 316648 195242 316704
rect 195298 316648 320220 316704
rect 195237 316646 320220 316648
rect 195237 316643 195303 316646
rect 320214 316644 320220 316646
rect 320284 316644 320290 316708
rect 67265 316434 67331 316437
rect 67265 316432 68908 316434
rect 67265 316376 67270 316432
rect 67326 316376 68908 316432
rect 67265 316374 68908 316376
rect 67265 316371 67331 316374
rect 156781 315890 156847 315893
rect 154652 315888 156847 315890
rect 154652 315832 156786 315888
rect 156842 315832 156847 315888
rect 154652 315830 156847 315832
rect 156781 315827 156847 315830
rect 66805 315346 66871 315349
rect 160829 315346 160895 315349
rect 182817 315346 182883 315349
rect 66805 315344 68908 315346
rect 66805 315288 66810 315344
rect 66866 315288 68908 315344
rect 66805 315286 68908 315288
rect 160829 315344 182883 315346
rect 160829 315288 160834 315344
rect 160890 315288 182822 315344
rect 182878 315288 182883 315344
rect 160829 315286 182883 315288
rect 66805 315283 66871 315286
rect 160829 315283 160895 315286
rect 182817 315283 182883 315286
rect 183001 315346 183067 315349
rect 222326 315346 222332 315348
rect 183001 315344 222332 315346
rect 183001 315288 183006 315344
rect 183062 315288 222332 315344
rect 183001 315286 222332 315288
rect 183001 315283 183067 315286
rect 222326 315284 222332 315286
rect 222396 315284 222402 315348
rect 157241 314802 157307 314805
rect 154652 314800 157307 314802
rect 154652 314744 157246 314800
rect 157302 314744 157307 314800
rect 154652 314742 157307 314744
rect 157241 314739 157307 314742
rect 196709 314802 196775 314805
rect 197261 314802 197327 314805
rect 294597 314802 294663 314805
rect 196709 314800 294663 314802
rect 196709 314744 196714 314800
rect 196770 314744 197266 314800
rect 197322 314744 294602 314800
rect 294658 314744 294663 314800
rect 196709 314742 294663 314744
rect 196709 314739 196775 314742
rect 197261 314739 197327 314742
rect 294597 314739 294663 314742
rect 66897 314258 66963 314261
rect 66897 314256 68908 314258
rect 66897 314200 66902 314256
rect 66958 314200 68908 314256
rect 66897 314198 68908 314200
rect 66897 314195 66963 314198
rect 215937 313986 216003 313989
rect 240777 313986 240843 313989
rect 215937 313984 240843 313986
rect 215937 313928 215942 313984
rect 215998 313928 240782 313984
rect 240838 313928 240843 313984
rect 215937 313926 240843 313928
rect 215937 313923 216003 313926
rect 240777 313923 240843 313926
rect 61653 313442 61719 313445
rect 61878 313442 61884 313444
rect 61653 313440 61884 313442
rect 61653 313384 61658 313440
rect 61714 313384 61884 313440
rect 61653 313382 61884 313384
rect 61653 313379 61719 313382
rect 61878 313380 61884 313382
rect 61948 313380 61954 313444
rect 154622 313306 154682 313684
rect 195237 313306 195303 313309
rect 154622 313304 195303 313306
rect 154622 313248 195242 313304
rect 195298 313248 195303 313304
rect 154622 313246 195303 313248
rect 195237 313243 195303 313246
rect 66805 313170 66871 313173
rect 66805 313168 68908 313170
rect 66805 313112 66810 313168
rect 66866 313112 68908 313168
rect 66805 313110 68908 313112
rect 66805 313107 66871 313110
rect 156413 312626 156479 312629
rect 154652 312624 156479 312626
rect 154652 312568 156418 312624
rect 156474 312568 156479 312624
rect 154652 312566 156479 312568
rect 156413 312563 156479 312566
rect 238017 312490 238083 312493
rect 256785 312490 256851 312493
rect 238017 312488 256851 312490
rect 238017 312432 238022 312488
rect 238078 312432 256790 312488
rect 256846 312432 256851 312488
rect 238017 312430 256851 312432
rect 238017 312427 238083 312430
rect 256785 312427 256851 312430
rect 66069 312082 66135 312085
rect 583109 312082 583175 312085
rect 583520 312082 584960 312172
rect 66069 312080 68908 312082
rect 66069 312024 66074 312080
rect 66130 312024 68908 312080
rect 66069 312022 68908 312024
rect 583109 312080 584960 312082
rect 583109 312024 583114 312080
rect 583170 312024 584960 312080
rect 583109 312022 584960 312024
rect 66069 312019 66135 312022
rect 583109 312019 583175 312022
rect 583520 311932 584960 312022
rect 157241 311538 157307 311541
rect 154652 311536 157307 311538
rect 154652 311480 157246 311536
rect 157302 311480 157307 311536
rect 154652 311478 157307 311480
rect 157241 311475 157307 311478
rect 66437 310994 66503 310997
rect 66437 310992 68908 310994
rect 66437 310936 66442 310992
rect 66498 310936 68908 310992
rect 66437 310934 68908 310936
rect 66437 310931 66503 310934
rect 230013 310722 230079 310725
rect 270718 310722 270724 310724
rect 230013 310720 270724 310722
rect 230013 310664 230018 310720
rect 230074 310664 270724 310720
rect 230013 310662 270724 310664
rect 230013 310659 230079 310662
rect 270718 310660 270724 310662
rect 270788 310660 270794 310724
rect 221549 310586 221615 310589
rect 315941 310586 316007 310589
rect 221549 310584 316007 310586
rect 221549 310528 221554 310584
rect 221610 310528 315946 310584
rect 316002 310528 316007 310584
rect 221549 310526 316007 310528
rect 221549 310523 221615 310526
rect 315941 310523 316007 310526
rect 156137 310450 156203 310453
rect 154652 310448 156203 310450
rect 154652 310392 156142 310448
rect 156198 310392 156203 310448
rect 154652 310390 156203 310392
rect 156137 310387 156203 310390
rect 66805 309906 66871 309909
rect 66805 309904 68908 309906
rect 66805 309848 66810 309904
rect 66866 309848 68908 309904
rect 66805 309846 68908 309848
rect 66805 309843 66871 309846
rect 157241 309634 157307 309637
rect 154652 309632 157307 309634
rect 154652 309576 157246 309632
rect 157302 309576 157307 309632
rect 154652 309574 157307 309576
rect 157241 309571 157307 309574
rect 209957 309362 210023 309365
rect 210509 309362 210575 309365
rect 269062 309362 269068 309364
rect 209957 309360 269068 309362
rect 209957 309304 209962 309360
rect 210018 309304 210514 309360
rect 210570 309304 269068 309360
rect 209957 309302 269068 309304
rect 209957 309299 210023 309302
rect 210509 309299 210575 309302
rect 269062 309300 269068 309302
rect 269132 309300 269138 309364
rect 209037 309226 209103 309229
rect 209405 309226 209471 309229
rect 339585 309226 339651 309229
rect 209037 309224 339651 309226
rect 209037 309168 209042 309224
rect 209098 309168 209410 309224
rect 209466 309168 339590 309224
rect 339646 309168 339651 309224
rect 209037 309166 339651 309168
rect 209037 309163 209103 309166
rect 209405 309163 209471 309166
rect 339585 309163 339651 309166
rect 67449 309090 67515 309093
rect 67633 309090 67699 309093
rect 206369 309090 206435 309093
rect 206921 309090 206987 309093
rect 67449 309088 68908 309090
rect 67449 309032 67454 309088
rect 67510 309032 67638 309088
rect 67694 309032 68908 309088
rect 67449 309030 68908 309032
rect 206369 309088 206987 309090
rect 206369 309032 206374 309088
rect 206430 309032 206926 309088
rect 206982 309032 206987 309088
rect 206369 309030 206987 309032
rect 67449 309027 67515 309030
rect 67633 309027 67699 309030
rect 206369 309027 206435 309030
rect 206921 309027 206987 309030
rect 156229 308546 156295 308549
rect 156689 308546 156755 308549
rect 154652 308544 156755 308546
rect 154652 308488 156234 308544
rect 156290 308488 156694 308544
rect 156750 308488 156755 308544
rect 154652 308486 156755 308488
rect 156229 308483 156295 308486
rect 156689 308483 156755 308486
rect 159449 308410 159515 308413
rect 197169 308410 197235 308413
rect 159449 308408 197235 308410
rect 159449 308352 159454 308408
rect 159510 308352 197174 308408
rect 197230 308352 197235 308408
rect 159449 308350 197235 308352
rect 159449 308347 159515 308350
rect 197169 308347 197235 308350
rect 66713 308002 66779 308005
rect 67214 308002 67220 308004
rect 66713 308000 67220 308002
rect 66713 307944 66718 308000
rect 66774 307944 67220 308000
rect 66713 307942 67220 307944
rect 66713 307939 66779 307942
rect 67214 307940 67220 307942
rect 67284 308002 67290 308004
rect 67284 307942 68908 308002
rect 67284 307940 67290 307942
rect 206921 307866 206987 307869
rect 258390 307866 258396 307868
rect 206921 307864 258396 307866
rect 206921 307808 206926 307864
rect 206982 307808 258396 307864
rect 206921 307806 258396 307808
rect 206921 307803 206987 307806
rect 258390 307804 258396 307806
rect 258460 307804 258466 307868
rect 67725 306914 67791 306917
rect 67725 306912 68908 306914
rect 67725 306856 67730 306912
rect 67786 306856 68908 306912
rect 67725 306854 68908 306856
rect 67725 306851 67791 306854
rect 154622 306778 154682 307428
rect 154622 306718 161490 306778
rect 161430 306506 161490 306718
rect 315941 306644 316007 306645
rect 315941 306642 315988 306644
rect 315896 306640 315988 306642
rect 316052 306642 316058 306644
rect 315896 306584 315946 306640
rect 315896 306582 315988 306584
rect 315941 306580 315988 306582
rect 316052 306582 316134 306642
rect 316052 306580 316058 306582
rect 315941 306579 316007 306580
rect 322054 306506 322060 306508
rect 161430 306446 322060 306506
rect 322054 306444 322060 306446
rect 322124 306444 322130 306508
rect 157241 306370 157307 306373
rect 315941 306372 316007 306373
rect 315941 306370 315988 306372
rect 154652 306368 157307 306370
rect -960 306234 480 306324
rect 154652 306312 157246 306368
rect 157302 306312 157307 306368
rect 154652 306310 157307 306312
rect 315896 306368 315988 306370
rect 316052 306370 316058 306372
rect 315896 306312 315946 306368
rect 315896 306310 315988 306312
rect 157241 306307 157307 306310
rect 315941 306308 315988 306310
rect 316052 306310 316134 306370
rect 316052 306308 316058 306310
rect 315941 306307 316007 306308
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 66897 305826 66963 305829
rect 66897 305824 68908 305826
rect 66897 305768 66902 305824
rect 66958 305768 68908 305824
rect 66897 305766 68908 305768
rect 66897 305763 66963 305766
rect 180057 305690 180123 305693
rect 189809 305690 189875 305693
rect 180057 305688 189875 305690
rect 180057 305632 180062 305688
rect 180118 305632 189814 305688
rect 189870 305632 189875 305688
rect 180057 305630 189875 305632
rect 180057 305627 180123 305630
rect 189809 305627 189875 305630
rect 157241 305282 157307 305285
rect 154652 305280 157307 305282
rect 154652 305224 157246 305280
rect 157302 305224 157307 305280
rect 154652 305222 157307 305224
rect 157241 305219 157307 305222
rect 210417 305010 210483 305013
rect 214741 305010 214807 305013
rect 583477 305010 583543 305013
rect 210417 305008 583543 305010
rect 210417 304952 210422 305008
rect 210478 304952 214746 305008
rect 214802 304952 583482 305008
rect 583538 304952 583543 305008
rect 210417 304950 583543 304952
rect 210417 304947 210483 304950
rect 214741 304947 214807 304950
rect 583477 304947 583543 304950
rect 66897 304738 66963 304741
rect 66897 304736 68908 304738
rect 66897 304680 66902 304736
rect 66958 304680 68908 304736
rect 66897 304678 68908 304680
rect 66897 304675 66963 304678
rect 157241 304194 157307 304197
rect 154652 304192 157307 304194
rect 154652 304136 157246 304192
rect 157302 304136 157307 304192
rect 154652 304134 157307 304136
rect 157241 304131 157307 304134
rect 160686 303724 160692 303788
rect 160756 303786 160762 303788
rect 160921 303786 160987 303789
rect 218646 303786 218652 303788
rect 160756 303784 218652 303786
rect 160756 303728 160926 303784
rect 160982 303728 218652 303784
rect 160756 303726 218652 303728
rect 160756 303724 160762 303726
rect 160921 303723 160987 303726
rect 218646 303724 218652 303726
rect 218716 303724 218722 303788
rect 66253 303650 66319 303653
rect 201677 303650 201743 303653
rect 583661 303650 583727 303653
rect 66253 303648 68908 303650
rect 66253 303592 66258 303648
rect 66314 303592 68908 303648
rect 66253 303590 68908 303592
rect 201677 303648 583727 303650
rect 201677 303592 201682 303648
rect 201738 303592 583666 303648
rect 583722 303592 583727 303648
rect 201677 303590 583727 303592
rect 66253 303587 66319 303590
rect 201677 303587 201743 303590
rect 583661 303587 583727 303590
rect 157241 303106 157307 303109
rect 154652 303104 157307 303106
rect 154652 303048 157246 303104
rect 157302 303048 157307 303104
rect 154652 303046 157307 303048
rect 157241 303043 157307 303046
rect 161974 302772 161980 302836
rect 162044 302834 162050 302836
rect 227846 302834 227852 302836
rect 162044 302774 227852 302834
rect 162044 302772 162050 302774
rect 227846 302772 227852 302774
rect 227916 302772 227922 302836
rect 66805 302562 66871 302565
rect 66805 302560 68908 302562
rect 66805 302504 66810 302560
rect 66866 302504 68908 302560
rect 66805 302502 68908 302504
rect 66805 302499 66871 302502
rect 239397 302426 239463 302429
rect 239581 302426 239647 302429
rect 287697 302426 287763 302429
rect 239397 302424 287763 302426
rect 239397 302368 239402 302424
rect 239458 302368 239586 302424
rect 239642 302368 287702 302424
rect 287758 302368 287763 302424
rect 239397 302366 287763 302368
rect 239397 302363 239463 302366
rect 239581 302363 239647 302366
rect 287697 302363 287763 302366
rect 206277 302290 206343 302293
rect 206645 302290 206711 302293
rect 582925 302290 582991 302293
rect 206277 302288 582991 302290
rect 206277 302232 206282 302288
rect 206338 302232 206650 302288
rect 206706 302232 582930 302288
rect 582986 302232 582991 302288
rect 206277 302230 582991 302232
rect 206277 302227 206343 302230
rect 206645 302227 206711 302230
rect 582925 302227 582991 302230
rect 199469 302154 199535 302157
rect 200941 302154 201007 302157
rect 199469 302152 201007 302154
rect 199469 302096 199474 302152
rect 199530 302096 200946 302152
rect 201002 302096 201007 302152
rect 199469 302094 201007 302096
rect 199469 302091 199535 302094
rect 200941 302091 201007 302094
rect 66805 301474 66871 301477
rect 154622 301474 154682 301988
rect 66805 301472 68908 301474
rect 66805 301416 66810 301472
rect 66866 301416 68908 301472
rect 66805 301414 68908 301416
rect 154622 301414 161490 301474
rect 66805 301411 66871 301414
rect 154622 300930 154682 301172
rect 161430 301066 161490 301414
rect 186814 301066 186820 301068
rect 161430 301006 186820 301066
rect 186814 301004 186820 301006
rect 186884 301004 186890 301068
rect 200941 301066 201007 301069
rect 201309 301066 201375 301069
rect 280797 301066 280863 301069
rect 200941 301064 280863 301066
rect 200941 301008 200946 301064
rect 201002 301008 201314 301064
rect 201370 301008 280802 301064
rect 280858 301008 280863 301064
rect 200941 301006 280863 301008
rect 200941 301003 201007 301006
rect 201309 301003 201375 301006
rect 280797 301003 280863 301006
rect 324957 300930 325023 300933
rect 154622 300928 325023 300930
rect 154622 300872 324962 300928
rect 325018 300872 325023 300928
rect 154622 300870 325023 300872
rect 324957 300867 325023 300870
rect 66253 300658 66319 300661
rect 66253 300656 68908 300658
rect 66253 300600 66258 300656
rect 66314 300600 68908 300656
rect 66253 300598 68908 300600
rect 66253 300595 66319 300598
rect 157241 300114 157307 300117
rect 154652 300112 157307 300114
rect 154652 300056 157246 300112
rect 157302 300056 157307 300112
rect 154652 300054 157307 300056
rect 157241 300051 157307 300054
rect 174537 300114 174603 300117
rect 174537 300112 180810 300114
rect 174537 300056 174542 300112
rect 174598 300056 180810 300112
rect 174537 300054 180810 300056
rect 174537 300051 174603 300054
rect 180750 299842 180810 300054
rect 193029 299842 193095 299845
rect 236821 299842 236887 299845
rect 180750 299840 236887 299842
rect 180750 299784 193034 299840
rect 193090 299784 236826 299840
rect 236882 299784 236887 299840
rect 180750 299782 236887 299784
rect 193029 299779 193095 299782
rect 236821 299779 236887 299782
rect 225597 299706 225663 299709
rect 227805 299706 227871 299709
rect 301221 299706 301287 299709
rect 225597 299704 301287 299706
rect 225597 299648 225602 299704
rect 225658 299648 227810 299704
rect 227866 299648 301226 299704
rect 301282 299648 301287 299704
rect 225597 299646 301287 299648
rect 225597 299643 225663 299646
rect 227805 299643 227871 299646
rect 301221 299643 301287 299646
rect 66805 299570 66871 299573
rect 236637 299570 236703 299573
rect 574737 299570 574803 299573
rect 66805 299568 68908 299570
rect 66805 299512 66810 299568
rect 66866 299512 68908 299568
rect 66805 299510 68908 299512
rect 236637 299568 574803 299570
rect 236637 299512 236642 299568
rect 236698 299512 574742 299568
rect 574798 299512 574803 299568
rect 236637 299510 574803 299512
rect 66805 299507 66871 299510
rect 236637 299507 236703 299510
rect 574737 299507 574803 299510
rect 157241 299026 157307 299029
rect 154652 299024 157307 299026
rect 154652 298968 157246 299024
rect 157302 298968 157307 299024
rect 154652 298966 157307 298968
rect 157241 298963 157307 298966
rect 582741 298754 582807 298757
rect 583520 298754 584960 298844
rect 582741 298752 584960 298754
rect 582741 298696 582746 298752
rect 582802 298696 584960 298752
rect 582741 298694 584960 298696
rect 582741 298691 582807 298694
rect 583520 298604 584960 298694
rect 67541 298482 67607 298485
rect 228357 298482 228423 298485
rect 229001 298482 229067 298485
rect 287094 298482 287100 298484
rect 67541 298480 68908 298482
rect 67541 298424 67546 298480
rect 67602 298424 68908 298480
rect 67541 298422 68908 298424
rect 228357 298480 287100 298482
rect 228357 298424 228362 298480
rect 228418 298424 229006 298480
rect 229062 298424 287100 298480
rect 228357 298422 287100 298424
rect 67541 298419 67607 298422
rect 228357 298419 228423 298422
rect 229001 298419 229067 298422
rect 287094 298420 287100 298422
rect 287164 298420 287170 298484
rect 170397 298346 170463 298349
rect 254117 298346 254183 298349
rect 170397 298344 254183 298346
rect 170397 298288 170402 298344
rect 170458 298288 254122 298344
rect 254178 298288 254183 298344
rect 170397 298286 254183 298288
rect 170397 298283 170463 298286
rect 254117 298283 254183 298286
rect 163589 298210 163655 298213
rect 249977 298210 250043 298213
rect 163589 298208 250043 298210
rect 163589 298152 163594 298208
rect 163650 298152 249982 298208
rect 250038 298152 250043 298208
rect 163589 298150 250043 298152
rect 163589 298147 163655 298150
rect 249977 298147 250043 298150
rect 156781 297938 156847 297941
rect 154652 297936 156847 297938
rect 154652 297880 156786 297936
rect 156842 297880 156847 297936
rect 154652 297878 156847 297880
rect 156781 297875 156847 297878
rect 176009 297530 176075 297533
rect 225965 297530 226031 297533
rect 176009 297528 226031 297530
rect 176009 297472 176014 297528
rect 176070 297472 225970 297528
rect 226026 297472 226031 297528
rect 176009 297470 226031 297472
rect 176009 297467 176075 297470
rect 225965 297467 226031 297470
rect 65926 297332 65932 297396
rect 65996 297394 66002 297396
rect 159357 297394 159423 297397
rect 237414 297394 237420 297396
rect 65996 297334 68908 297394
rect 159357 297392 237420 297394
rect 159357 297336 159362 297392
rect 159418 297336 237420 297392
rect 159357 297334 237420 297336
rect 65996 297332 66002 297334
rect 159357 297331 159423 297334
rect 237414 297332 237420 297334
rect 237484 297332 237490 297396
rect 156597 296850 156663 296853
rect 154652 296848 156663 296850
rect 154652 296792 156602 296848
rect 156658 296792 156663 296848
rect 154652 296790 156663 296792
rect 156597 296787 156663 296790
rect 222929 296850 222995 296853
rect 273294 296850 273300 296852
rect 222929 296848 273300 296850
rect 222929 296792 222934 296848
rect 222990 296792 273300 296848
rect 222929 296790 273300 296792
rect 222929 296787 222995 296790
rect 273294 296788 273300 296790
rect 273364 296788 273370 296852
rect 315941 296850 316007 296853
rect 316166 296850 316172 296852
rect 315896 296848 316172 296850
rect 315896 296792 315946 296848
rect 316002 296792 316172 296848
rect 315896 296790 316172 296792
rect 315941 296787 316007 296790
rect 316166 296788 316172 296790
rect 316236 296788 316242 296852
rect 315941 296714 316007 296717
rect 315896 296712 316050 296714
rect 315896 296656 315946 296712
rect 316002 296656 316050 296712
rect 315896 296654 316050 296656
rect 315941 296651 316050 296654
rect 315990 296580 316050 296651
rect 315982 296516 315988 296580
rect 316052 296516 316058 296580
rect 66437 296306 66503 296309
rect 66437 296304 68908 296306
rect 66437 296248 66442 296304
rect 66498 296248 68908 296304
rect 66437 296246 68908 296248
rect 66437 296243 66503 296246
rect 162761 296034 162827 296037
rect 180006 296034 180012 296036
rect 162761 296032 180012 296034
rect 162761 295976 162766 296032
rect 162822 295976 180012 296032
rect 162761 295974 180012 295976
rect 162761 295971 162827 295974
rect 180006 295972 180012 295974
rect 180076 295972 180082 296036
rect 157241 295762 157307 295765
rect 154652 295760 157307 295762
rect 154652 295704 157246 295760
rect 157302 295704 157307 295760
rect 154652 295702 157307 295704
rect 157241 295699 157307 295702
rect 154849 295626 154915 295629
rect 251449 295626 251515 295629
rect 154849 295624 251515 295626
rect 154849 295568 154854 295624
rect 154910 295568 251454 295624
rect 251510 295568 251515 295624
rect 154849 295566 251515 295568
rect 154849 295563 154915 295566
rect 251449 295563 251515 295566
rect 69422 295428 69428 295492
rect 69492 295428 69498 295492
rect 187049 295490 187115 295493
rect 241421 295490 241487 295493
rect 187049 295488 241487 295490
rect 187049 295432 187054 295488
rect 187110 295432 241426 295488
rect 241482 295432 241487 295488
rect 187049 295430 241487 295432
rect 67541 295218 67607 295221
rect 69430 295218 69490 295428
rect 187049 295427 187115 295430
rect 241421 295427 241487 295430
rect 67541 295216 69490 295218
rect 67541 295160 67546 295216
rect 67602 295188 69490 295216
rect 67602 295160 69460 295188
rect 67541 295158 69460 295160
rect 67541 295155 67607 295158
rect 156413 294674 156479 294677
rect 154652 294672 156479 294674
rect 154652 294616 156418 294672
rect 156474 294616 156479 294672
rect 154652 294614 156479 294616
rect 156413 294611 156479 294614
rect 160737 294538 160803 294541
rect 245929 294538 245995 294541
rect 160737 294536 245995 294538
rect 160737 294480 160742 294536
rect 160798 294480 245934 294536
rect 245990 294480 245995 294536
rect 160737 294478 245995 294480
rect 160737 294475 160803 294478
rect 245929 294475 245995 294478
rect 66253 294130 66319 294133
rect 66253 294128 68908 294130
rect 66253 294072 66258 294128
rect 66314 294072 68908 294128
rect 66253 294070 68908 294072
rect 66253 294067 66319 294070
rect 178677 293994 178743 293997
rect 211981 293994 212047 293997
rect 178677 293992 212047 293994
rect 178677 293936 178682 293992
rect 178738 293936 211986 293992
rect 212042 293936 212047 293992
rect 178677 293934 212047 293936
rect 178677 293931 178743 293934
rect 211981 293931 212047 293934
rect 216673 293994 216739 293997
rect 217685 293994 217751 293997
rect 255957 293994 256023 293997
rect 216673 293992 256023 293994
rect 216673 293936 216678 293992
rect 216734 293936 217690 293992
rect 217746 293936 255962 293992
rect 256018 293936 256023 293992
rect 216673 293934 256023 293936
rect 216673 293931 216739 293934
rect 217685 293931 217751 293934
rect 255957 293931 256023 293934
rect 161974 293586 161980 293588
rect 154652 293526 161980 293586
rect 161974 293524 161980 293526
rect 162044 293524 162050 293588
rect -960 293178 480 293268
rect 2773 293178 2839 293181
rect -960 293176 2839 293178
rect -960 293120 2778 293176
rect 2834 293120 2839 293176
rect -960 293118 2839 293120
rect -960 293028 480 293118
rect 2773 293115 2839 293118
rect 236821 293178 236887 293181
rect 242934 293178 242940 293180
rect 236821 293176 242940 293178
rect 236821 293120 236826 293176
rect 236882 293120 242940 293176
rect 236821 293118 242940 293120
rect 236821 293115 236887 293118
rect 242934 293116 242940 293118
rect 243004 293116 243010 293180
rect 66897 293042 66963 293045
rect 66897 293040 68908 293042
rect 66897 292984 66902 293040
rect 66958 292984 68908 293040
rect 66897 292982 68908 292984
rect 66897 292979 66963 292982
rect 211981 292906 212047 292909
rect 313273 292906 313339 292909
rect 211981 292904 313339 292906
rect 211981 292848 211986 292904
rect 212042 292848 313278 292904
rect 313334 292848 313339 292904
rect 211981 292846 313339 292848
rect 211981 292843 212047 292846
rect 313273 292843 313339 292846
rect 157241 292770 157307 292773
rect 154652 292768 157307 292770
rect 154652 292712 157246 292768
rect 157302 292712 157307 292768
rect 154652 292710 157307 292712
rect 157241 292707 157307 292710
rect 203517 292770 203583 292773
rect 204161 292770 204227 292773
rect 284334 292770 284340 292772
rect 203517 292768 284340 292770
rect 203517 292712 203522 292768
rect 203578 292712 204166 292768
rect 204222 292712 284340 292768
rect 203517 292710 284340 292712
rect 203517 292707 203583 292710
rect 204161 292707 204227 292710
rect 284334 292708 284340 292710
rect 284404 292708 284410 292772
rect 178534 292572 178540 292636
rect 178604 292634 178610 292636
rect 218605 292634 218671 292637
rect 178604 292632 218671 292634
rect 178604 292576 218610 292632
rect 218666 292576 218671 292632
rect 178604 292574 218671 292576
rect 178604 292572 178610 292574
rect 218605 292571 218671 292574
rect 197997 292498 198063 292501
rect 200389 292498 200455 292501
rect 201125 292498 201191 292501
rect 197997 292496 201191 292498
rect 197997 292440 198002 292496
rect 198058 292440 200394 292496
rect 200450 292440 201130 292496
rect 201186 292440 201191 292496
rect 197997 292438 201191 292440
rect 197997 292435 198063 292438
rect 200389 292435 200455 292438
rect 201125 292435 201191 292438
rect 66662 292164 66668 292228
rect 66732 292226 66738 292228
rect 66805 292226 66871 292229
rect 66732 292224 68908 292226
rect 66732 292168 66810 292224
rect 66866 292168 68908 292224
rect 66732 292166 68908 292168
rect 66732 292164 66738 292166
rect 66805 292163 66871 292166
rect 222837 291954 222903 291957
rect 223614 291954 223620 291956
rect 222837 291952 223620 291954
rect 222837 291896 222842 291952
rect 222898 291896 223620 291952
rect 222837 291894 223620 291896
rect 222837 291891 222903 291894
rect 223614 291892 223620 291894
rect 223684 291892 223690 291956
rect 201125 291818 201191 291821
rect 583385 291818 583451 291821
rect 201125 291816 583451 291818
rect 201125 291760 201130 291816
rect 201186 291760 583390 291816
rect 583446 291760 583451 291816
rect 201125 291758 583451 291760
rect 201125 291755 201191 291758
rect 583385 291755 583451 291758
rect 157241 291682 157307 291685
rect 154652 291680 157307 291682
rect 154652 291624 157246 291680
rect 157302 291624 157307 291680
rect 154652 291622 157307 291624
rect 157241 291619 157307 291622
rect 181621 291274 181687 291277
rect 239949 291274 240015 291277
rect 302877 291274 302943 291277
rect 181621 291272 302943 291274
rect 181621 291216 181626 291272
rect 181682 291216 239954 291272
rect 240010 291216 302882 291272
rect 302938 291216 302943 291272
rect 181621 291214 302943 291216
rect 181621 291211 181687 291214
rect 239949 291211 240015 291214
rect 302877 291211 302943 291214
rect 68878 290458 68938 291108
rect 157241 290594 157307 290597
rect 154652 290592 157307 290594
rect 154652 290536 157246 290592
rect 157302 290536 157307 290592
rect 154652 290534 157307 290536
rect 157241 290531 157307 290534
rect 64830 290398 68938 290458
rect 155217 290458 155283 290461
rect 200573 290458 200639 290461
rect 155217 290456 200639 290458
rect 155217 290400 155222 290456
rect 155278 290400 200578 290456
rect 200634 290400 200639 290456
rect 155217 290398 200639 290400
rect 53741 290050 53807 290053
rect 64830 290050 64890 290398
rect 155217 290395 155283 290398
rect 200573 290395 200639 290398
rect 197997 290186 198063 290189
rect 231117 290186 231183 290189
rect 197997 290184 231183 290186
rect 197997 290128 198002 290184
rect 198058 290128 231122 290184
rect 231178 290128 231183 290184
rect 197997 290126 231183 290128
rect 197997 290123 198063 290126
rect 231117 290123 231183 290126
rect 238569 290186 238635 290189
rect 253933 290186 253999 290189
rect 238569 290184 253999 290186
rect 238569 290128 238574 290184
rect 238630 290128 253938 290184
rect 253994 290128 253999 290184
rect 238569 290126 253999 290128
rect 238569 290123 238635 290126
rect 253933 290123 253999 290126
rect 53741 290048 64890 290050
rect 53741 289992 53746 290048
rect 53802 289992 64890 290048
rect 53741 289990 64890 289992
rect 66805 290050 66871 290053
rect 210877 290050 210943 290053
rect 270534 290050 270540 290052
rect 66805 290048 68908 290050
rect 66805 289992 66810 290048
rect 66866 289992 68908 290048
rect 66805 289990 68908 289992
rect 210877 290048 270540 290050
rect 210877 289992 210882 290048
rect 210938 289992 270540 290048
rect 210877 289990 270540 289992
rect 53741 289987 53807 289990
rect 66805 289987 66871 289990
rect 210877 289987 210943 289990
rect 270534 289988 270540 289990
rect 270604 289988 270610 290052
rect 202137 289914 202203 289917
rect 309133 289914 309199 289917
rect 202137 289912 309199 289914
rect 202137 289856 202142 289912
rect 202198 289856 309138 289912
rect 309194 289856 309199 289912
rect 202137 289854 309199 289856
rect 202137 289851 202203 289854
rect 309133 289851 309199 289854
rect 157241 289506 157307 289509
rect 154652 289504 157307 289506
rect 154652 289448 157246 289504
rect 157302 289448 157307 289504
rect 154652 289446 157307 289448
rect 157241 289443 157307 289446
rect 164969 289098 165035 289101
rect 178033 289098 178099 289101
rect 213453 289098 213519 289101
rect 583017 289098 583083 289101
rect 164969 289096 583083 289098
rect 164969 289040 164974 289096
rect 165030 289040 178038 289096
rect 178094 289040 213458 289096
rect 213514 289040 583022 289096
rect 583078 289040 583083 289096
rect 164969 289038 583083 289040
rect 164969 289035 165035 289038
rect 178033 289035 178099 289038
rect 213453 289035 213519 289038
rect 583017 289035 583083 289038
rect 66253 288962 66319 288965
rect 66253 288960 68908 288962
rect 66253 288904 66258 288960
rect 66314 288904 68908 288960
rect 66253 288902 68908 288904
rect 66253 288899 66319 288902
rect 198273 288554 198339 288557
rect 248505 288554 248571 288557
rect 198273 288552 248571 288554
rect 198273 288496 198278 288552
rect 198334 288496 248510 288552
rect 248566 288496 248571 288552
rect 198273 288494 248571 288496
rect 198273 288491 198339 288494
rect 248505 288491 248571 288494
rect 239489 288418 239555 288421
rect 243813 288418 243879 288421
rect 239489 288416 243879 288418
rect 66805 287874 66871 287877
rect 66805 287872 68908 287874
rect 66805 287816 66810 287872
rect 66866 287816 68908 287872
rect 66805 287814 68908 287816
rect 66805 287811 66871 287814
rect 154622 287738 154682 288388
rect 239489 288360 239494 288416
rect 239550 288360 243818 288416
rect 243874 288360 243879 288416
rect 239489 288358 243879 288360
rect 239489 288355 239555 288358
rect 243813 288355 243879 288358
rect 262949 287738 263015 287741
rect 306414 287738 306420 287740
rect 154622 287678 161490 287738
rect 161430 287466 161490 287678
rect 262949 287736 306420 287738
rect 262949 287680 262954 287736
rect 263010 287680 306420 287736
rect 262949 287678 306420 287680
rect 262949 287675 263015 287678
rect 306414 287676 306420 287678
rect 306484 287676 306490 287740
rect 192569 287602 192635 287605
rect 238109 287602 238175 287605
rect 192569 287600 238175 287602
rect 192569 287544 192574 287600
rect 192630 287544 238114 287600
rect 238170 287544 238175 287600
rect 192569 287542 238175 287544
rect 192569 287539 192635 287542
rect 238109 287539 238175 287542
rect 161430 287406 219450 287466
rect 191046 287330 191052 287332
rect 154652 287270 191052 287330
rect 191046 287268 191052 287270
rect 191116 287268 191122 287332
rect 219390 287194 219450 287406
rect 236453 287330 236519 287333
rect 261569 287330 261635 287333
rect 236453 287328 261635 287330
rect 236453 287272 236458 287328
rect 236514 287272 261574 287328
rect 261630 287272 261635 287328
rect 236453 287270 261635 287272
rect 236453 287267 236519 287270
rect 261569 287267 261635 287270
rect 231301 287194 231367 287197
rect 263961 287194 264027 287197
rect 315941 287196 316007 287197
rect 315941 287194 315988 287196
rect 219390 287192 264027 287194
rect 219390 287136 231306 287192
rect 231362 287136 263966 287192
rect 264022 287136 264027 287192
rect 219390 287134 264027 287136
rect 315896 287192 315988 287194
rect 316052 287194 316058 287196
rect 315896 287136 315946 287192
rect 315896 287134 315988 287136
rect 231301 287131 231367 287134
rect 263961 287131 264027 287134
rect 315941 287132 315988 287134
rect 316052 287134 316134 287194
rect 316052 287132 316058 287134
rect 315941 287131 316007 287132
rect 315941 287060 316007 287061
rect 315941 287058 315988 287060
rect 315896 287056 315988 287058
rect 316052 287058 316058 287060
rect 315896 287000 315946 287056
rect 315896 286998 315988 287000
rect 315941 286996 315988 286998
rect 316052 286998 316134 287058
rect 316052 286996 316058 286998
rect 315941 286995 316007 286996
rect 66989 286786 67055 286789
rect 66989 286784 68908 286786
rect 66989 286728 66994 286784
rect 67050 286728 68908 286784
rect 66989 286726 68908 286728
rect 66989 286723 67055 286726
rect 164233 286378 164299 286381
rect 218237 286378 218303 286381
rect 164233 286376 218303 286378
rect 164233 286320 164238 286376
rect 164294 286320 218242 286376
rect 218298 286320 218303 286376
rect 164233 286318 218303 286320
rect 164233 286315 164299 286318
rect 218237 286315 218303 286318
rect 156137 286242 156203 286245
rect 154652 286240 156203 286242
rect 154652 286184 156142 286240
rect 156198 286184 156203 286240
rect 154652 286182 156203 286184
rect 156137 286179 156203 286182
rect 242341 285970 242407 285973
rect 309225 285970 309291 285973
rect 242341 285968 309291 285970
rect 242341 285912 242346 285968
rect 242402 285912 309230 285968
rect 309286 285912 309291 285968
rect 242341 285910 309291 285912
rect 242341 285907 242407 285910
rect 309225 285907 309291 285910
rect 198733 285834 198799 285837
rect 218697 285834 218763 285837
rect 198733 285832 218763 285834
rect 198733 285776 198738 285832
rect 198794 285776 218702 285832
rect 218758 285776 218763 285832
rect 198733 285774 218763 285776
rect 198733 285771 198799 285774
rect 218697 285771 218763 285774
rect 221457 285834 221523 285837
rect 223798 285834 223804 285836
rect 221457 285832 223804 285834
rect 221457 285776 221462 285832
rect 221518 285776 223804 285832
rect 221457 285774 223804 285776
rect 221457 285771 221523 285774
rect 223798 285772 223804 285774
rect 223868 285772 223874 285836
rect 232497 285834 232563 285837
rect 276657 285834 276723 285837
rect 232497 285832 276723 285834
rect 232497 285776 232502 285832
rect 232558 285776 276662 285832
rect 276718 285776 276723 285832
rect 232497 285774 276723 285776
rect 232497 285771 232563 285774
rect 276657 285771 276723 285774
rect 66805 285698 66871 285701
rect 204253 285698 204319 285701
rect 205173 285698 205239 285701
rect 66805 285696 68908 285698
rect 66805 285640 66810 285696
rect 66866 285640 68908 285696
rect 66805 285638 68908 285640
rect 204253 285696 205239 285698
rect 204253 285640 204258 285696
rect 204314 285640 205178 285696
rect 205234 285640 205239 285696
rect 204253 285638 205239 285640
rect 66805 285635 66871 285638
rect 204253 285635 204319 285638
rect 205173 285635 205239 285638
rect 220721 285698 220787 285701
rect 222101 285698 222167 285701
rect 220721 285696 222167 285698
rect 220721 285640 220726 285696
rect 220782 285640 222106 285696
rect 222162 285640 222167 285696
rect 220721 285638 222167 285640
rect 220721 285635 220787 285638
rect 222101 285635 222167 285638
rect 223614 285636 223620 285700
rect 223684 285698 223690 285700
rect 223941 285698 224007 285701
rect 223684 285696 224007 285698
rect 223684 285640 223946 285696
rect 224002 285640 224007 285696
rect 223684 285638 224007 285640
rect 223684 285636 223690 285638
rect 223941 285635 224007 285638
rect 583520 285276 584960 285516
rect 157241 285154 157307 285157
rect 154652 285152 157307 285154
rect 154652 285096 157246 285152
rect 157302 285096 157307 285152
rect 154652 285094 157307 285096
rect 157241 285091 157307 285094
rect 211797 284882 211863 284885
rect 212349 284882 212415 284885
rect 216673 284882 216739 284885
rect 211797 284880 216739 284882
rect 211797 284824 211802 284880
rect 211858 284824 212354 284880
rect 212410 284824 216678 284880
rect 216734 284824 216739 284880
rect 211797 284822 216739 284824
rect 211797 284819 211863 284822
rect 212349 284819 212415 284822
rect 216673 284819 216739 284822
rect 197302 284684 197308 284748
rect 197372 284746 197378 284748
rect 232773 284746 232839 284749
rect 197372 284744 232839 284746
rect 197372 284688 232778 284744
rect 232834 284688 232839 284744
rect 197372 284686 232839 284688
rect 197372 284684 197378 284686
rect 232773 284683 232839 284686
rect 67081 284610 67147 284613
rect 176009 284610 176075 284613
rect 204253 284610 204319 284613
rect 67081 284608 68908 284610
rect 67081 284552 67086 284608
rect 67142 284552 68908 284608
rect 67081 284550 68908 284552
rect 176009 284608 204319 284610
rect 176009 284552 176014 284608
rect 176070 284552 204258 284608
rect 204314 284552 204319 284608
rect 176009 284550 204319 284552
rect 67081 284547 67147 284550
rect 176009 284547 176075 284550
rect 204253 284547 204319 284550
rect 238109 284610 238175 284613
rect 245694 284610 245700 284612
rect 238109 284608 245700 284610
rect 238109 284552 238114 284608
rect 238170 284552 245700 284608
rect 238109 284550 245700 284552
rect 238109 284547 238175 284550
rect 245694 284548 245700 284550
rect 245764 284548 245770 284612
rect 230473 284474 230539 284477
rect 231669 284474 231735 284477
rect 290457 284474 290523 284477
rect 230473 284472 290523 284474
rect 230473 284416 230478 284472
rect 230534 284416 231674 284472
rect 231730 284416 290462 284472
rect 290518 284416 290523 284472
rect 230473 284414 290523 284416
rect 230473 284411 230539 284414
rect 231669 284411 231735 284414
rect 290457 284411 290523 284414
rect 156781 284338 156847 284341
rect 154652 284336 156847 284338
rect 154652 284280 156786 284336
rect 156842 284280 156847 284336
rect 154652 284278 156847 284280
rect 156781 284275 156847 284278
rect 159357 284338 159423 284341
rect 206093 284338 206159 284341
rect 159357 284336 206159 284338
rect 159357 284280 159362 284336
rect 159418 284280 206098 284336
rect 206154 284280 206159 284336
rect 159357 284278 206159 284280
rect 159357 284275 159423 284278
rect 206093 284275 206159 284278
rect 217542 284276 217548 284340
rect 217612 284338 217618 284340
rect 220077 284338 220143 284341
rect 217612 284336 220143 284338
rect 217612 284280 220082 284336
rect 220138 284280 220143 284336
rect 217612 284278 220143 284280
rect 217612 284276 217618 284278
rect 220077 284275 220143 284278
rect 224217 284338 224283 284341
rect 224902 284338 224908 284340
rect 224217 284336 224908 284338
rect 224217 284280 224222 284336
rect 224278 284280 224908 284336
rect 224217 284278 224908 284280
rect 224217 284275 224283 284278
rect 224902 284276 224908 284278
rect 224972 284276 224978 284340
rect 226977 284338 227043 284341
rect 238518 284338 238524 284340
rect 226977 284336 238524 284338
rect 226977 284280 226982 284336
rect 227038 284280 238524 284336
rect 226977 284278 238524 284280
rect 226977 284275 227043 284278
rect 238518 284276 238524 284278
rect 238588 284276 238594 284340
rect 240041 284338 240107 284341
rect 583017 284338 583083 284341
rect 240041 284336 583083 284338
rect 240041 284280 240046 284336
rect 240102 284280 583022 284336
rect 583078 284280 583083 284336
rect 240041 284278 583083 284280
rect 240041 284275 240107 284278
rect 583017 284275 583083 284278
rect 243169 284202 243235 284205
rect 243169 284200 243554 284202
rect 243169 284144 243174 284200
rect 243230 284144 243554 284200
rect 243169 284142 243554 284144
rect 243169 284139 243235 284142
rect 201953 284066 202019 284069
rect 180750 284064 202019 284066
rect 180750 284008 201958 284064
rect 202014 284008 202019 284064
rect 180750 284006 202019 284008
rect 66621 283794 66687 283797
rect 66621 283792 68908 283794
rect 66621 283736 66626 283792
rect 66682 283736 68908 283792
rect 66621 283734 68908 283736
rect 66621 283731 66687 283734
rect 160829 283522 160895 283525
rect 180750 283522 180810 284006
rect 201953 284003 202019 284006
rect 216029 284066 216095 284069
rect 216438 284066 216444 284068
rect 216029 284064 216444 284066
rect 216029 284008 216034 284064
rect 216090 284008 216444 284064
rect 216029 284006 216444 284008
rect 216029 284003 216095 284006
rect 216438 284004 216444 284006
rect 216508 284004 216514 284068
rect 205357 283932 205423 283933
rect 205357 283930 205404 283932
rect 205312 283928 205404 283930
rect 205312 283872 205362 283928
rect 205312 283870 205404 283872
rect 205357 283868 205404 283870
rect 205468 283868 205474 283932
rect 211613 283930 211679 283933
rect 214465 283932 214531 283933
rect 212390 283930 212396 283932
rect 211613 283928 212396 283930
rect 211613 283872 211618 283928
rect 211674 283872 212396 283928
rect 211613 283870 212396 283872
rect 205357 283867 205423 283868
rect 211613 283867 211679 283870
rect 212390 283868 212396 283870
rect 212460 283868 212466 283932
rect 214414 283930 214420 283932
rect 214374 283870 214420 283930
rect 214484 283928 214531 283932
rect 214526 283872 214531 283928
rect 214414 283868 214420 283870
rect 214484 283868 214531 283872
rect 215518 283868 215524 283932
rect 215588 283930 215594 283932
rect 215937 283930 216003 283933
rect 215588 283928 216003 283930
rect 215588 283872 215942 283928
rect 215998 283872 216003 283928
rect 215588 283870 216003 283872
rect 215588 283868 215594 283870
rect 214465 283867 214531 283868
rect 215937 283867 216003 283870
rect 226793 283930 226859 283933
rect 227478 283930 227484 283932
rect 226793 283928 227484 283930
rect 226793 283872 226798 283928
rect 226854 283872 227484 283928
rect 226793 283870 227484 283872
rect 226793 283867 226859 283870
rect 227478 283868 227484 283870
rect 227548 283868 227554 283932
rect 236269 283930 236335 283933
rect 237230 283930 237236 283932
rect 236269 283928 237236 283930
rect 236269 283872 236274 283928
rect 236330 283872 237236 283928
rect 236269 283870 237236 283872
rect 236269 283867 236335 283870
rect 237230 283868 237236 283870
rect 237300 283868 237306 283932
rect 195329 283794 195395 283797
rect 195329 283792 200284 283794
rect 195329 283736 195334 283792
rect 195390 283736 200284 283792
rect 243494 283764 243554 284142
rect 244222 284140 244228 284204
rect 244292 284202 244298 284204
rect 244292 284142 248430 284202
rect 244292 284140 244298 284142
rect 243629 284066 243695 284069
rect 244222 284066 244228 284068
rect 243629 284064 244228 284066
rect 243629 284008 243634 284064
rect 243690 284008 244228 284064
rect 243629 284006 244228 284008
rect 243629 284003 243695 284006
rect 244222 284004 244228 284006
rect 244292 284004 244298 284068
rect 248370 284066 248430 284142
rect 307017 284066 307083 284069
rect 248370 284064 307083 284066
rect 248370 284008 307022 284064
rect 307078 284008 307083 284064
rect 248370 284006 307083 284008
rect 307017 284003 307083 284006
rect 195329 283734 200284 283736
rect 195329 283731 195395 283734
rect 160829 283520 180810 283522
rect 160829 283464 160834 283520
rect 160890 283464 180810 283520
rect 160829 283462 180810 283464
rect 160829 283459 160895 283462
rect 157149 283250 157215 283253
rect 244273 283250 244339 283253
rect 245377 283250 245443 283253
rect 154652 283248 157215 283250
rect 154652 283192 157154 283248
rect 157210 283192 157215 283248
rect 154652 283190 157215 283192
rect 244076 283248 245443 283250
rect 244076 283192 244278 283248
rect 244334 283192 245382 283248
rect 245438 283192 245443 283248
rect 244076 283190 245443 283192
rect 157149 283187 157215 283190
rect 244273 283187 244339 283190
rect 245377 283187 245443 283190
rect 198181 282978 198247 282981
rect 198181 282976 200284 282978
rect 198181 282920 198186 282976
rect 198242 282920 200284 282976
rect 198181 282918 200284 282920
rect 198181 282915 198247 282918
rect 66345 282706 66411 282709
rect 66345 282704 68908 282706
rect 66345 282648 66350 282704
rect 66406 282648 68908 282704
rect 66345 282646 68908 282648
rect 66345 282643 66411 282646
rect 197353 282434 197419 282437
rect 245653 282434 245719 282437
rect 197353 282432 200284 282434
rect 197353 282376 197358 282432
rect 197414 282376 200284 282432
rect 197353 282374 200284 282376
rect 244076 282432 245719 282434
rect 244076 282376 245658 282432
rect 245714 282376 245719 282432
rect 244076 282374 245719 282376
rect 197353 282371 197419 282374
rect 245653 282371 245719 282374
rect 157241 282162 157307 282165
rect 154652 282160 157307 282162
rect 154652 282104 157246 282160
rect 157302 282104 157307 282160
rect 154652 282102 157307 282104
rect 157241 282099 157307 282102
rect 245694 282100 245700 282164
rect 245764 282162 245770 282164
rect 258717 282162 258783 282165
rect 245764 282160 258783 282162
rect 245764 282104 258722 282160
rect 258778 282104 258783 282160
rect 245764 282102 258783 282104
rect 245764 282100 245770 282102
rect 258717 282099 258783 282102
rect 67449 281618 67515 281621
rect 185577 281618 185643 281621
rect 246113 281618 246179 281621
rect 67449 281616 68908 281618
rect 67449 281560 67454 281616
rect 67510 281560 68908 281616
rect 67449 281558 68908 281560
rect 185577 281616 200284 281618
rect 185577 281560 185582 281616
rect 185638 281560 200284 281616
rect 185577 281558 200284 281560
rect 244076 281616 246179 281618
rect 244076 281560 246118 281616
rect 246174 281560 246179 281616
rect 244076 281558 246179 281560
rect 67449 281555 67515 281558
rect 185577 281555 185643 281558
rect 246113 281555 246179 281558
rect 157241 281074 157307 281077
rect 244406 281074 244412 281076
rect 154652 281072 157307 281074
rect 154652 281016 157246 281072
rect 157302 281016 157307 281072
rect 154652 281014 157307 281016
rect 244076 281014 244412 281074
rect 157241 281011 157307 281014
rect 244406 281012 244412 281014
rect 244476 281074 244482 281076
rect 245653 281074 245719 281077
rect 244476 281072 245719 281074
rect 244476 281016 245658 281072
rect 245714 281016 245719 281072
rect 244476 281014 245719 281016
rect 244476 281012 244482 281014
rect 245653 281011 245719 281014
rect 182909 280938 182975 280941
rect 197302 280938 197308 280940
rect 182909 280936 197308 280938
rect 182909 280880 182914 280936
rect 182970 280880 197308 280936
rect 182909 280878 197308 280880
rect 182909 280875 182975 280878
rect 197302 280876 197308 280878
rect 197372 280876 197378 280940
rect 197353 280802 197419 280805
rect 197353 280800 200284 280802
rect 197353 280744 197358 280800
rect 197414 280744 200284 280800
rect 197353 280742 200284 280744
rect 197353 280739 197419 280742
rect 66805 280530 66871 280533
rect 66805 280528 68908 280530
rect 66805 280472 66810 280528
rect 66866 280472 68908 280528
rect 66805 280470 68908 280472
rect 66805 280467 66871 280470
rect 197445 280258 197511 280261
rect 246113 280258 246179 280261
rect 197445 280256 200284 280258
rect -960 279972 480 280212
rect 197445 280200 197450 280256
rect 197506 280200 200284 280256
rect 197445 280198 200284 280200
rect 244076 280256 246179 280258
rect 244076 280200 246118 280256
rect 246174 280200 246179 280256
rect 244076 280198 246179 280200
rect 197445 280195 197511 280198
rect 246113 280195 246179 280198
rect 157057 279986 157123 279989
rect 154652 279984 157123 279986
rect 154652 279928 157062 279984
rect 157118 279928 157123 279984
rect 154652 279926 157123 279928
rect 157057 279923 157123 279926
rect 66621 279442 66687 279445
rect 67766 279442 67772 279444
rect 66621 279440 67772 279442
rect 66621 279384 66626 279440
rect 66682 279384 67772 279440
rect 66621 279382 67772 279384
rect 66621 279379 66687 279382
rect 67766 279380 67772 279382
rect 67836 279442 67842 279444
rect 197353 279442 197419 279445
rect 246113 279442 246179 279445
rect 67836 279382 68908 279442
rect 197353 279440 200284 279442
rect 197353 279384 197358 279440
rect 197414 279384 200284 279440
rect 197353 279382 200284 279384
rect 244076 279440 246179 279442
rect 244076 279384 246118 279440
rect 246174 279384 246179 279440
rect 244076 279382 246179 279384
rect 67836 279380 67842 279382
rect 197353 279379 197419 279382
rect 246113 279379 246179 279382
rect 156965 278898 157031 278901
rect 244641 278898 244707 278901
rect 154652 278896 157031 278898
rect 154652 278840 156970 278896
rect 157026 278840 157031 278896
rect 154652 278838 157031 278840
rect 244076 278896 244707 278898
rect 244076 278840 244646 278896
rect 244702 278840 244707 278896
rect 244076 278838 244707 278840
rect 156965 278835 157031 278838
rect 244641 278835 244707 278838
rect 197353 278626 197419 278629
rect 197353 278624 200284 278626
rect 197353 278568 197358 278624
rect 197414 278568 200284 278624
rect 197353 278566 200284 278568
rect 197353 278563 197419 278566
rect 67357 278354 67423 278357
rect 67357 278352 68908 278354
rect 67357 278296 67362 278352
rect 67418 278296 68908 278352
rect 67357 278294 68908 278296
rect 67357 278291 67423 278294
rect 167729 278082 167795 278085
rect 195973 278082 196039 278085
rect 167729 278080 196039 278082
rect 167729 278024 167734 278080
rect 167790 278024 195978 278080
rect 196034 278024 196039 278080
rect 167729 278022 196039 278024
rect 167729 278019 167795 278022
rect 195973 278019 196039 278022
rect 198089 278082 198155 278085
rect 247125 278082 247191 278085
rect 198089 278080 200284 278082
rect 198089 278024 198094 278080
rect 198150 278024 200284 278080
rect 198089 278022 200284 278024
rect 244076 278080 247191 278082
rect 244076 278024 247130 278080
rect 247186 278024 247191 278080
rect 244076 278022 247191 278024
rect 198089 278019 198155 278022
rect 247125 278019 247191 278022
rect 156505 277810 156571 277813
rect 154652 277808 156571 277810
rect 154652 277752 156510 277808
rect 156566 277752 156571 277808
rect 154652 277750 156571 277752
rect 156505 277747 156571 277750
rect 246113 277538 246179 277541
rect 315941 277538 316007 277541
rect 316166 277538 316172 277540
rect 244076 277536 246179 277538
rect 244076 277480 246118 277536
rect 246174 277480 246179 277536
rect 244076 277478 246179 277480
rect 315896 277536 316172 277538
rect 315896 277480 315946 277536
rect 316002 277480 316172 277536
rect 315896 277478 316172 277480
rect 246113 277475 246179 277478
rect 315941 277475 316007 277478
rect 316166 277476 316172 277478
rect 316236 277476 316242 277540
rect 315941 277404 316007 277405
rect 315941 277402 315988 277404
rect 315896 277400 315988 277402
rect 316052 277402 316058 277404
rect 315896 277344 315946 277400
rect 315896 277342 315988 277344
rect 315941 277340 315988 277342
rect 316052 277342 316134 277402
rect 316052 277340 316058 277342
rect 315941 277339 316007 277340
rect 66253 277266 66319 277269
rect 66253 277264 68908 277266
rect 66253 277208 66258 277264
rect 66314 277208 68908 277264
rect 66253 277206 68908 277208
rect 66253 277203 66319 277206
rect 154665 276994 154731 276997
rect 154622 276992 154731 276994
rect 154622 276936 154670 276992
rect 154726 276936 154731 276992
rect 154622 276931 154731 276936
rect 193029 276994 193095 276997
rect 200254 276994 200314 277236
rect 193029 276992 200314 276994
rect 193029 276936 193034 276992
rect 193090 276936 200314 276992
rect 193029 276934 200314 276936
rect 193029 276931 193095 276934
rect 66161 276178 66227 276181
rect 154622 276178 154682 276931
rect 197353 276722 197419 276725
rect 246021 276722 246087 276725
rect 197353 276720 200284 276722
rect 197353 276664 197358 276720
rect 197414 276664 200284 276720
rect 197353 276662 200284 276664
rect 244076 276720 246087 276722
rect 244076 276664 246026 276720
rect 246082 276664 246087 276720
rect 244076 276662 246087 276664
rect 197353 276659 197419 276662
rect 246021 276659 246087 276662
rect 66161 276176 68908 276178
rect 66161 276120 66166 276176
rect 66222 276120 68908 276176
rect 66161 276118 68908 276120
rect 154622 276118 161490 276178
rect 66161 276115 66227 276118
rect 161430 276042 161490 276118
rect 187141 276042 187207 276045
rect 161430 276040 187207 276042
rect 161430 275984 187146 276040
rect 187202 275984 187207 276040
rect 161430 275982 187207 275984
rect 187141 275979 187207 275982
rect 157241 275906 157307 275909
rect 245929 275906 245995 275909
rect 154652 275904 157307 275906
rect 154652 275848 157246 275904
rect 157302 275848 157307 275904
rect 244076 275904 245995 275906
rect 154652 275846 157307 275848
rect 157241 275843 157307 275846
rect 67357 275362 67423 275365
rect 160921 275362 160987 275365
rect 200254 275362 200314 275876
rect 244076 275848 245934 275904
rect 245990 275848 245995 275904
rect 244076 275846 245995 275848
rect 245929 275843 245995 275846
rect 248454 275362 248460 275364
rect 67357 275360 68908 275362
rect 67357 275304 67362 275360
rect 67418 275304 68908 275360
rect 67357 275302 68908 275304
rect 160921 275360 200314 275362
rect 160921 275304 160926 275360
rect 160982 275304 200314 275360
rect 160921 275302 200314 275304
rect 244076 275302 248460 275362
rect 67357 275299 67423 275302
rect 160921 275299 160987 275302
rect 248454 275300 248460 275302
rect 248524 275300 248530 275364
rect 197445 275090 197511 275093
rect 197445 275088 200284 275090
rect 197445 275032 197450 275088
rect 197506 275032 200284 275088
rect 197445 275030 200284 275032
rect 197445 275027 197511 275030
rect 157241 274818 157307 274821
rect 154652 274816 157307 274818
rect 154652 274760 157246 274816
rect 157302 274760 157307 274816
rect 154652 274758 157307 274760
rect 157241 274755 157307 274758
rect 197353 274546 197419 274549
rect 245929 274546 245995 274549
rect 197353 274544 200284 274546
rect 197353 274488 197358 274544
rect 197414 274488 200284 274544
rect 197353 274486 200284 274488
rect 244076 274544 245995 274546
rect 244076 274488 245934 274544
rect 245990 274488 245995 274544
rect 244076 274486 245995 274488
rect 197353 274483 197419 274486
rect 245929 274483 245995 274486
rect 67081 274274 67147 274277
rect 67081 274272 68908 274274
rect 67081 274216 67086 274272
rect 67142 274216 68908 274272
rect 67081 274214 68908 274216
rect 67081 274211 67147 274214
rect 157241 273730 157307 273733
rect 154652 273728 157307 273730
rect 154652 273672 157246 273728
rect 157302 273672 157307 273728
rect 154652 273670 157307 273672
rect 157241 273667 157307 273670
rect 197353 273730 197419 273733
rect 245837 273730 245903 273733
rect 197353 273728 200284 273730
rect 197353 273672 197358 273728
rect 197414 273672 200284 273728
rect 197353 273670 200284 273672
rect 244076 273728 245903 273730
rect 244076 273672 245842 273728
rect 245898 273672 245903 273728
rect 244076 273670 245903 273672
rect 197353 273667 197419 273670
rect 245837 273667 245903 273670
rect 66989 273186 67055 273189
rect 245929 273186 245995 273189
rect 66989 273184 68908 273186
rect 66989 273128 66994 273184
rect 67050 273128 68908 273184
rect 66989 273126 68908 273128
rect 244076 273184 245995 273186
rect 244076 273128 245934 273184
rect 245990 273128 245995 273184
rect 244076 273126 245995 273128
rect 66989 273123 67055 273126
rect 245929 273123 245995 273126
rect 197353 272914 197419 272917
rect 197353 272912 200284 272914
rect 197353 272856 197358 272912
rect 197414 272856 200284 272912
rect 197353 272854 200284 272856
rect 197353 272851 197419 272854
rect 157241 272642 157307 272645
rect 154652 272640 157307 272642
rect 154652 272584 157246 272640
rect 157302 272584 157307 272640
rect 154652 272582 157307 272584
rect 157241 272579 157307 272582
rect 245837 272370 245903 272373
rect 244076 272368 245903 272370
rect 66805 272098 66871 272101
rect 66805 272096 68908 272098
rect 66805 272040 66810 272096
rect 66866 272040 68908 272096
rect 66805 272038 68908 272040
rect 66805 272035 66871 272038
rect 188337 271962 188403 271965
rect 200254 271962 200314 272340
rect 244076 272312 245842 272368
rect 245898 272312 245903 272368
rect 244076 272310 245903 272312
rect 245837 272307 245903 272310
rect 580257 272234 580323 272237
rect 583520 272234 584960 272324
rect 580257 272232 584960 272234
rect 580257 272176 580262 272232
rect 580318 272176 584960 272232
rect 580257 272174 584960 272176
rect 580257 272171 580323 272174
rect 583520 272084 584960 272174
rect 188337 271960 200314 271962
rect 188337 271904 188342 271960
rect 188398 271904 200314 271960
rect 188337 271902 200314 271904
rect 188337 271899 188403 271902
rect 157241 271554 157307 271557
rect 154652 271552 157307 271554
rect 154652 271496 157246 271552
rect 157302 271496 157307 271552
rect 154652 271494 157307 271496
rect 157241 271491 157307 271494
rect 197353 271554 197419 271557
rect 245745 271554 245811 271557
rect 197353 271552 200284 271554
rect 197353 271496 197358 271552
rect 197414 271496 200284 271552
rect 197353 271494 200284 271496
rect 244076 271552 245811 271554
rect 244076 271496 245750 271552
rect 245806 271496 245811 271552
rect 244076 271494 245811 271496
rect 197353 271491 197419 271494
rect 245745 271491 245811 271494
rect 66805 271010 66871 271013
rect 197445 271010 197511 271013
rect 245653 271010 245719 271013
rect 246297 271010 246363 271013
rect 66805 271008 68908 271010
rect 66805 270952 66810 271008
rect 66866 270952 68908 271008
rect 66805 270950 68908 270952
rect 197445 271008 200284 271010
rect 197445 270952 197450 271008
rect 197506 270952 200284 271008
rect 197445 270950 200284 270952
rect 244076 271008 246363 271010
rect 244076 270952 245658 271008
rect 245714 270952 246302 271008
rect 246358 270952 246363 271008
rect 244076 270950 246363 270952
rect 66805 270947 66871 270950
rect 197445 270947 197511 270950
rect 245653 270947 245719 270950
rect 246297 270947 246363 270950
rect 156781 270466 156847 270469
rect 154652 270464 156847 270466
rect 154652 270408 156786 270464
rect 156842 270408 156847 270464
rect 154652 270406 156847 270408
rect 156781 270403 156847 270406
rect 197353 270194 197419 270197
rect 245653 270194 245719 270197
rect 197353 270192 200284 270194
rect 197353 270136 197358 270192
rect 197414 270136 200284 270192
rect 197353 270134 200284 270136
rect 244076 270192 245719 270194
rect 244076 270136 245658 270192
rect 245714 270136 245719 270192
rect 244076 270134 245719 270136
rect 197353 270131 197419 270134
rect 245653 270131 245719 270134
rect 66437 269922 66503 269925
rect 66437 269920 68908 269922
rect 66437 269864 66442 269920
rect 66498 269864 68908 269920
rect 66437 269862 68908 269864
rect 66437 269859 66503 269862
rect 245929 269650 245995 269653
rect 244076 269648 245995 269650
rect 244076 269592 245934 269648
rect 245990 269592 245995 269648
rect 244076 269590 245995 269592
rect 245929 269587 245995 269590
rect 157241 269378 157307 269381
rect 154652 269376 157307 269378
rect 154652 269320 157246 269376
rect 157302 269320 157307 269376
rect 154652 269318 157307 269320
rect 157241 269315 157307 269318
rect 200070 269318 200284 269378
rect 200070 269242 200130 269318
rect 165478 269182 200130 269242
rect 162117 269106 162183 269109
rect 164233 269106 164299 269109
rect 165478 269106 165538 269182
rect 162117 269104 165538 269106
rect 162117 269048 162122 269104
rect 162178 269048 164238 269104
rect 164294 269048 165538 269104
rect 162117 269046 165538 269048
rect 162117 269043 162183 269046
rect 164233 269043 164299 269046
rect 67766 268772 67772 268836
rect 67836 268834 67842 268836
rect 197353 268834 197419 268837
rect 244457 268834 244523 268837
rect 67836 268774 68908 268834
rect 197353 268832 200284 268834
rect 197353 268776 197358 268832
rect 197414 268776 200284 268832
rect 197353 268774 200284 268776
rect 244076 268832 244523 268834
rect 244076 268776 244462 268832
rect 244518 268776 244523 268832
rect 244076 268774 244523 268776
rect 67836 268772 67842 268774
rect 197353 268771 197419 268774
rect 244457 268771 244523 268774
rect 156505 268290 156571 268293
rect 154652 268288 156571 268290
rect 154652 268232 156510 268288
rect 156566 268232 156571 268288
rect 154652 268230 156571 268232
rect 156505 268227 156571 268230
rect 245929 268018 245995 268021
rect 200070 267958 200284 268018
rect 244076 268016 245995 268018
rect 244076 267960 245934 268016
rect 245990 267960 245995 268016
rect 244076 267958 245995 267960
rect 172421 267882 172487 267885
rect 200070 267882 200130 267958
rect 245929 267955 245995 267958
rect 315941 267882 316007 267885
rect 316166 267882 316172 267884
rect 172421 267880 200130 267882
rect 172421 267824 172426 267880
rect 172482 267824 200130 267880
rect 172421 267822 200130 267824
rect 315896 267880 316172 267882
rect 315896 267824 315946 267880
rect 316002 267824 316172 267880
rect 315896 267822 316172 267824
rect 172421 267819 172487 267822
rect 315941 267819 316007 267822
rect 316166 267820 316172 267822
rect 316236 267820 316242 267884
rect 66437 267746 66503 267749
rect 67950 267746 67956 267748
rect 66437 267744 67956 267746
rect 66437 267688 66442 267744
rect 66498 267688 67956 267744
rect 66437 267686 67956 267688
rect 66437 267683 66503 267686
rect 67950 267684 67956 267686
rect 68020 267746 68026 267748
rect 315941 267746 316007 267749
rect 316166 267746 316172 267748
rect 68020 267686 68908 267746
rect 315896 267744 316172 267746
rect 315896 267688 315946 267744
rect 316002 267688 316172 267744
rect 315896 267686 316172 267688
rect 68020 267684 68026 267686
rect 315941 267683 316007 267686
rect 316166 267684 316172 267686
rect 316236 267684 316242 267748
rect 157241 267474 157307 267477
rect 246021 267474 246087 267477
rect 154652 267472 157307 267474
rect 154652 267416 157246 267472
rect 157302 267416 157307 267472
rect 154652 267414 157307 267416
rect 244076 267472 246087 267474
rect 244076 267416 246026 267472
rect 246082 267416 246087 267472
rect 244076 267414 246087 267416
rect 157241 267411 157307 267414
rect 246021 267411 246087 267414
rect -960 267202 480 267292
rect 3417 267202 3483 267205
rect -960 267200 3483 267202
rect -960 267144 3422 267200
rect 3478 267144 3483 267200
rect -960 267142 3483 267144
rect -960 267052 480 267142
rect 3417 267139 3483 267142
rect 197118 267140 197124 267204
rect 197188 267202 197194 267204
rect 197188 267142 200284 267202
rect 197188 267140 197194 267142
rect 244222 267004 244228 267068
rect 244292 267066 244298 267068
rect 328453 267066 328519 267069
rect 244292 267064 328519 267066
rect 244292 267008 328458 267064
rect 328514 267008 328519 267064
rect 244292 267006 328519 267008
rect 244292 267004 244298 267006
rect 328453 267003 328519 267006
rect 66662 266868 66668 266932
rect 66732 266930 66738 266932
rect 66732 266870 68908 266930
rect 66732 266868 66738 266870
rect 197353 266658 197419 266661
rect 245929 266658 245995 266661
rect 197353 266656 200284 266658
rect 197353 266600 197358 266656
rect 197414 266600 200284 266656
rect 197353 266598 200284 266600
rect 244076 266656 245995 266658
rect 244076 266600 245934 266656
rect 245990 266600 245995 266656
rect 244076 266598 245995 266600
rect 197353 266595 197419 266598
rect 245929 266595 245995 266598
rect 188337 266386 188403 266389
rect 154652 266384 188403 266386
rect 154652 266328 188342 266384
rect 188398 266328 188403 266384
rect 154652 266326 188403 266328
rect 188337 266323 188403 266326
rect 66805 265842 66871 265845
rect 197353 265842 197419 265845
rect 245837 265842 245903 265845
rect 66805 265840 68908 265842
rect 66805 265784 66810 265840
rect 66866 265784 68908 265840
rect 66805 265782 68908 265784
rect 197353 265840 200284 265842
rect 197353 265784 197358 265840
rect 197414 265784 200284 265840
rect 197353 265782 200284 265784
rect 244076 265840 245903 265842
rect 244076 265784 245842 265840
rect 245898 265784 245903 265840
rect 244076 265782 245903 265784
rect 66805 265779 66871 265782
rect 197353 265779 197419 265782
rect 245837 265779 245903 265782
rect 157241 265298 157307 265301
rect 154652 265296 157307 265298
rect 154652 265240 157246 265296
rect 157302 265240 157307 265296
rect 154652 265238 157307 265240
rect 157241 265235 157307 265238
rect 199878 265236 199884 265300
rect 199948 265298 199954 265300
rect 245745 265298 245811 265301
rect 199948 265238 200284 265298
rect 244076 265296 245811 265298
rect 244076 265240 245750 265296
rect 245806 265240 245811 265296
rect 244076 265238 245811 265240
rect 199948 265236 199954 265238
rect 245745 265235 245811 265238
rect 66805 264754 66871 264757
rect 154757 264754 154823 264757
rect 66805 264752 68908 264754
rect 66805 264696 66810 264752
rect 66866 264696 68908 264752
rect 66805 264694 68908 264696
rect 154622 264752 154823 264754
rect 154622 264696 154762 264752
rect 154818 264696 154823 264752
rect 154622 264694 154823 264696
rect 66805 264691 66871 264694
rect 154622 264180 154682 264694
rect 154757 264691 154823 264694
rect 197353 264482 197419 264485
rect 245837 264482 245903 264485
rect 197353 264480 200284 264482
rect 197353 264424 197358 264480
rect 197414 264424 200284 264480
rect 197353 264422 200284 264424
rect 244076 264480 245903 264482
rect 244076 264424 245842 264480
rect 245898 264424 245903 264480
rect 244076 264422 245903 264424
rect 197353 264419 197419 264422
rect 245837 264419 245903 264422
rect 262213 264210 262279 264213
rect 583109 264210 583175 264213
rect 262213 264208 583175 264210
rect 262213 264152 262218 264208
rect 262274 264152 583114 264208
rect 583170 264152 583175 264208
rect 262213 264150 583175 264152
rect 262213 264147 262279 264150
rect 583109 264147 583175 264150
rect 245929 263938 245995 263941
rect 244076 263936 245995 263938
rect 244076 263880 245934 263936
rect 245990 263880 245995 263936
rect 244076 263878 245995 263880
rect 245929 263875 245995 263878
rect 66437 263666 66503 263669
rect 197353 263666 197419 263669
rect 66437 263664 68908 263666
rect 66437 263608 66442 263664
rect 66498 263608 68908 263664
rect 66437 263606 68908 263608
rect 197353 263664 200284 263666
rect 197353 263608 197358 263664
rect 197414 263608 200284 263664
rect 197353 263606 200284 263608
rect 66437 263603 66503 263606
rect 197353 263603 197419 263606
rect 157241 263122 157307 263125
rect 154652 263120 157307 263122
rect 154652 263064 157246 263120
rect 157302 263064 157307 263120
rect 154652 263062 157307 263064
rect 157241 263059 157307 263062
rect 199469 263122 199535 263125
rect 245745 263122 245811 263125
rect 199469 263120 200284 263122
rect 199469 263064 199474 263120
rect 199530 263064 200284 263120
rect 199469 263062 200284 263064
rect 244076 263120 245811 263122
rect 244076 263064 245750 263120
rect 245806 263064 245811 263120
rect 244076 263062 245811 263064
rect 199469 263059 199535 263062
rect 245745 263059 245811 263062
rect 66805 262578 66871 262581
rect 66805 262576 68908 262578
rect 66805 262520 66810 262576
rect 66866 262520 68908 262576
rect 66805 262518 68908 262520
rect 66805 262515 66871 262518
rect 197353 262306 197419 262309
rect 245929 262306 245995 262309
rect 197353 262304 200284 262306
rect 197353 262248 197358 262304
rect 197414 262248 200284 262304
rect 197353 262246 200284 262248
rect 244076 262304 245995 262306
rect 244076 262248 245934 262304
rect 245990 262248 245995 262304
rect 244076 262246 245995 262248
rect 197353 262243 197419 262246
rect 245929 262243 245995 262246
rect 154849 262034 154915 262037
rect 154652 262032 154915 262034
rect 154652 261976 154854 262032
rect 154910 261976 154915 262032
rect 154652 261974 154915 261976
rect 154849 261971 154915 261974
rect 245837 261762 245903 261765
rect 244076 261760 245903 261762
rect 244076 261704 245842 261760
rect 245898 261704 245903 261760
rect 244076 261702 245903 261704
rect 245837 261699 245903 261702
rect 66805 261490 66871 261493
rect 197445 261490 197511 261493
rect 66805 261488 68908 261490
rect 66805 261432 66810 261488
rect 66866 261432 68908 261488
rect 66805 261430 68908 261432
rect 197445 261488 200284 261490
rect 197445 261432 197450 261488
rect 197506 261432 200284 261488
rect 197445 261430 200284 261432
rect 66805 261427 66871 261430
rect 197445 261427 197511 261430
rect 156781 260946 156847 260949
rect 154652 260944 156847 260946
rect 154652 260916 156786 260944
rect 154622 260888 156786 260916
rect 156842 260888 156847 260944
rect 154622 260886 156847 260888
rect 154622 260812 154682 260886
rect 156781 260883 156847 260886
rect 197353 260946 197419 260949
rect 244549 260946 244615 260949
rect 244917 260946 244983 260949
rect 197353 260944 200284 260946
rect 197353 260888 197358 260944
rect 197414 260888 200284 260944
rect 197353 260886 200284 260888
rect 244076 260944 244983 260946
rect 244076 260888 244554 260944
rect 244610 260888 244922 260944
rect 244978 260888 244983 260944
rect 244076 260886 244983 260888
rect 197353 260883 197419 260886
rect 244549 260883 244615 260886
rect 244917 260883 244983 260886
rect 154614 260748 154620 260812
rect 154684 260748 154690 260812
rect 67541 260402 67607 260405
rect 67541 260400 68908 260402
rect 67541 260344 67546 260400
rect 67602 260344 68908 260400
rect 67541 260342 68908 260344
rect 67541 260339 67607 260342
rect 197353 260130 197419 260133
rect 197353 260128 200284 260130
rect 197353 260072 197358 260128
rect 197414 260072 200284 260128
rect 197353 260070 200284 260072
rect 197353 260067 197419 260070
rect 156689 259858 156755 259861
rect 154652 259856 156755 259858
rect 154652 259800 156694 259856
rect 156750 259800 156755 259856
rect 154652 259798 156755 259800
rect 244046 259858 244106 260100
rect 251449 259858 251515 259861
rect 244046 259856 251515 259858
rect 244046 259800 251454 259856
rect 251510 259800 251515 259856
rect 244046 259798 251515 259800
rect 156689 259795 156755 259798
rect 251449 259795 251515 259798
rect 245929 259586 245995 259589
rect 244076 259584 245995 259586
rect 244076 259528 245934 259584
rect 245990 259528 245995 259584
rect 244076 259526 245995 259528
rect 245929 259523 245995 259526
rect 197353 259314 197419 259317
rect 197353 259312 200284 259314
rect 68093 258770 68159 258773
rect 68878 258770 68938 259284
rect 197353 259256 197358 259312
rect 197414 259256 200284 259312
rect 197353 259254 200284 259256
rect 197353 259251 197419 259254
rect 156597 259042 156663 259045
rect 154652 259040 156663 259042
rect 154652 258984 156602 259040
rect 156658 258984 156663 259040
rect 154652 258982 156663 258984
rect 156597 258979 156663 258982
rect 583017 258906 583083 258909
rect 583520 258906 584960 258996
rect 583017 258904 584960 258906
rect 583017 258848 583022 258904
rect 583078 258848 584960 258904
rect 583017 258846 584960 258848
rect 583017 258843 583083 258846
rect 68093 258768 68938 258770
rect 68093 258712 68098 258768
rect 68154 258712 68938 258768
rect 68093 258710 68938 258712
rect 197445 258770 197511 258773
rect 245929 258770 245995 258773
rect 197445 258768 200284 258770
rect 197445 258712 197450 258768
rect 197506 258712 200284 258768
rect 197445 258710 200284 258712
rect 244076 258768 245995 258770
rect 244076 258712 245934 258768
rect 245990 258712 245995 258768
rect 583520 258756 584960 258846
rect 244076 258710 245995 258712
rect 68093 258707 68159 258710
rect 197445 258707 197511 258710
rect 245929 258707 245995 258710
rect 66805 258498 66871 258501
rect 66805 258496 68908 258498
rect 66805 258440 66810 258496
rect 66866 258440 68908 258496
rect 66805 258438 68908 258440
rect 66805 258435 66871 258438
rect 245837 258226 245903 258229
rect 244076 258224 245903 258226
rect 244076 258168 245842 258224
rect 245898 258168 245903 258224
rect 244076 258166 245903 258168
rect 245837 258163 245903 258166
rect 157241 257954 157307 257957
rect 154652 257952 157307 257954
rect 154652 257896 157246 257952
rect 157302 257896 157307 257952
rect 154652 257894 157307 257896
rect 157241 257891 157307 257894
rect 197353 257954 197419 257957
rect 197353 257952 200284 257954
rect 197353 257896 197358 257952
rect 197414 257896 200284 257952
rect 197353 257894 200284 257896
rect 197353 257891 197419 257894
rect 66437 257410 66503 257413
rect 199653 257410 199719 257413
rect 199929 257410 199995 257413
rect 247217 257410 247283 257413
rect 66437 257408 68908 257410
rect 66437 257352 66442 257408
rect 66498 257352 68908 257408
rect 66437 257350 68908 257352
rect 199653 257408 200284 257410
rect 199653 257352 199658 257408
rect 199714 257352 199934 257408
rect 199990 257352 200284 257408
rect 199653 257350 200284 257352
rect 244076 257408 247283 257410
rect 244076 257352 247222 257408
rect 247278 257352 247283 257408
rect 244076 257350 247283 257352
rect 66437 257347 66503 257350
rect 199653 257347 199719 257350
rect 199929 257347 199995 257350
rect 247217 257347 247283 257350
rect 157241 256866 157307 256869
rect 154652 256864 157307 256866
rect 154652 256808 157246 256864
rect 157302 256808 157307 256864
rect 154652 256806 157307 256808
rect 157241 256803 157307 256806
rect 197353 256594 197419 256597
rect 245653 256594 245719 256597
rect 197353 256592 200284 256594
rect 197353 256536 197358 256592
rect 197414 256536 200284 256592
rect 197353 256534 200284 256536
rect 244076 256592 245719 256594
rect 244076 256536 245658 256592
rect 245714 256536 245719 256592
rect 244076 256534 245719 256536
rect 197353 256531 197419 256534
rect 245653 256531 245719 256534
rect 66069 256322 66135 256325
rect 66069 256320 68908 256322
rect 66069 256264 66074 256320
rect 66130 256264 68908 256320
rect 66069 256262 68908 256264
rect 66069 256259 66135 256262
rect 61878 255988 61884 256052
rect 61948 256050 61954 256052
rect 66989 256050 67055 256053
rect 244457 256050 244523 256053
rect 61948 256048 67055 256050
rect 61948 255992 66994 256048
rect 67050 255992 67055 256048
rect 61948 255990 67055 255992
rect 244076 256048 244523 256050
rect 244076 255992 244462 256048
rect 244518 255992 244523 256048
rect 244076 255990 244523 255992
rect 61948 255988 61954 255990
rect 66989 255987 67055 255990
rect 244457 255987 244523 255990
rect 157241 255778 157307 255781
rect 154652 255776 157307 255778
rect 154652 255720 157246 255776
rect 157302 255720 157307 255776
rect 154652 255718 157307 255720
rect 157241 255715 157307 255718
rect 173157 255506 173223 255509
rect 200254 255506 200314 255748
rect 173157 255504 200314 255506
rect 173157 255448 173162 255504
rect 173218 255448 200314 255504
rect 173157 255446 200314 255448
rect 173157 255443 173223 255446
rect 66437 255234 66503 255237
rect 197997 255234 198063 255237
rect 246021 255234 246087 255237
rect 66437 255232 68908 255234
rect 66437 255176 66442 255232
rect 66498 255176 68908 255232
rect 66437 255174 68908 255176
rect 197997 255232 200284 255234
rect 197997 255176 198002 255232
rect 198058 255176 200284 255232
rect 197997 255174 200284 255176
rect 244076 255232 246087 255234
rect 244076 255176 246026 255232
rect 246082 255176 246087 255232
rect 244076 255174 246087 255176
rect 66437 255171 66503 255174
rect 197997 255171 198063 255174
rect 246021 255171 246087 255174
rect 156045 254690 156111 254693
rect 157241 254690 157307 254693
rect 154652 254688 157307 254690
rect 154652 254632 156050 254688
rect 156106 254632 157246 254688
rect 157302 254632 157307 254688
rect 154652 254630 157307 254632
rect 156045 254627 156111 254630
rect 157241 254627 157307 254630
rect 197353 254418 197419 254421
rect 248413 254418 248479 254421
rect 197353 254416 200284 254418
rect 197353 254360 197358 254416
rect 197414 254360 200284 254416
rect 197353 254358 200284 254360
rect 244076 254416 248479 254418
rect 244076 254360 248418 254416
rect 248474 254360 248479 254416
rect 244076 254358 248479 254360
rect 197353 254355 197419 254358
rect 248413 254355 248479 254358
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 69430 254012 69490 254116
rect 69422 253948 69428 254012
rect 69492 253948 69498 254012
rect 245929 253874 245995 253877
rect 244076 253872 245995 253874
rect 244076 253816 245934 253872
rect 245990 253816 245995 253872
rect 244076 253814 245995 253816
rect 245929 253811 245995 253814
rect 157241 253602 157307 253605
rect 154652 253600 157307 253602
rect 154652 253544 157246 253600
rect 157302 253544 157307 253600
rect 154652 253542 157307 253544
rect 157241 253539 157307 253542
rect 197445 253602 197511 253605
rect 197445 253600 200284 253602
rect 197445 253544 197450 253600
rect 197506 253544 200284 253600
rect 197445 253542 200284 253544
rect 197445 253539 197511 253542
rect 156781 253194 156847 253197
rect 170489 253194 170555 253197
rect 156781 253192 170555 253194
rect 156781 253136 156786 253192
rect 156842 253136 170494 253192
rect 170550 253136 170555 253192
rect 156781 253134 170555 253136
rect 156781 253131 156847 253134
rect 170489 253131 170555 253134
rect 66621 253058 66687 253061
rect 200021 253058 200087 253061
rect 245929 253058 245995 253061
rect 66621 253056 68908 253058
rect 66621 253000 66626 253056
rect 66682 253000 68908 253056
rect 66621 252998 68908 253000
rect 200021 253056 200284 253058
rect 200021 253000 200026 253056
rect 200082 253000 200284 253056
rect 200021 252998 200284 253000
rect 244076 253056 245995 253058
rect 244076 253000 245934 253056
rect 245990 253000 245995 253056
rect 244076 252998 245995 253000
rect 66621 252995 66687 252998
rect 200021 252995 200087 252998
rect 245929 252995 245995 252998
rect 156137 252514 156203 252517
rect 154652 252512 156203 252514
rect 154652 252456 156142 252512
rect 156198 252456 156203 252512
rect 154652 252454 156203 252456
rect 156137 252451 156203 252454
rect 197445 252242 197511 252245
rect 246941 252242 247007 252245
rect 197445 252240 200284 252242
rect 197445 252184 197450 252240
rect 197506 252184 200284 252240
rect 197445 252182 200284 252184
rect 244076 252240 247007 252242
rect 244076 252184 246946 252240
rect 247002 252184 247007 252240
rect 244076 252182 247007 252184
rect 197445 252179 197511 252182
rect 246941 252179 247007 252182
rect 67398 251908 67404 251972
rect 67468 251970 67474 251972
rect 67468 251910 68908 251970
rect 67468 251908 67474 251910
rect 197353 251698 197419 251701
rect 245745 251698 245811 251701
rect 197353 251696 200284 251698
rect 197353 251640 197358 251696
rect 197414 251640 200284 251696
rect 197353 251638 200284 251640
rect 244076 251696 245811 251698
rect 244076 251640 245750 251696
rect 245806 251640 245811 251696
rect 244076 251638 245811 251640
rect 197353 251635 197419 251638
rect 245745 251635 245811 251638
rect 157241 251426 157307 251429
rect 154652 251424 157307 251426
rect 154652 251368 157246 251424
rect 157302 251368 157307 251424
rect 154652 251366 157307 251368
rect 157241 251363 157307 251366
rect 67909 250882 67975 250885
rect 197445 250882 197511 250885
rect 245745 250882 245811 250885
rect 67909 250880 68908 250882
rect 67909 250824 67914 250880
rect 67970 250824 68908 250880
rect 67909 250822 68908 250824
rect 197445 250880 200284 250882
rect 197445 250824 197450 250880
rect 197506 250824 200284 250880
rect 197445 250822 200284 250824
rect 244076 250880 245811 250882
rect 244076 250824 245750 250880
rect 245806 250824 245811 250880
rect 244076 250822 245811 250824
rect 67909 250819 67975 250822
rect 197445 250819 197511 250822
rect 245745 250819 245811 250822
rect 157241 250610 157307 250613
rect 154652 250608 157307 250610
rect 154652 250552 157246 250608
rect 157302 250552 157307 250608
rect 154652 250550 157307 250552
rect 157241 250547 157307 250550
rect 244365 250338 244431 250341
rect 244076 250336 244431 250338
rect 244076 250280 244370 250336
rect 244426 250280 244431 250336
rect 244076 250278 244431 250280
rect 244365 250275 244431 250278
rect 67725 250066 67791 250069
rect 197353 250066 197419 250069
rect 67725 250064 68908 250066
rect 67725 250008 67730 250064
rect 67786 250008 68908 250064
rect 67725 250006 68908 250008
rect 197353 250064 200284 250066
rect 197353 250008 197358 250064
rect 197414 250008 200284 250064
rect 197353 250006 200284 250008
rect 67725 250003 67791 250006
rect 197353 250003 197419 250006
rect 157149 249522 157215 249525
rect 154652 249520 157215 249522
rect 154652 249464 157154 249520
rect 157210 249464 157215 249520
rect 154652 249462 157215 249464
rect 157149 249459 157215 249462
rect 197445 249522 197511 249525
rect 245929 249522 245995 249525
rect 197445 249520 200284 249522
rect 197445 249464 197450 249520
rect 197506 249464 200284 249520
rect 197445 249462 200284 249464
rect 244076 249520 245995 249522
rect 244076 249464 245934 249520
rect 245990 249464 245995 249520
rect 244076 249462 245995 249464
rect 197445 249459 197511 249462
rect 245929 249459 245995 249462
rect 181529 249114 181595 249117
rect 197169 249114 197235 249117
rect 181529 249112 200314 249114
rect 181529 249056 181534 249112
rect 181590 249056 197174 249112
rect 197230 249056 200314 249112
rect 181529 249054 200314 249056
rect 181529 249051 181595 249054
rect 197169 249051 197235 249054
rect 66805 248978 66871 248981
rect 66805 248976 68908 248978
rect 66805 248920 66810 248976
rect 66866 248920 68908 248976
rect 66805 248918 68908 248920
rect 66805 248915 66871 248918
rect 200254 248676 200314 249054
rect 244917 248706 244983 248709
rect 244076 248704 244983 248706
rect 244076 248648 244922 248704
rect 244978 248648 244983 248704
rect 244076 248646 244983 248648
rect 244917 248643 244983 248646
rect 200021 248570 200087 248573
rect 199976 248568 200130 248570
rect 199976 248512 200026 248568
rect 200082 248512 200130 248568
rect 199976 248510 200130 248512
rect 200021 248507 200130 248510
rect 157241 248434 157307 248437
rect 154652 248432 157307 248434
rect 154652 248376 157246 248432
rect 157302 248376 157307 248432
rect 154652 248374 157307 248376
rect 157241 248371 157307 248374
rect 192937 248434 193003 248437
rect 200070 248436 200130 248507
rect 315941 248436 316007 248437
rect 199510 248434 199516 248436
rect 192937 248432 199516 248434
rect 192937 248376 192942 248432
rect 192998 248376 199516 248432
rect 192937 248374 199516 248376
rect 192937 248371 193003 248374
rect 199510 248372 199516 248374
rect 199580 248372 199586 248436
rect 200062 248372 200068 248436
rect 200132 248372 200138 248436
rect 315941 248434 315988 248436
rect 315896 248432 315988 248434
rect 316052 248434 316058 248436
rect 315896 248376 315946 248432
rect 315896 248374 315988 248376
rect 315941 248372 315988 248374
rect 316052 248374 316134 248434
rect 316052 248372 316058 248374
rect 315941 248371 316007 248372
rect 315941 248298 316007 248301
rect 316166 248298 316172 248300
rect 315896 248296 316172 248298
rect 315896 248240 315946 248296
rect 316002 248240 316172 248296
rect 315896 248238 316172 248240
rect 315941 248235 316007 248238
rect 316166 248236 316172 248238
rect 316236 248236 316242 248300
rect 245929 248162 245995 248165
rect 244076 248160 245995 248162
rect 244076 248104 245934 248160
rect 245990 248104 245995 248160
rect 244076 248102 245995 248104
rect 245929 248099 245995 248102
rect 66805 247890 66871 247893
rect 197353 247890 197419 247893
rect 66805 247888 68908 247890
rect 66805 247832 66810 247888
rect 66866 247832 68908 247888
rect 66805 247830 68908 247832
rect 197353 247888 200284 247890
rect 197353 247832 197358 247888
rect 197414 247832 200284 247888
rect 197353 247830 200284 247832
rect 66805 247827 66871 247830
rect 197353 247827 197419 247830
rect 186957 247618 187023 247621
rect 200062 247618 200068 247620
rect 186957 247616 200068 247618
rect 186957 247560 186962 247616
rect 187018 247560 200068 247616
rect 186957 247558 200068 247560
rect 186957 247555 187023 247558
rect 200062 247556 200068 247558
rect 200132 247556 200138 247620
rect 157241 247346 157307 247349
rect 154652 247344 157307 247346
rect 154652 247288 157246 247344
rect 157302 247288 157307 247344
rect 154652 247286 157307 247288
rect 157241 247283 157307 247286
rect 196709 247346 196775 247349
rect 244365 247346 244431 247349
rect 196709 247344 200284 247346
rect 196709 247288 196714 247344
rect 196770 247288 200284 247344
rect 196709 247286 200284 247288
rect 244076 247344 244431 247346
rect 244076 247288 244370 247344
rect 244426 247288 244431 247344
rect 244076 247286 244431 247288
rect 196709 247283 196775 247286
rect 244365 247283 244431 247286
rect 165521 247074 165587 247077
rect 170949 247074 171015 247077
rect 171133 247074 171199 247077
rect 165521 247072 171199 247074
rect 165521 247016 165526 247072
rect 165582 247016 170954 247072
rect 171010 247016 171138 247072
rect 171194 247016 171199 247072
rect 165521 247014 171199 247016
rect 165521 247011 165587 247014
rect 170949 247011 171015 247014
rect 171133 247011 171199 247014
rect 67265 246802 67331 246805
rect 67265 246800 68908 246802
rect 67265 246744 67270 246800
rect 67326 246744 68908 246800
rect 67265 246742 68908 246744
rect 67265 246739 67331 246742
rect 197353 246530 197419 246533
rect 197353 246528 200284 246530
rect 197353 246472 197358 246528
rect 197414 246472 200284 246528
rect 197353 246470 200284 246472
rect 197353 246467 197419 246470
rect 157241 246258 157307 246261
rect 243494 246260 243554 246500
rect 154652 246256 157307 246258
rect 154652 246200 157246 246256
rect 157302 246200 157307 246256
rect 154652 246198 157307 246200
rect 157241 246195 157307 246198
rect 243486 246196 243492 246260
rect 243556 246196 243562 246260
rect 69422 245924 69428 245988
rect 69492 245924 69498 245988
rect 197445 245986 197511 245989
rect 246389 245986 246455 245989
rect 197445 245984 200284 245986
rect 197445 245928 197450 245984
rect 197506 245928 200284 245984
rect 197445 245926 200284 245928
rect 244076 245984 246455 245986
rect 244076 245928 246394 245984
rect 246450 245928 246455 245984
rect 244076 245926 246455 245928
rect 69430 245684 69490 245924
rect 197445 245923 197511 245926
rect 246389 245923 246455 245926
rect 155585 245850 155651 245853
rect 199469 245850 199535 245853
rect 155585 245848 199535 245850
rect 155585 245792 155590 245848
rect 155646 245792 199474 245848
rect 199530 245792 199535 245848
rect 155585 245790 199535 245792
rect 155585 245787 155651 245790
rect 199469 245787 199535 245790
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 156597 245170 156663 245173
rect 154652 245168 156663 245170
rect 154652 245112 156602 245168
rect 156658 245112 156663 245168
rect 154652 245110 156663 245112
rect 156597 245107 156663 245110
rect 197445 245170 197511 245173
rect 245837 245170 245903 245173
rect 197445 245168 200284 245170
rect 197445 245112 197450 245168
rect 197506 245112 200284 245168
rect 197445 245110 200284 245112
rect 244076 245168 245903 245170
rect 244076 245112 245842 245168
rect 245898 245112 245903 245168
rect 244076 245110 245903 245112
rect 197445 245107 197511 245110
rect 245837 245107 245903 245110
rect 246297 244898 246363 244901
rect 298134 244898 298140 244900
rect 246297 244896 298140 244898
rect 246297 244840 246302 244896
rect 246358 244840 298140 244896
rect 246297 244838 298140 244840
rect 246297 244835 246363 244838
rect 298134 244836 298140 244838
rect 298204 244836 298210 244900
rect 67173 244626 67239 244629
rect 67173 244624 69276 244626
rect 67173 244568 67178 244624
rect 67234 244596 69276 244624
rect 67234 244568 69306 244596
rect 67173 244566 69306 244568
rect 67173 244563 67239 244566
rect 69246 244356 69306 244566
rect 154246 244564 154252 244628
rect 154316 244626 154322 244628
rect 199837 244626 199903 244629
rect 245929 244626 245995 244629
rect 154316 244624 199903 244626
rect 154316 244568 199842 244624
rect 199898 244568 199903 244624
rect 154316 244566 199903 244568
rect 244076 244624 245995 244626
rect 244076 244568 245934 244624
rect 245990 244568 245995 244624
rect 244076 244566 245995 244568
rect 154316 244564 154322 244566
rect 199837 244563 199903 244566
rect 245929 244563 245995 244566
rect 69238 244292 69244 244356
rect 69308 244292 69314 244356
rect 197353 244354 197419 244357
rect 197353 244352 200284 244354
rect 197353 244296 197358 244352
rect 197414 244296 200284 244352
rect 197353 244294 200284 244296
rect 197353 244291 197419 244294
rect 157241 244082 157307 244085
rect 154652 244080 157307 244082
rect 154652 244024 157246 244080
rect 157302 244024 157307 244080
rect 154652 244022 157307 244024
rect 157241 244019 157307 244022
rect 196709 243810 196775 243813
rect 246389 243810 246455 243813
rect 196709 243808 200284 243810
rect 196709 243752 196714 243808
rect 196770 243752 200284 243808
rect 196709 243750 200284 243752
rect 244076 243808 246455 243810
rect 244076 243752 246394 243808
rect 246450 243752 246455 243808
rect 244076 243750 246455 243752
rect 196709 243747 196775 243750
rect 246389 243747 246455 243750
rect 67766 243476 67772 243540
rect 67836 243538 67842 243540
rect 67836 243478 68908 243538
rect 67836 243476 67842 243478
rect 155166 243476 155172 243540
rect 155236 243538 155242 243540
rect 159449 243538 159515 243541
rect 155236 243536 159515 243538
rect 155236 243480 159454 243536
rect 159510 243480 159515 243536
rect 155236 243478 159515 243480
rect 155236 243476 155242 243478
rect 159449 243475 159515 243478
rect 159725 243130 159791 243133
rect 192477 243130 192543 243133
rect 159725 243128 192543 243130
rect 159725 243072 159730 243128
rect 159786 243072 192482 243128
rect 192538 243072 192543 243128
rect 159725 243070 192543 243072
rect 159725 243067 159791 243070
rect 192477 243067 192543 243070
rect 156137 242994 156203 242997
rect 154652 242992 156203 242994
rect 154652 242936 156142 242992
rect 156198 242936 156203 242992
rect 154652 242934 156203 242936
rect 156137 242931 156203 242934
rect 189073 242994 189139 242997
rect 245878 242994 245884 242996
rect 189073 242992 200284 242994
rect 189073 242936 189078 242992
rect 189134 242936 200284 242992
rect 189073 242934 200284 242936
rect 244076 242934 245884 242994
rect 189073 242931 189139 242934
rect 245878 242932 245884 242934
rect 245948 242932 245954 242996
rect 246297 242450 246363 242453
rect 244076 242448 246363 242450
rect 69430 241906 69490 242420
rect 244076 242392 246302 242448
rect 246358 242392 246363 242448
rect 244076 242390 246363 242392
rect 246297 242387 246363 242390
rect 156781 242178 156847 242181
rect 154652 242176 156847 242178
rect 154652 242120 156786 242176
rect 156842 242120 156847 242176
rect 154652 242118 156847 242120
rect 156781 242115 156847 242118
rect 197905 242178 197971 242181
rect 197905 242176 200284 242178
rect 197905 242120 197910 242176
rect 197966 242120 200284 242176
rect 197905 242118 200284 242120
rect 197905 242115 197971 242118
rect 135989 242044 136055 242045
rect 135989 242042 136036 242044
rect 135944 242040 136036 242042
rect 135944 241984 135994 242040
rect 135944 241982 136036 241984
rect 135989 241980 136036 241982
rect 136100 241980 136106 242044
rect 138054 241980 138060 242044
rect 138124 242042 138130 242044
rect 138197 242042 138263 242045
rect 138124 242040 138263 242042
rect 138124 241984 138202 242040
rect 138258 241984 138263 242040
rect 138124 241982 138263 241984
rect 138124 241980 138130 241982
rect 135989 241979 136055 241980
rect 138197 241979 138263 241982
rect 150249 242042 150315 242045
rect 164969 242042 165035 242045
rect 150249 242040 165035 242042
rect 150249 241984 150254 242040
rect 150310 241984 164974 242040
rect 165030 241984 165035 242040
rect 150249 241982 165035 241984
rect 150249 241979 150315 241982
rect 164969 241979 165035 241982
rect 69749 241906 69815 241909
rect 69430 241904 69815 241906
rect 69430 241848 69754 241904
rect 69810 241848 69815 241904
rect 69430 241846 69815 241848
rect 69749 241843 69815 241846
rect 151854 241844 151860 241908
rect 151924 241906 151930 241908
rect 152549 241906 152615 241909
rect 151924 241904 152615 241906
rect 151924 241848 152554 241904
rect 152610 241848 152615 241904
rect 151924 241846 152615 241848
rect 151924 241844 151930 241846
rect 152549 241843 152615 241846
rect 69238 241708 69244 241772
rect 69308 241770 69314 241772
rect 69657 241770 69723 241773
rect 69308 241768 69723 241770
rect 69308 241712 69662 241768
rect 69718 241712 69723 241768
rect 69308 241710 69723 241712
rect 69308 241708 69314 241710
rect 69657 241707 69723 241710
rect 155493 241770 155559 241773
rect 172513 241772 172579 241773
rect 172462 241770 172468 241772
rect 155493 241768 172468 241770
rect 172532 241770 172579 241772
rect 172532 241768 172660 241770
rect 155493 241712 155498 241768
rect 155554 241712 172468 241768
rect 172574 241712 172660 241768
rect 155493 241710 172468 241712
rect 155493 241707 155559 241710
rect 172462 241708 172468 241710
rect 172532 241710 172660 241712
rect 172532 241708 172579 241710
rect 172513 241707 172579 241708
rect 195329 241634 195395 241637
rect 195329 241632 200284 241634
rect 195329 241576 195334 241632
rect 195390 241576 200284 241632
rect 195329 241574 200284 241576
rect 195329 241571 195395 241574
rect 57789 241498 57855 241501
rect 82951 241498 83017 241501
rect 84101 241498 84167 241501
rect 148133 241500 148199 241501
rect 148133 241498 148180 241500
rect 57789 241496 84167 241498
rect 57789 241440 57794 241496
rect 57850 241440 82956 241496
rect 83012 241440 84106 241496
rect 84162 241440 84167 241496
rect 57789 241438 84167 241440
rect 148088 241496 148180 241498
rect 148088 241440 148138 241496
rect 148088 241438 148180 241440
rect 57789 241435 57855 241438
rect 82951 241435 83017 241438
rect 84101 241435 84167 241438
rect 148133 241436 148180 241438
rect 148244 241436 148250 241500
rect 150663 241498 150729 241501
rect 170397 241498 170463 241501
rect 150663 241496 170463 241498
rect 150663 241440 150668 241496
rect 150724 241440 170402 241496
rect 170458 241440 170463 241496
rect 150663 241438 170463 241440
rect 148133 241435 148199 241436
rect 150663 241435 150729 241438
rect 170397 241435 170463 241438
rect 193949 241498 194015 241501
rect 194501 241498 194567 241501
rect 193949 241496 194567 241498
rect 193949 241440 193954 241496
rect 194010 241440 194506 241496
rect 194562 241440 194567 241496
rect 193949 241438 194567 241440
rect 193949 241435 194015 241438
rect 194501 241435 194567 241438
rect 195830 241436 195836 241500
rect 195900 241498 195906 241500
rect 197997 241498 198063 241501
rect 195900 241496 198063 241498
rect 195900 241440 198002 241496
rect 198058 241440 198063 241496
rect 195900 241438 198063 241440
rect 195900 241436 195906 241438
rect 197997 241435 198063 241438
rect 244046 241365 244106 241604
rect 67173 241362 67239 241365
rect 67398 241362 67404 241364
rect 67173 241360 67404 241362
rect 67173 241304 67178 241360
rect 67234 241304 67404 241360
rect 67173 241302 67404 241304
rect 67173 241299 67239 241302
rect 67398 241300 67404 241302
rect 67468 241300 67474 241364
rect 243997 241360 244106 241365
rect 243997 241304 244002 241360
rect 244058 241304 244106 241360
rect 243997 241302 244106 241304
rect 243997 241299 244063 241302
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 245745 240818 245811 240821
rect 244076 240816 245811 240818
rect 195830 240682 195836 240684
rect 180750 240622 195836 240682
rect 148133 240546 148199 240549
rect 180750 240546 180810 240622
rect 195830 240620 195836 240622
rect 195900 240620 195906 240684
rect 148133 240544 180810 240546
rect 148133 240488 148138 240544
rect 148194 240488 180810 240544
rect 148133 240486 180810 240488
rect 194501 240546 194567 240549
rect 200254 240546 200314 240788
rect 244076 240760 245750 240816
rect 245806 240760 245811 240816
rect 244076 240758 245811 240760
rect 245745 240755 245811 240758
rect 194501 240544 200314 240546
rect 194501 240488 194506 240544
rect 194562 240488 200314 240544
rect 194501 240486 200314 240488
rect 148133 240483 148199 240486
rect 194501 240483 194567 240486
rect 71681 240410 71747 240413
rect 199929 240410 199995 240413
rect 71681 240408 199995 240410
rect 71681 240352 71686 240408
rect 71742 240352 199934 240408
rect 199990 240352 199995 240408
rect 71681 240350 199995 240352
rect 71681 240347 71747 240350
rect 199929 240347 199995 240350
rect 199878 240212 199884 240276
rect 199948 240274 199954 240276
rect 200113 240274 200179 240277
rect 245694 240274 245700 240276
rect 199948 240272 200179 240274
rect 199948 240216 200118 240272
rect 200174 240216 200179 240272
rect 199948 240214 200179 240216
rect 244076 240214 245700 240274
rect 199948 240212 199954 240214
rect 200113 240211 200179 240214
rect 245694 240212 245700 240214
rect 245764 240212 245770 240276
rect 199837 240138 199903 240141
rect 200573 240138 200639 240141
rect 199837 240136 200639 240138
rect 199837 240080 199842 240136
rect 199898 240080 200578 240136
rect 200634 240080 200639 240136
rect 199837 240078 200639 240080
rect 199837 240075 199903 240078
rect 200573 240075 200639 240078
rect 224902 240076 224908 240140
rect 224972 240138 224978 240140
rect 225229 240138 225295 240141
rect 224972 240136 225295 240138
rect 224972 240080 225234 240136
rect 225290 240080 225295 240136
rect 224972 240078 225295 240080
rect 224972 240076 224978 240078
rect 225229 240075 225295 240078
rect 227846 240076 227852 240140
rect 227916 240138 227922 240140
rect 228173 240138 228239 240141
rect 231945 240140 232011 240141
rect 227916 240136 228239 240138
rect 227916 240080 228178 240136
rect 228234 240080 228239 240136
rect 227916 240078 228239 240080
rect 227916 240076 227922 240078
rect 228173 240075 228239 240078
rect 231894 240076 231900 240140
rect 231964 240138 232011 240140
rect 231964 240136 232056 240138
rect 232006 240080 232056 240136
rect 231964 240078 232056 240080
rect 231964 240076 232011 240078
rect 237414 240076 237420 240140
rect 237484 240138 237490 240140
rect 237925 240138 237991 240141
rect 252553 240138 252619 240141
rect 580165 240138 580231 240141
rect 237484 240136 237991 240138
rect 237484 240080 237930 240136
rect 237986 240080 237991 240136
rect 237484 240078 237991 240080
rect 237484 240076 237490 240078
rect 231945 240075 232011 240076
rect 237925 240075 237991 240078
rect 248370 240136 580231 240138
rect 248370 240080 252558 240136
rect 252614 240080 580170 240136
rect 580226 240080 580231 240136
rect 248370 240078 580231 240080
rect 126145 240002 126211 240005
rect 228725 240002 228791 240005
rect 232681 240002 232747 240005
rect 126145 240000 232747 240002
rect 126145 239944 126150 240000
rect 126206 239944 228730 240000
rect 228786 239944 232686 240000
rect 232742 239944 232747 240000
rect 126145 239942 232747 239944
rect 126145 239939 126211 239942
rect 228725 239939 228791 239942
rect 232681 239939 232747 239942
rect 239213 240002 239279 240005
rect 248370 240002 248430 240078
rect 252553 240075 252619 240078
rect 580165 240075 580231 240078
rect 239213 240000 248430 240002
rect 239213 239944 239218 240000
rect 239274 239944 248430 240000
rect 239213 239942 248430 239944
rect 239213 239939 239279 239942
rect 117221 239866 117287 239869
rect 224309 239866 224375 239869
rect 117221 239864 224375 239866
rect 117221 239808 117226 239864
rect 117282 239808 224314 239864
rect 224370 239808 224375 239864
rect 117221 239806 224375 239808
rect 117221 239803 117287 239806
rect 224309 239803 224375 239806
rect 50889 239594 50955 239597
rect 74441 239594 74507 239597
rect 50889 239592 74507 239594
rect 50889 239536 50894 239592
rect 50950 239536 74446 239592
rect 74502 239536 74507 239592
rect 50889 239534 74507 239536
rect 50889 239531 50955 239534
rect 74441 239531 74507 239534
rect 232497 239594 232563 239597
rect 246021 239594 246087 239597
rect 232497 239592 246087 239594
rect 232497 239536 232502 239592
rect 232558 239536 246026 239592
rect 246082 239536 246087 239592
rect 232497 239534 246087 239536
rect 232497 239531 232563 239534
rect 246021 239531 246087 239534
rect 43989 239458 44055 239461
rect 77201 239458 77267 239461
rect 43989 239456 77267 239458
rect 43989 239400 43994 239456
rect 44050 239400 77206 239456
rect 77262 239400 77267 239456
rect 43989 239398 77267 239400
rect 43989 239395 44055 239398
rect 77201 239395 77267 239398
rect 84745 239458 84811 239461
rect 106917 239458 106983 239461
rect 84745 239456 106983 239458
rect 84745 239400 84750 239456
rect 84806 239400 106922 239456
rect 106978 239400 106983 239456
rect 84745 239398 106983 239400
rect 84745 239395 84811 239398
rect 106917 239395 106983 239398
rect 112529 239458 112595 239461
rect 220813 239458 220879 239461
rect 112529 239456 220879 239458
rect 112529 239400 112534 239456
rect 112590 239400 220818 239456
rect 220874 239400 220879 239456
rect 112529 239398 220879 239400
rect 112529 239395 112595 239398
rect 220813 239395 220879 239398
rect 224309 239458 224375 239461
rect 242249 239458 242315 239461
rect 224309 239456 242315 239458
rect 224309 239400 224314 239456
rect 224370 239400 242254 239456
rect 242310 239400 242315 239456
rect 224309 239398 242315 239400
rect 224309 239395 224375 239398
rect 242249 239395 242315 239398
rect 315941 238780 316007 238781
rect 315941 238778 315988 238780
rect 315896 238776 315988 238778
rect 316052 238778 316058 238780
rect 315896 238720 315946 238776
rect 315896 238718 315988 238720
rect 315941 238716 315988 238718
rect 316052 238718 316134 238778
rect 316052 238716 316058 238718
rect 315941 238715 316007 238716
rect 70301 238642 70367 238645
rect 200205 238642 200271 238645
rect 70301 238640 200271 238642
rect 70301 238584 70306 238640
rect 70362 238584 200210 238640
rect 200266 238584 200271 238640
rect 70301 238582 200271 238584
rect 70301 238579 70367 238582
rect 200205 238579 200271 238582
rect 202045 238642 202111 238645
rect 203006 238642 203012 238644
rect 202045 238640 203012 238642
rect 202045 238584 202050 238640
rect 202106 238584 203012 238640
rect 202045 238582 203012 238584
rect 202045 238579 202111 238582
rect 203006 238580 203012 238582
rect 203076 238580 203082 238644
rect 212574 238580 212580 238644
rect 212644 238642 212650 238644
rect 213637 238642 213703 238645
rect 212644 238640 213703 238642
rect 212644 238584 213642 238640
rect 213698 238584 213703 238640
rect 212644 238582 213703 238584
rect 212644 238580 212650 238582
rect 213637 238579 213703 238582
rect 222326 238580 222332 238644
rect 222396 238642 222402 238644
rect 223389 238642 223455 238645
rect 222396 238640 223455 238642
rect 222396 238584 223394 238640
rect 223450 238584 223455 238640
rect 222396 238582 223455 238584
rect 222396 238580 222402 238582
rect 223389 238579 223455 238582
rect 227621 238642 227687 238645
rect 229686 238642 229692 238644
rect 227621 238640 229692 238642
rect 227621 238584 227626 238640
rect 227682 238584 229692 238640
rect 227621 238582 229692 238584
rect 227621 238579 227687 238582
rect 229686 238580 229692 238582
rect 229756 238580 229762 238644
rect 233734 238580 233740 238644
rect 233804 238642 233810 238644
rect 236453 238642 236519 238645
rect 233804 238640 236519 238642
rect 233804 238584 236458 238640
rect 236514 238584 236519 238640
rect 233804 238582 236519 238584
rect 233804 238580 233810 238582
rect 236453 238579 236519 238582
rect 241278 238580 241284 238644
rect 241348 238642 241354 238644
rect 241789 238642 241855 238645
rect 315941 238644 316007 238645
rect 315941 238642 315988 238644
rect 241348 238640 241855 238642
rect 241348 238584 241794 238640
rect 241850 238584 241855 238640
rect 241348 238582 241855 238584
rect 315896 238640 315988 238642
rect 316052 238642 316058 238644
rect 315896 238584 315946 238640
rect 315896 238582 315988 238584
rect 241348 238580 241354 238582
rect 241789 238579 241855 238582
rect 315941 238580 315988 238582
rect 316052 238582 316134 238642
rect 316052 238580 316058 238582
rect 315941 238579 316007 238580
rect 73153 238506 73219 238509
rect 202229 238506 202295 238509
rect 73153 238504 202295 238506
rect 73153 238448 73158 238504
rect 73214 238448 202234 238504
rect 202290 238448 202295 238504
rect 73153 238446 202295 238448
rect 73153 238443 73219 238446
rect 202229 238443 202295 238446
rect 218646 238444 218652 238508
rect 218716 238506 218722 238508
rect 232589 238506 232655 238509
rect 218716 238504 232655 238506
rect 218716 238448 232594 238504
rect 232650 238448 232655 238504
rect 218716 238446 232655 238448
rect 218716 238444 218722 238446
rect 232589 238443 232655 238446
rect 235349 238506 235415 238509
rect 259453 238506 259519 238509
rect 235349 238504 259519 238506
rect 235349 238448 235354 238504
rect 235410 238448 259458 238504
rect 259514 238448 259519 238504
rect 235349 238446 259519 238448
rect 235349 238443 235415 238446
rect 259453 238443 259519 238446
rect 124305 238370 124371 238373
rect 148133 238370 148199 238373
rect 124305 238368 148199 238370
rect 124305 238312 124310 238368
rect 124366 238312 148138 238368
rect 148194 238312 148199 238368
rect 124305 238310 148199 238312
rect 124305 238307 124371 238310
rect 148133 238307 148199 238310
rect 242157 238370 242223 238373
rect 252645 238370 252711 238373
rect 242157 238368 252711 238370
rect 242157 238312 242162 238368
rect 242218 238312 252650 238368
rect 252706 238312 252711 238368
rect 242157 238310 252711 238312
rect 242157 238307 242223 238310
rect 252645 238307 252711 238310
rect 230565 238234 230631 238237
rect 230974 238234 230980 238236
rect 230565 238232 230980 238234
rect 230565 238176 230570 238232
rect 230626 238176 230980 238232
rect 230565 238174 230980 238176
rect 230565 238171 230631 238174
rect 230974 238172 230980 238174
rect 231044 238234 231050 238236
rect 287697 238234 287763 238237
rect 231044 238232 287763 238234
rect 231044 238176 287702 238232
rect 287758 238176 287763 238232
rect 231044 238174 287763 238176
rect 231044 238172 231050 238174
rect 287697 238171 287763 238174
rect 218053 238098 218119 238101
rect 223614 238098 223620 238100
rect 218053 238096 223620 238098
rect 218053 238040 218058 238096
rect 218114 238040 223620 238096
rect 218053 238038 223620 238040
rect 218053 238035 218119 238038
rect 223614 238036 223620 238038
rect 223684 238036 223690 238100
rect 60457 237962 60523 237965
rect 73797 237962 73863 237965
rect 60457 237960 73863 237962
rect 60457 237904 60462 237960
rect 60518 237904 73802 237960
rect 73858 237904 73863 237960
rect 60457 237902 73863 237904
rect 60457 237899 60523 237902
rect 73797 237899 73863 237902
rect 200297 237962 200363 237965
rect 224769 237962 224835 237965
rect 200297 237960 224835 237962
rect 200297 237904 200302 237960
rect 200358 237904 224774 237960
rect 224830 237904 224835 237960
rect 200297 237902 224835 237904
rect 200297 237899 200363 237902
rect 224769 237899 224835 237902
rect 259453 237962 259519 237965
rect 582833 237962 582899 237965
rect 259453 237960 582899 237962
rect 259453 237904 259458 237960
rect 259514 237904 582838 237960
rect 582894 237904 582899 237960
rect 259453 237902 582899 237904
rect 259453 237899 259519 237902
rect 582833 237899 582899 237902
rect 147673 237690 147739 237693
rect 152457 237690 152523 237693
rect 147673 237688 152523 237690
rect 147673 237632 147678 237688
rect 147734 237632 152462 237688
rect 152518 237632 152523 237688
rect 147673 237630 152523 237632
rect 147673 237627 147739 237630
rect 152457 237627 152523 237630
rect 167637 237418 167703 237421
rect 168465 237418 168531 237421
rect 167637 237416 168531 237418
rect 167637 237360 167642 237416
rect 167698 237360 168470 237416
rect 168526 237360 168531 237416
rect 167637 237358 168531 237360
rect 167637 237355 167703 237358
rect 168465 237355 168531 237358
rect 200573 237418 200639 237421
rect 201401 237418 201467 237421
rect 200573 237416 201467 237418
rect 200573 237360 200578 237416
rect 200634 237360 201406 237416
rect 201462 237360 201467 237416
rect 200573 237358 201467 237360
rect 200573 237355 200639 237358
rect 201401 237355 201467 237358
rect 209037 237418 209103 237421
rect 211245 237418 211311 237421
rect 209037 237416 211311 237418
rect 209037 237360 209042 237416
rect 209098 237360 211250 237416
rect 211306 237360 211311 237416
rect 209037 237358 211311 237360
rect 209037 237355 209103 237358
rect 211245 237355 211311 237358
rect 212574 237356 212580 237420
rect 212644 237418 212650 237420
rect 213085 237418 213151 237421
rect 212644 237416 213151 237418
rect 212644 237360 213090 237416
rect 213146 237360 213151 237416
rect 212644 237358 213151 237360
rect 212644 237356 212650 237358
rect 213085 237355 213151 237358
rect 237925 237418 237991 237421
rect 238661 237418 238727 237421
rect 237925 237416 238727 237418
rect 237925 237360 237930 237416
rect 237986 237360 238666 237416
rect 238722 237360 238727 237416
rect 237925 237358 238727 237360
rect 237925 237355 237991 237358
rect 238661 237355 238727 237358
rect 252645 237418 252711 237421
rect 253197 237418 253263 237421
rect 252645 237416 253263 237418
rect 252645 237360 252650 237416
rect 252706 237360 253202 237416
rect 253258 237360 253263 237416
rect 252645 237358 253263 237360
rect 252645 237355 252711 237358
rect 253197 237355 253263 237358
rect 103513 237282 103579 237285
rect 137134 237282 137140 237284
rect 103513 237280 137140 237282
rect 103513 237224 103518 237280
rect 103574 237224 137140 237280
rect 103513 237222 137140 237224
rect 103513 237219 103579 237222
rect 137134 237220 137140 237222
rect 137204 237220 137210 237284
rect 180006 237220 180012 237284
rect 180076 237282 180082 237284
rect 204437 237282 204503 237285
rect 180076 237280 204503 237282
rect 180076 237224 204442 237280
rect 204498 237224 204503 237280
rect 180076 237222 204503 237224
rect 180076 237220 180082 237222
rect 204437 237219 204503 237222
rect 207974 237220 207980 237284
rect 208044 237282 208050 237284
rect 214557 237282 214623 237285
rect 208044 237280 214623 237282
rect 208044 237224 214562 237280
rect 214618 237224 214623 237280
rect 208044 237222 214623 237224
rect 208044 237220 208050 237222
rect 214557 237219 214623 237222
rect 223614 237220 223620 237284
rect 223684 237282 223690 237284
rect 582741 237282 582807 237285
rect 223684 237280 582807 237282
rect 223684 237224 582746 237280
rect 582802 237224 582807 237280
rect 223684 237222 582807 237224
rect 223684 237220 223690 237222
rect 582741 237219 582807 237222
rect 127065 237146 127131 237149
rect 160093 237146 160159 237149
rect 240685 237146 240751 237149
rect 127065 237144 240751 237146
rect 127065 237088 127070 237144
rect 127126 237088 160098 237144
rect 160154 237088 240690 237144
rect 240746 237088 240751 237144
rect 127065 237086 240751 237088
rect 127065 237083 127131 237086
rect 160093 237083 160159 237086
rect 240685 237083 240751 237086
rect 137134 236948 137140 237012
rect 137204 237010 137210 237012
rect 178953 237010 179019 237013
rect 137204 237008 179019 237010
rect 137204 236952 178958 237008
rect 179014 236952 179019 237008
rect 137204 236950 179019 236952
rect 137204 236948 137210 236950
rect 178953 236947 179019 236950
rect 52085 236602 52151 236605
rect 128353 236602 128419 236605
rect 52085 236600 128419 236602
rect 52085 236544 52090 236600
rect 52146 236544 128358 236600
rect 128414 236544 128419 236600
rect 52085 236542 128419 236544
rect 52085 236539 52151 236542
rect 128353 236539 128419 236542
rect 177389 236602 177455 236605
rect 186262 236602 186268 236604
rect 177389 236600 186268 236602
rect 177389 236544 177394 236600
rect 177450 236544 186268 236600
rect 177389 236542 186268 236544
rect 177389 236539 177455 236542
rect 186262 236540 186268 236542
rect 186332 236540 186338 236604
rect 67950 235860 67956 235924
rect 68020 235922 68026 235924
rect 245929 235922 245995 235925
rect 68020 235920 245995 235922
rect 68020 235864 245934 235920
rect 245990 235864 245995 235920
rect 68020 235862 245995 235864
rect 68020 235860 68026 235862
rect 245929 235859 245995 235862
rect 120073 235786 120139 235789
rect 157333 235786 157399 235789
rect 173249 235786 173315 235789
rect 244641 235786 244707 235789
rect 120073 235784 173315 235786
rect 120073 235728 120078 235784
rect 120134 235728 157338 235784
rect 157394 235728 173254 235784
rect 173310 235728 173315 235784
rect 120073 235726 173315 235728
rect 120073 235723 120139 235726
rect 157333 235723 157399 235726
rect 173249 235723 173315 235726
rect 180750 235784 244707 235786
rect 180750 235728 244646 235784
rect 244702 235728 244707 235784
rect 180750 235726 244707 235728
rect 151813 235650 151879 235653
rect 179413 235650 179479 235653
rect 180750 235650 180810 235726
rect 244641 235723 244707 235726
rect 151813 235648 180810 235650
rect 151813 235592 151818 235648
rect 151874 235592 179418 235648
rect 179474 235592 180810 235648
rect 151813 235590 180810 235592
rect 151813 235587 151879 235590
rect 179413 235587 179479 235590
rect 186262 235588 186268 235652
rect 186332 235650 186338 235652
rect 210325 235650 210391 235653
rect 186332 235648 210391 235650
rect 186332 235592 210330 235648
rect 210386 235592 210391 235648
rect 186332 235590 210391 235592
rect 186332 235588 186338 235590
rect 210325 235587 210391 235590
rect 242341 235242 242407 235245
rect 249701 235242 249767 235245
rect 291929 235242 291995 235245
rect 242341 235240 291995 235242
rect 242341 235184 242346 235240
rect 242402 235184 249706 235240
rect 249762 235184 291934 235240
rect 291990 235184 291995 235240
rect 242341 235182 291995 235184
rect 242341 235179 242407 235182
rect 249701 235179 249767 235182
rect 291929 235179 291995 235182
rect 135989 234698 136055 234701
rect 153009 234698 153075 234701
rect 135989 234696 153075 234698
rect 135989 234640 135994 234696
rect 136050 234640 153014 234696
rect 153070 234640 153075 234696
rect 135989 234638 153075 234640
rect 135989 234635 136055 234638
rect 153009 234635 153075 234638
rect 64689 234562 64755 234565
rect 216029 234562 216095 234565
rect 244089 234562 244155 234565
rect 64689 234560 244155 234562
rect 64689 234504 64694 234560
rect 64750 234504 216034 234560
rect 216090 234504 244094 234560
rect 244150 234504 244155 234560
rect 64689 234502 244155 234504
rect 64689 234499 64755 234502
rect 216029 234499 216095 234502
rect 244089 234499 244155 234502
rect 71773 234426 71839 234429
rect 160829 234426 160895 234429
rect 71773 234424 160895 234426
rect 71773 234368 71778 234424
rect 71834 234368 160834 234424
rect 160890 234368 160895 234424
rect 71773 234366 160895 234368
rect 71773 234363 71839 234366
rect 160829 234363 160895 234366
rect 187141 234426 187207 234429
rect 208853 234426 208919 234429
rect 187141 234424 208919 234426
rect 187141 234368 187146 234424
rect 187202 234368 208858 234424
rect 208914 234368 208919 234424
rect 187141 234366 208919 234368
rect 187141 234363 187207 234366
rect 208853 234363 208919 234366
rect 146385 234290 146451 234293
rect 162301 234290 162367 234293
rect 146385 234288 162367 234290
rect 146385 234232 146390 234288
rect 146446 234232 162306 234288
rect 162362 234232 162367 234288
rect 146385 234230 162367 234232
rect 146385 234227 146451 234230
rect 162301 234227 162367 234230
rect 139209 234018 139275 234021
rect 139710 234018 139716 234020
rect 139209 234016 139716 234018
rect 139209 233960 139214 234016
rect 139270 233960 139716 234016
rect 139209 233958 139716 233960
rect 139209 233955 139275 233958
rect 139710 233956 139716 233958
rect 139780 233956 139786 234020
rect 216673 234018 216739 234021
rect 230197 234018 230263 234021
rect 216673 234016 230263 234018
rect 216673 233960 216678 234016
rect 216734 233960 230202 234016
rect 230258 233960 230263 234016
rect 216673 233958 230263 233960
rect 216673 233955 216739 233958
rect 230197 233955 230263 233958
rect 170949 233882 171015 233885
rect 203517 233882 203583 233885
rect 170949 233880 203583 233882
rect 170949 233824 170954 233880
rect 171010 233824 203522 233880
rect 203578 233824 203583 233880
rect 170949 233822 203583 233824
rect 170949 233819 171015 233822
rect 203517 233819 203583 233822
rect 209681 233882 209747 233885
rect 215518 233882 215524 233884
rect 209681 233880 215524 233882
rect 209681 233824 209686 233880
rect 209742 233824 215524 233880
rect 209681 233822 215524 233824
rect 209681 233819 209747 233822
rect 215518 233820 215524 233822
rect 215588 233820 215594 233884
rect 222101 233882 222167 233885
rect 316033 233882 316099 233885
rect 222101 233880 316099 233882
rect 222101 233824 222106 233880
rect 222162 233824 316038 233880
rect 316094 233824 316099 233880
rect 222101 233822 316099 233824
rect 222101 233819 222167 233822
rect 316033 233819 316099 233822
rect 67633 233202 67699 233205
rect 231485 233202 231551 233205
rect 67633 233200 231551 233202
rect 67633 233144 67638 233200
rect 67694 233144 231490 233200
rect 231546 233144 231551 233200
rect 67633 233142 231551 233144
rect 67633 233139 67699 233142
rect 231485 233139 231551 233142
rect 140773 233066 140839 233069
rect 234061 233066 234127 233069
rect 140773 233064 234127 233066
rect 140773 233008 140778 233064
rect 140834 233008 234066 233064
rect 234122 233008 234127 233064
rect 140773 233006 234127 233008
rect 140773 233003 140839 233006
rect 234061 233003 234127 233006
rect 113173 232930 113239 232933
rect 143574 232930 143580 232932
rect 113173 232928 143580 232930
rect 113173 232872 113178 232928
rect 113234 232872 143580 232928
rect 113173 232870 143580 232872
rect 113173 232867 113239 232870
rect 143574 232868 143580 232870
rect 143644 232930 143650 232932
rect 209221 232930 209287 232933
rect 143644 232928 209287 232930
rect 143644 232872 209226 232928
rect 209282 232872 209287 232928
rect 143644 232870 209287 232872
rect 143644 232868 143650 232870
rect 209221 232867 209287 232870
rect 211797 232930 211863 232933
rect 212625 232930 212691 232933
rect 211797 232928 212691 232930
rect 211797 232872 211802 232928
rect 211858 232872 212630 232928
rect 212686 232872 212691 232928
rect 211797 232870 212691 232872
rect 211797 232867 211863 232870
rect 212625 232867 212691 232870
rect 251817 232658 251883 232661
rect 266445 232658 266511 232661
rect 251817 232656 266511 232658
rect 251817 232600 251822 232656
rect 251878 232600 266450 232656
rect 266506 232600 266511 232656
rect 251817 232598 266511 232600
rect 251817 232595 251883 232598
rect 266445 232595 266511 232598
rect 223389 232522 223455 232525
rect 280337 232522 280403 232525
rect 223389 232520 280403 232522
rect 223389 232464 223394 232520
rect 223450 232464 280342 232520
rect 280398 232464 280403 232520
rect 223389 232462 280403 232464
rect 223389 232459 223455 232462
rect 280337 232459 280403 232462
rect 582649 232386 582715 232389
rect 583520 232386 584960 232476
rect 582649 232384 584960 232386
rect 582649 232328 582654 232384
rect 582710 232328 584960 232384
rect 582649 232326 584960 232328
rect 582649 232323 582715 232326
rect 583520 232236 584960 232326
rect 103329 231842 103395 231845
rect 166993 231842 167059 231845
rect 232957 231842 233023 231845
rect 103329 231840 233023 231842
rect 103329 231784 103334 231840
rect 103390 231784 166998 231840
rect 167054 231784 232962 231840
rect 233018 231784 233023 231840
rect 103329 231782 233023 231784
rect 103329 231779 103395 231782
rect 166993 231779 167059 231782
rect 232957 231779 233023 231782
rect 143441 231706 143507 231709
rect 163589 231706 163655 231709
rect 143441 231704 163655 231706
rect 143441 231648 143446 231704
rect 143502 231648 163594 231704
rect 163650 231648 163655 231704
rect 143441 231646 163655 231648
rect 143441 231643 143507 231646
rect 163589 231643 163655 231646
rect 182817 231706 182883 231709
rect 224217 231706 224283 231709
rect 224861 231706 224927 231709
rect 182817 231704 224927 231706
rect 182817 231648 182822 231704
rect 182878 231648 224222 231704
rect 224278 231648 224866 231704
rect 224922 231648 224927 231704
rect 182817 231646 224927 231648
rect 182817 231643 182883 231646
rect 224217 231643 224283 231646
rect 224861 231643 224927 231646
rect 145925 231570 145991 231573
rect 158161 231570 158227 231573
rect 197077 231572 197143 231573
rect 197077 231570 197124 231572
rect 145925 231568 158227 231570
rect 145925 231512 145930 231568
rect 145986 231512 158166 231568
rect 158222 231512 158227 231568
rect 145925 231510 158227 231512
rect 197032 231568 197124 231570
rect 197032 231512 197082 231568
rect 197032 231510 197124 231512
rect 145925 231507 145991 231510
rect 158161 231507 158227 231510
rect 197077 231508 197124 231510
rect 197188 231508 197194 231572
rect 197077 231507 197143 231508
rect 154614 231372 154620 231436
rect 154684 231434 154690 231436
rect 155861 231434 155927 231437
rect 154684 231432 155927 231434
rect 154684 231376 155866 231432
rect 155922 231376 155927 231432
rect 154684 231374 155927 231376
rect 154684 231372 154690 231374
rect 155861 231371 155927 231374
rect 56317 231162 56383 231165
rect 146201 231162 146267 231165
rect 56317 231160 146267 231162
rect 56317 231104 56322 231160
rect 56378 231104 146206 231160
rect 146262 231104 146267 231160
rect 56317 231102 146267 231104
rect 56317 231099 56383 231102
rect 146201 231099 146267 231102
rect 197077 230618 197143 230621
rect 325785 230618 325851 230621
rect 197077 230616 325851 230618
rect 197077 230560 197082 230616
rect 197138 230560 325790 230616
rect 325846 230560 325851 230616
rect 197077 230558 325851 230560
rect 197077 230555 197143 230558
rect 325785 230555 325851 230558
rect 59077 230482 59143 230485
rect 245878 230482 245884 230484
rect 59077 230480 245884 230482
rect 59077 230424 59082 230480
rect 59138 230424 245884 230480
rect 59077 230422 245884 230424
rect 59077 230419 59143 230422
rect 245878 230420 245884 230422
rect 245948 230420 245954 230484
rect 108297 230346 108363 230349
rect 154062 230346 154068 230348
rect 108297 230344 154068 230346
rect 108297 230288 108302 230344
rect 108358 230288 154068 230344
rect 108297 230286 154068 230288
rect 108297 230283 108363 230286
rect 154062 230284 154068 230286
rect 154132 230284 154138 230348
rect 172421 230346 172487 230349
rect 195329 230346 195395 230349
rect 172421 230344 195395 230346
rect 172421 230288 172426 230344
rect 172482 230288 195334 230344
rect 195390 230288 195395 230344
rect 172421 230286 195395 230288
rect 172421 230283 172487 230286
rect 195329 230283 195395 230286
rect 135161 230210 135227 230213
rect 167637 230210 167703 230213
rect 135161 230208 167703 230210
rect 135161 230152 135166 230208
rect 135222 230152 167642 230208
rect 167698 230152 167703 230208
rect 135161 230150 167703 230152
rect 135161 230147 135227 230150
rect 167637 230147 167703 230150
rect 195881 229938 195947 229941
rect 232589 229938 232655 229941
rect 195881 229936 232655 229938
rect 195881 229880 195886 229936
rect 195942 229880 232594 229936
rect 232650 229880 232655 229936
rect 195881 229878 232655 229880
rect 195881 229875 195947 229878
rect 232589 229875 232655 229878
rect 233877 229938 233943 229941
rect 278814 229938 278820 229940
rect 233877 229936 278820 229938
rect 233877 229880 233882 229936
rect 233938 229880 278820 229936
rect 233877 229878 278820 229880
rect 233877 229875 233943 229878
rect 278814 229876 278820 229878
rect 278884 229876 278890 229940
rect 195830 229740 195836 229804
rect 195900 229802 195906 229804
rect 583293 229802 583359 229805
rect 195900 229800 583359 229802
rect 195900 229744 583298 229800
rect 583354 229744 583359 229800
rect 195900 229742 583359 229744
rect 195900 229740 195906 229742
rect 583293 229739 583359 229742
rect 315941 229122 316007 229125
rect 316166 229122 316172 229124
rect 315896 229120 316172 229122
rect 315896 229064 315946 229120
rect 316002 229064 316172 229120
rect 315896 229062 316172 229064
rect 315941 229059 316007 229062
rect 316166 229060 316172 229062
rect 316236 229060 316242 229124
rect 123477 228986 123543 228989
rect 155166 228986 155172 228988
rect 123477 228984 155172 228986
rect 123477 228928 123482 228984
rect 123538 228928 155172 228984
rect 123477 228926 155172 228928
rect 123477 228923 123543 228926
rect 155166 228924 155172 228926
rect 155236 228924 155242 228988
rect 200113 228986 200179 228989
rect 245653 228986 245719 228989
rect 315941 228986 316007 228989
rect 316166 228986 316172 228988
rect 200113 228984 245719 228986
rect 200113 228928 200118 228984
rect 200174 228928 245658 228984
rect 245714 228928 245719 228984
rect 200113 228926 245719 228928
rect 315896 228984 316172 228986
rect 315896 228928 315946 228984
rect 316002 228928 316172 228984
rect 315896 228926 316172 228928
rect 200113 228923 200179 228926
rect 245653 228923 245719 228926
rect 315941 228923 316007 228926
rect 316166 228924 316172 228926
rect 316236 228924 316242 228988
rect 146201 228850 146267 228853
rect 162393 228850 162459 228853
rect 146201 228848 162459 228850
rect 146201 228792 146206 228848
rect 146262 228792 162398 228848
rect 162454 228792 162459 228848
rect 146201 228790 162459 228792
rect 146201 228787 146267 228790
rect 162393 228787 162459 228790
rect 172421 228442 172487 228445
rect 197077 228442 197143 228445
rect 172421 228440 197143 228442
rect 172421 228384 172426 228440
rect 172482 228384 197082 228440
rect 197138 228384 197143 228440
rect 172421 228382 197143 228384
rect 172421 228379 172487 228382
rect 197077 228379 197143 228382
rect 90909 228306 90975 228309
rect 151077 228306 151143 228309
rect 90909 228304 151143 228306
rect 90909 228248 90914 228304
rect 90970 228248 151082 228304
rect 151138 228248 151143 228304
rect 90909 228246 151143 228248
rect 90909 228243 90975 228246
rect 151077 228243 151143 228246
rect 188981 228306 189047 228309
rect 332685 228306 332751 228309
rect 188981 228304 332751 228306
rect 188981 228248 188986 228304
rect 189042 228248 332690 228304
rect 332746 228248 332751 228304
rect 188981 228246 332751 228248
rect 188981 228243 189047 228246
rect 332685 228243 332751 228246
rect -960 227884 480 228124
rect 173709 227762 173775 227765
rect 200205 227762 200271 227765
rect 200849 227762 200915 227765
rect 173709 227760 200915 227762
rect 173709 227704 173714 227760
rect 173770 227704 200210 227760
rect 200266 227704 200854 227760
rect 200910 227704 200915 227760
rect 173709 227702 200915 227704
rect 173709 227699 173775 227702
rect 200205 227699 200271 227702
rect 200849 227699 200915 227702
rect 245653 227762 245719 227765
rect 246297 227762 246363 227765
rect 245653 227760 246363 227762
rect 245653 227704 245658 227760
rect 245714 227704 246302 227760
rect 246358 227704 246363 227760
rect 245653 227702 246363 227704
rect 245653 227699 245719 227702
rect 246297 227699 246363 227702
rect 50797 227626 50863 227629
rect 218697 227626 218763 227629
rect 50797 227624 218763 227626
rect 50797 227568 50802 227624
rect 50858 227568 218702 227624
rect 218758 227568 218763 227624
rect 50797 227566 218763 227568
rect 50797 227563 50863 227566
rect 218697 227563 218763 227566
rect 84694 227428 84700 227492
rect 84764 227490 84770 227492
rect 245694 227490 245700 227492
rect 84764 227430 245700 227490
rect 84764 227428 84770 227430
rect 245694 227428 245700 227430
rect 245764 227428 245770 227492
rect 129549 227354 129615 227357
rect 163497 227354 163563 227357
rect 244365 227354 244431 227357
rect 129549 227352 244431 227354
rect 129549 227296 129554 227352
rect 129610 227296 163502 227352
rect 163558 227296 244370 227352
rect 244426 227296 244431 227352
rect 129549 227294 244431 227296
rect 129549 227291 129615 227294
rect 163497 227291 163563 227294
rect 244365 227291 244431 227294
rect 84101 226266 84167 226269
rect 239765 226266 239831 226269
rect 84101 226264 239831 226266
rect 84101 226208 84106 226264
rect 84162 226208 239770 226264
rect 239826 226208 239831 226264
rect 84101 226206 239831 226208
rect 84101 226203 84167 226206
rect 239765 226203 239831 226206
rect 67725 226130 67791 226133
rect 159633 226130 159699 226133
rect 67725 226128 159699 226130
rect 67725 226072 67730 226128
rect 67786 226072 159638 226128
rect 159694 226072 159699 226128
rect 67725 226070 159699 226072
rect 67725 226067 67791 226070
rect 159633 226067 159699 226070
rect 167637 226130 167703 226133
rect 204989 226130 205055 226133
rect 167637 226128 205055 226130
rect 167637 226072 167642 226128
rect 167698 226072 204994 226128
rect 205050 226072 205055 226128
rect 167637 226070 205055 226072
rect 167637 226067 167703 226070
rect 204989 226067 205055 226070
rect 79317 225994 79383 225997
rect 166533 225994 166599 225997
rect 79317 225992 166599 225994
rect 79317 225936 79322 225992
rect 79378 225936 166538 225992
rect 166594 225936 166599 225992
rect 79317 225934 166599 225936
rect 79317 225931 79383 225934
rect 166533 225931 166599 225934
rect 195053 225586 195119 225589
rect 242341 225586 242407 225589
rect 195053 225584 242407 225586
rect 195053 225528 195058 225584
rect 195114 225528 242346 225584
rect 242402 225528 242407 225584
rect 195053 225526 242407 225528
rect 195053 225523 195119 225526
rect 242341 225523 242407 225526
rect 53557 224906 53623 224909
rect 234981 224906 235047 224909
rect 53557 224904 235047 224906
rect 53557 224848 53562 224904
rect 53618 224848 234986 224904
rect 235042 224848 235047 224904
rect 53557 224846 235047 224848
rect 53557 224843 53623 224846
rect 234981 224843 235047 224846
rect 107469 224770 107535 224773
rect 140814 224770 140820 224772
rect 107469 224768 140820 224770
rect 107469 224712 107474 224768
rect 107530 224712 140820 224768
rect 107469 224710 140820 224712
rect 107469 224707 107535 224710
rect 140814 224708 140820 224710
rect 140884 224770 140890 224772
rect 251357 224770 251423 224773
rect 140884 224768 251423 224770
rect 140884 224712 251362 224768
rect 251418 224712 251423 224768
rect 140884 224710 251423 224712
rect 140884 224708 140890 224710
rect 251357 224707 251423 224710
rect 185669 224226 185735 224229
rect 205081 224226 205147 224229
rect 185669 224224 205147 224226
rect 185669 224168 185674 224224
rect 185730 224168 205086 224224
rect 205142 224168 205147 224224
rect 185669 224166 205147 224168
rect 185669 224163 185735 224166
rect 205081 224163 205147 224166
rect 63309 223546 63375 223549
rect 173709 223546 173775 223549
rect 63309 223544 173775 223546
rect 63309 223488 63314 223544
rect 63370 223488 173714 223544
rect 173770 223488 173775 223544
rect 63309 223486 173775 223488
rect 63309 223483 63375 223486
rect 173709 223483 173775 223486
rect 276013 223546 276079 223549
rect 276238 223546 276244 223548
rect 276013 223544 276244 223546
rect 276013 223488 276018 223544
rect 276074 223488 276244 223544
rect 276013 223486 276244 223488
rect 276013 223483 276079 223486
rect 276238 223484 276244 223486
rect 276308 223484 276314 223548
rect 137277 223410 137343 223413
rect 196709 223410 196775 223413
rect 137277 223408 196775 223410
rect 137277 223352 137282 223408
rect 137338 223352 196714 223408
rect 196770 223352 196775 223408
rect 137277 223350 196775 223352
rect 137277 223347 137343 223350
rect 196709 223347 196775 223350
rect 199510 222940 199516 223004
rect 199580 223002 199586 223004
rect 258717 223002 258783 223005
rect 199580 223000 258783 223002
rect 199580 222944 258722 223000
rect 258778 222944 258783 223000
rect 199580 222942 258783 222944
rect 199580 222940 199586 222942
rect 258717 222939 258783 222942
rect 156689 222866 156755 222869
rect 353293 222866 353359 222869
rect 156689 222864 353359 222866
rect 156689 222808 156694 222864
rect 156750 222808 353298 222864
rect 353354 222808 353359 222864
rect 156689 222806 353359 222808
rect 156689 222803 156755 222806
rect 353293 222803 353359 222806
rect 4797 222322 4863 222325
rect 155861 222322 155927 222325
rect 4797 222320 155927 222322
rect 4797 222264 4802 222320
rect 4858 222264 155866 222320
rect 155922 222264 155927 222320
rect 4797 222262 155927 222264
rect 4797 222259 4863 222262
rect 155861 222259 155927 222262
rect 217317 222322 217383 222325
rect 217542 222322 217548 222324
rect 217317 222320 217548 222322
rect 217317 222264 217322 222320
rect 217378 222264 217548 222320
rect 217317 222262 217548 222264
rect 217317 222259 217383 222262
rect 217542 222260 217548 222262
rect 217612 222322 217618 222324
rect 283005 222322 283071 222325
rect 217612 222320 283071 222322
rect 217612 222264 283010 222320
rect 283066 222264 283071 222320
rect 217612 222262 283071 222264
rect 217612 222260 217618 222262
rect 283005 222259 283071 222262
rect 69790 222124 69796 222188
rect 69860 222186 69866 222188
rect 205633 222186 205699 222189
rect 69860 222184 205699 222186
rect 69860 222128 205638 222184
rect 205694 222128 205699 222184
rect 69860 222126 205699 222128
rect 69860 222124 69866 222126
rect 205633 222123 205699 222126
rect 118877 222050 118943 222053
rect 193857 222050 193923 222053
rect 118877 222048 193923 222050
rect 118877 221992 118882 222048
rect 118938 221992 193862 222048
rect 193918 221992 193923 222048
rect 118877 221990 193923 221992
rect 118877 221987 118943 221990
rect 193857 221987 193923 221990
rect 194685 221778 194751 221781
rect 209865 221778 209931 221781
rect 194685 221776 209931 221778
rect 194685 221720 194690 221776
rect 194746 221720 209870 221776
rect 209926 221720 209931 221776
rect 194685 221718 209931 221720
rect 194685 221715 194751 221718
rect 209865 221715 209931 221718
rect 205633 221642 205699 221645
rect 206461 221642 206527 221645
rect 238017 221642 238083 221645
rect 205633 221640 238083 221642
rect 205633 221584 205638 221640
rect 205694 221584 206466 221640
rect 206522 221584 238022 221640
rect 238078 221584 238083 221640
rect 205633 221582 238083 221584
rect 205633 221579 205699 221582
rect 206461 221579 206527 221582
rect 238017 221579 238083 221582
rect 67265 221506 67331 221509
rect 356053 221506 356119 221509
rect 67265 221504 356119 221506
rect 67265 221448 67270 221504
rect 67326 221448 356058 221504
rect 356114 221448 356119 221504
rect 67265 221446 356119 221448
rect 67265 221443 67331 221446
rect 356053 221443 356119 221446
rect 88977 220826 89043 220829
rect 206369 220826 206435 220829
rect 253933 220826 253999 220829
rect 254577 220826 254643 220829
rect 88977 220824 206435 220826
rect 88977 220768 88982 220824
rect 89038 220768 206374 220824
rect 206430 220768 206435 220824
rect 88977 220766 206435 220768
rect 88977 220763 89043 220766
rect 206369 220763 206435 220766
rect 238710 220824 254643 220826
rect 238710 220768 253938 220824
rect 253994 220768 254582 220824
rect 254638 220768 254643 220824
rect 238710 220766 254643 220768
rect 73797 220690 73863 220693
rect 188521 220690 188587 220693
rect 73797 220688 188587 220690
rect 73797 220632 73802 220688
rect 73858 220632 188526 220688
rect 188582 220632 188587 220688
rect 73797 220630 188587 220632
rect 73797 220627 73863 220630
rect 188521 220627 188587 220630
rect 142153 220554 142219 220557
rect 238710 220554 238770 220766
rect 253933 220763 253999 220766
rect 254577 220763 254643 220766
rect 142153 220552 238770 220554
rect 142153 220496 142158 220552
rect 142214 220496 238770 220552
rect 142153 220494 238770 220496
rect 142153 220491 142219 220494
rect 266997 220282 267063 220285
rect 273478 220282 273484 220284
rect 266997 220280 273484 220282
rect 266997 220224 267002 220280
rect 267058 220224 273484 220280
rect 266997 220222 273484 220224
rect 266997 220219 267063 220222
rect 273478 220220 273484 220222
rect 273548 220220 273554 220284
rect 260097 220146 260163 220149
rect 318977 220146 319043 220149
rect 260097 220144 319043 220146
rect 260097 220088 260102 220144
rect 260158 220088 318982 220144
rect 319038 220088 319043 220144
rect 260097 220086 319043 220088
rect 260097 220083 260163 220086
rect 318977 220083 319043 220086
rect 315941 219468 316007 219469
rect 315941 219466 315988 219468
rect 315896 219464 315988 219466
rect 316052 219466 316058 219468
rect 315896 219408 315946 219464
rect 315896 219406 315988 219408
rect 315941 219404 315988 219406
rect 316052 219406 316134 219466
rect 316052 219404 316058 219406
rect 315941 219403 316007 219404
rect 64597 219330 64663 219333
rect 182909 219330 182975 219333
rect 64597 219328 182975 219330
rect 64597 219272 64602 219328
rect 64658 219272 182914 219328
rect 182970 219272 182975 219328
rect 64597 219270 182975 219272
rect 64597 219267 64663 219270
rect 182909 219267 182975 219270
rect 191833 219330 191899 219333
rect 195789 219330 195855 219333
rect 191833 219328 195855 219330
rect 191833 219272 191838 219328
rect 191894 219272 195794 219328
rect 195850 219272 195855 219328
rect 191833 219270 195855 219272
rect 191833 219267 191899 219270
rect 195789 219267 195855 219270
rect 203517 219330 203583 219333
rect 244457 219330 244523 219333
rect 315941 219330 316007 219333
rect 583477 219330 583543 219333
rect 203517 219328 244523 219330
rect 203517 219272 203522 219328
rect 203578 219272 244462 219328
rect 244518 219272 244523 219328
rect 203517 219270 244523 219272
rect 315896 219328 316050 219330
rect 315896 219272 315946 219328
rect 316002 219272 316050 219328
rect 315896 219270 316050 219272
rect 203517 219267 203583 219270
rect 244457 219267 244523 219270
rect 315941 219267 316050 219270
rect 583477 219328 583586 219330
rect 583477 219272 583482 219328
rect 583538 219272 583586 219328
rect 583477 219267 583586 219272
rect 55029 219194 55095 219197
rect 159725 219194 159791 219197
rect 315990 219196 316050 219267
rect 55029 219192 159791 219194
rect 55029 219136 55034 219192
rect 55090 219136 159730 219192
rect 159786 219136 159791 219192
rect 55029 219134 159791 219136
rect 55029 219131 55095 219134
rect 159725 219131 159791 219134
rect 315982 219132 315988 219196
rect 316052 219132 316058 219196
rect 583526 219194 583586 219267
rect 583342 219148 583586 219194
rect 583342 219134 584960 219148
rect 583342 219058 583402 219134
rect 583520 219058 584960 219134
rect 583342 218998 584960 219058
rect 583520 218908 584960 218998
rect 77150 218588 77156 218652
rect 77220 218650 77226 218652
rect 324313 218650 324379 218653
rect 77220 218648 324379 218650
rect 77220 218592 324318 218648
rect 324374 218592 324379 218648
rect 77220 218590 324379 218592
rect 77220 218588 77226 218590
rect 324313 218587 324379 218590
rect 224861 218106 224927 218109
rect 225781 218106 225847 218109
rect 224861 218104 225847 218106
rect 224861 218048 224866 218104
rect 224922 218048 225786 218104
rect 225842 218048 225847 218104
rect 224861 218046 225847 218048
rect 224861 218043 224927 218046
rect 225781 218043 225847 218046
rect 56409 217970 56475 217973
rect 217225 217970 217291 217973
rect 56409 217968 217291 217970
rect 56409 217912 56414 217968
rect 56470 217912 217230 217968
rect 217286 217912 217291 217968
rect 56409 217910 217291 217912
rect 56409 217907 56475 217910
rect 217225 217907 217291 217910
rect 155861 217834 155927 217837
rect 221457 217834 221523 217837
rect 155861 217832 221523 217834
rect 155861 217776 155866 217832
rect 155922 217776 221462 217832
rect 221518 217776 221523 217832
rect 155861 217774 221523 217776
rect 155861 217771 155927 217774
rect 221457 217771 221523 217774
rect 92289 217290 92355 217293
rect 181529 217290 181595 217293
rect 92289 217288 181595 217290
rect 92289 217232 92294 217288
rect 92350 217232 181534 217288
rect 181590 217232 181595 217288
rect 92289 217230 181595 217232
rect 92289 217227 92355 217230
rect 181529 217227 181595 217230
rect 217225 217290 217291 217293
rect 260097 217290 260163 217293
rect 217225 217288 260163 217290
rect 217225 217232 217230 217288
rect 217286 217232 260102 217288
rect 260158 217232 260163 217288
rect 217225 217230 260163 217232
rect 217225 217227 217291 217230
rect 260097 217227 260163 217230
rect 192477 216746 192543 216749
rect 197997 216746 198063 216749
rect 192477 216744 198063 216746
rect 192477 216688 192482 216744
rect 192538 216688 198002 216744
rect 198058 216688 198063 216744
rect 192477 216686 198063 216688
rect 192477 216683 192543 216686
rect 197997 216683 198063 216686
rect 207381 216746 207447 216749
rect 207749 216746 207815 216749
rect 302182 216746 302188 216748
rect 207381 216744 302188 216746
rect 207381 216688 207386 216744
rect 207442 216688 207754 216744
rect 207810 216688 302188 216744
rect 207381 216686 302188 216688
rect 207381 216683 207447 216686
rect 207749 216683 207815 216686
rect 302182 216684 302188 216686
rect 302252 216684 302258 216748
rect 60549 216610 60615 216613
rect 205357 216610 205423 216613
rect 60549 216608 205423 216610
rect 60549 216552 60554 216608
rect 60610 216552 205362 216608
rect 205418 216552 205423 216608
rect 60549 216550 205423 216552
rect 60549 216547 60615 216550
rect 205357 216547 205423 216550
rect 69657 216474 69723 216477
rect 178534 216474 178540 216476
rect 69657 216472 178540 216474
rect 69657 216416 69662 216472
rect 69718 216416 178540 216472
rect 69657 216414 178540 216416
rect 69657 216411 69723 216414
rect 178534 216412 178540 216414
rect 178604 216412 178610 216476
rect 153101 216338 153167 216341
rect 238293 216338 238359 216341
rect 153101 216336 238770 216338
rect 153101 216280 153106 216336
rect 153162 216280 238298 216336
rect 238354 216280 238770 216336
rect 153101 216278 238770 216280
rect 153101 216275 153167 216278
rect 238293 216275 238359 216278
rect 200757 215930 200823 215933
rect 226977 215930 227043 215933
rect 200757 215928 227043 215930
rect 200757 215872 200762 215928
rect 200818 215872 226982 215928
rect 227038 215872 227043 215928
rect 200757 215870 227043 215872
rect 238710 215930 238770 216278
rect 276606 215930 276612 215932
rect 238710 215870 276612 215930
rect 200757 215867 200823 215870
rect 226977 215867 227043 215870
rect 276606 215868 276612 215870
rect 276676 215868 276682 215932
rect 178033 215386 178099 215389
rect 195329 215386 195395 215389
rect 178033 215384 195395 215386
rect 178033 215328 178038 215384
rect 178094 215328 195334 215384
rect 195390 215328 195395 215384
rect 178033 215326 195395 215328
rect 178033 215323 178099 215326
rect 195329 215323 195395 215326
rect 204897 215386 204963 215389
rect 205357 215386 205423 215389
rect 204897 215384 205423 215386
rect 204897 215328 204902 215384
rect 204958 215328 205362 215384
rect 205418 215328 205423 215384
rect 204897 215326 205423 215328
rect 204897 215323 204963 215326
rect 205357 215323 205423 215326
rect 235993 215386 236059 215389
rect 236729 215386 236795 215389
rect 336733 215386 336799 215389
rect 235993 215384 336799 215386
rect 235993 215328 235998 215384
rect 236054 215328 236734 215384
rect 236790 215328 336738 215384
rect 336794 215328 336799 215384
rect 235993 215326 336799 215328
rect 235993 215323 236059 215326
rect 236729 215323 236795 215326
rect 336733 215323 336799 215326
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 77385 214842 77451 214845
rect 152457 214842 152523 214845
rect 77385 214840 152523 214842
rect 77385 214784 77390 214840
rect 77446 214784 152462 214840
rect 152518 214784 152523 214840
rect 77385 214782 152523 214784
rect 77385 214779 77451 214782
rect 152457 214779 152523 214782
rect 154389 214842 154455 214845
rect 178677 214842 178743 214845
rect 154389 214840 178743 214842
rect 154389 214784 154394 214840
rect 154450 214784 178682 214840
rect 178738 214784 178743 214840
rect 154389 214782 178743 214784
rect 154389 214779 154455 214782
rect 178677 214779 178743 214782
rect 107561 214706 107627 214709
rect 187049 214706 187115 214709
rect 107561 214704 187115 214706
rect 107561 214648 107566 214704
rect 107622 214648 187054 214704
rect 187110 214648 187115 214704
rect 107561 214646 187115 214648
rect 107561 214643 107627 214646
rect 187049 214643 187115 214646
rect 187233 214706 187299 214709
rect 296069 214706 296135 214709
rect 187233 214704 296135 214706
rect 187233 214648 187238 214704
rect 187294 214648 296074 214704
rect 296130 214648 296135 214704
rect 187233 214646 296135 214648
rect 187233 214643 187299 214646
rect 296069 214643 296135 214646
rect 65926 214508 65932 214572
rect 65996 214570 66002 214572
rect 342253 214570 342319 214573
rect 65996 214568 342319 214570
rect 65996 214512 342258 214568
rect 342314 214512 342319 214568
rect 65996 214510 342319 214512
rect 65996 214508 66002 214510
rect 342253 214507 342319 214510
rect 184289 214026 184355 214029
rect 218973 214026 219039 214029
rect 184289 214024 219039 214026
rect 184289 213968 184294 214024
rect 184350 213968 218978 214024
rect 219034 213968 219039 214024
rect 184289 213966 219039 213968
rect 184289 213963 184355 213966
rect 218973 213963 219039 213966
rect 75177 213890 75243 213893
rect 194685 213890 194751 213893
rect 75177 213888 194751 213890
rect 75177 213832 75182 213888
rect 75238 213832 194690 213888
rect 194746 213832 194751 213888
rect 75177 213830 194751 213832
rect 75177 213827 75243 213830
rect 194685 213827 194751 213830
rect 269113 213890 269179 213893
rect 269246 213890 269252 213892
rect 269113 213888 269252 213890
rect 269113 213832 269118 213888
rect 269174 213832 269252 213888
rect 269113 213830 269252 213832
rect 269113 213827 269179 213830
rect 269246 213828 269252 213830
rect 269316 213828 269322 213892
rect 99281 213346 99347 213349
rect 170397 213346 170463 213349
rect 99281 213344 170463 213346
rect 99281 213288 99286 213344
rect 99342 213288 170402 213344
rect 170458 213288 170463 213344
rect 99281 213286 170463 213288
rect 99281 213283 99347 213286
rect 170397 213283 170463 213286
rect 202229 213346 202295 213349
rect 304349 213346 304415 213349
rect 202229 213344 304415 213346
rect 202229 213288 202234 213344
rect 202290 213288 304354 213344
rect 304410 213288 304415 213344
rect 202229 213286 304415 213288
rect 202229 213283 202295 213286
rect 304349 213283 304415 213286
rect 104893 213210 104959 213213
rect 193029 213210 193095 213213
rect 194041 213210 194107 213213
rect 104893 213208 194107 213210
rect 104893 213152 104898 213208
rect 104954 213152 193034 213208
rect 193090 213152 194046 213208
rect 194102 213152 194107 213208
rect 104893 213150 194107 213152
rect 104893 213147 104959 213150
rect 193029 213147 193095 213150
rect 194041 213147 194107 213150
rect 205081 213210 205147 213213
rect 317597 213210 317663 213213
rect 205081 213208 317663 213210
rect 205081 213152 205086 213208
rect 205142 213152 317602 213208
rect 317658 213152 317663 213208
rect 205081 213150 317663 213152
rect 205081 213147 205147 213150
rect 317597 213147 317663 213150
rect 95233 212530 95299 212533
rect 255313 212530 255379 212533
rect 256049 212530 256115 212533
rect 95233 212528 256115 212530
rect 95233 212472 95238 212528
rect 95294 212472 255318 212528
rect 255374 212472 256054 212528
rect 256110 212472 256115 212528
rect 95233 212470 256115 212472
rect 95233 212467 95299 212470
rect 255313 212467 255379 212470
rect 256049 212467 256115 212470
rect 77109 212394 77175 212397
rect 203149 212394 203215 212397
rect 77109 212392 203215 212394
rect 77109 212336 77114 212392
rect 77170 212336 203154 212392
rect 203210 212336 203215 212392
rect 77109 212334 203215 212336
rect 77109 212331 77175 212334
rect 203149 212331 203215 212334
rect 166257 211850 166323 211853
rect 335445 211850 335511 211853
rect 166257 211848 335511 211850
rect 166257 211792 166262 211848
rect 166318 211792 335450 211848
rect 335506 211792 335511 211848
rect 166257 211790 335511 211792
rect 166257 211787 166323 211790
rect 335445 211787 335511 211790
rect 104801 211034 104867 211037
rect 217501 211034 217567 211037
rect 104801 211032 217567 211034
rect 104801 210976 104806 211032
rect 104862 210976 217506 211032
rect 217562 210976 217567 211032
rect 104801 210974 217567 210976
rect 104801 210971 104867 210974
rect 217501 210971 217567 210974
rect 126881 210898 126947 210901
rect 227253 210898 227319 210901
rect 126881 210896 227319 210898
rect 126881 210840 126886 210896
rect 126942 210840 227258 210896
rect 227314 210840 227319 210896
rect 126881 210838 227319 210840
rect 126881 210835 126947 210838
rect 227253 210835 227319 210838
rect 248321 210626 248387 210629
rect 277526 210626 277532 210628
rect 248321 210624 277532 210626
rect 248321 210568 248326 210624
rect 248382 210568 277532 210624
rect 248321 210566 277532 210568
rect 248321 210563 248387 210566
rect 277526 210564 277532 210566
rect 277596 210564 277602 210628
rect 223021 210490 223087 210493
rect 284518 210490 284524 210492
rect 223021 210488 284524 210490
rect 223021 210432 223026 210488
rect 223082 210432 284524 210488
rect 223021 210430 284524 210432
rect 223021 210427 223087 210430
rect 284518 210428 284524 210430
rect 284588 210428 284594 210492
rect 200849 210354 200915 210357
rect 310462 210354 310468 210356
rect 200849 210352 310468 210354
rect 200849 210296 200854 210352
rect 200910 210296 310468 210352
rect 200849 210294 310468 210296
rect 200849 210291 200915 210294
rect 310462 210292 310468 210294
rect 310532 210292 310538 210356
rect 315941 209812 316007 209813
rect 315941 209810 315988 209812
rect 315896 209808 315988 209810
rect 316052 209810 316058 209812
rect 315896 209752 315946 209808
rect 315896 209750 315988 209752
rect 315941 209748 315988 209750
rect 316052 209750 316134 209810
rect 316052 209748 316058 209750
rect 315941 209747 316007 209748
rect 126789 209674 126855 209677
rect 243997 209674 244063 209677
rect 315941 209674 316007 209677
rect 126789 209672 244063 209674
rect 126789 209616 126794 209672
rect 126850 209616 244002 209672
rect 244058 209616 244063 209672
rect 126789 209614 244063 209616
rect 315896 209672 316050 209674
rect 315896 209616 315946 209672
rect 316002 209616 316050 209672
rect 315896 209614 316050 209616
rect 126789 209611 126855 209614
rect 243997 209611 244063 209614
rect 315941 209611 316050 209614
rect 171961 209538 172027 209541
rect 210417 209538 210483 209541
rect 315990 209540 316050 209611
rect 171961 209536 210483 209538
rect 171961 209480 171966 209536
rect 172022 209480 210422 209536
rect 210478 209480 210483 209536
rect 171961 209478 210483 209480
rect 171961 209475 172027 209478
rect 210417 209475 210483 209478
rect 315982 209476 315988 209540
rect 316052 209476 316058 209540
rect 66662 208932 66668 208996
rect 66732 208994 66738 208996
rect 583477 208994 583543 208997
rect 66732 208992 583543 208994
rect 66732 208936 583482 208992
rect 583538 208936 583543 208992
rect 66732 208934 583543 208936
rect 66732 208932 66738 208934
rect 583477 208931 583543 208934
rect 101949 207770 102015 207773
rect 177389 207770 177455 207773
rect 101949 207768 177455 207770
rect 101949 207712 101954 207768
rect 102010 207712 177394 207768
rect 177450 207712 177455 207768
rect 101949 207710 177455 207712
rect 101949 207707 102015 207710
rect 177389 207707 177455 207710
rect 181437 207770 181503 207773
rect 247677 207770 247743 207773
rect 181437 207768 247743 207770
rect 181437 207712 181442 207768
rect 181498 207712 247682 207768
rect 247738 207712 247743 207768
rect 181437 207710 247743 207712
rect 181437 207707 181503 207710
rect 247677 207707 247743 207710
rect 140681 207634 140747 207637
rect 332593 207634 332659 207637
rect 140681 207632 332659 207634
rect 140681 207576 140686 207632
rect 140742 207576 332598 207632
rect 332654 207576 332659 207632
rect 140681 207574 332659 207576
rect 140681 207571 140747 207574
rect 332593 207571 332659 207574
rect 214414 207028 214420 207092
rect 214484 207090 214490 207092
rect 214649 207090 214715 207093
rect 214484 207088 214715 207090
rect 214484 207032 214654 207088
rect 214710 207032 214715 207088
rect 214484 207030 214715 207032
rect 214484 207028 214490 207030
rect 214649 207027 214715 207030
rect 128261 206954 128327 206957
rect 229737 206954 229803 206957
rect 128261 206952 229803 206954
rect 128261 206896 128266 206952
rect 128322 206896 229742 206952
rect 229798 206896 229803 206952
rect 128261 206894 229803 206896
rect 128261 206891 128327 206894
rect 229737 206891 229803 206894
rect 152457 206818 152523 206821
rect 208393 206818 208459 206821
rect 152457 206816 208459 206818
rect 152457 206760 152462 206816
rect 152518 206760 208398 206816
rect 208454 206760 208459 206816
rect 152457 206758 208459 206760
rect 152457 206755 152523 206758
rect 208393 206755 208459 206758
rect 3509 206274 3575 206277
rect 154614 206274 154620 206276
rect 3509 206272 154620 206274
rect 3509 206216 3514 206272
rect 3570 206216 154620 206272
rect 3509 206214 154620 206216
rect 3509 206211 3575 206214
rect 154614 206212 154620 206214
rect 154684 206212 154690 206276
rect 161974 206212 161980 206276
rect 162044 206274 162050 206276
rect 345013 206274 345079 206277
rect 583753 206274 583819 206277
rect 162044 206272 345079 206274
rect 162044 206216 345018 206272
rect 345074 206216 345079 206272
rect 162044 206214 345079 206216
rect 162044 206212 162050 206214
rect 345013 206211 345079 206214
rect 583710 206272 583819 206274
rect 583710 206216 583758 206272
rect 583814 206216 583819 206272
rect 583710 206211 583819 206216
rect 583710 205866 583770 206211
rect 583342 205820 583770 205866
rect 583342 205806 584960 205820
rect 583342 205730 583402 205806
rect 583520 205730 584960 205806
rect 583342 205670 584960 205730
rect 74533 205594 74599 205597
rect 202965 205594 203031 205597
rect 203609 205594 203675 205597
rect 74533 205592 203675 205594
rect 74533 205536 74538 205592
rect 74594 205536 202970 205592
rect 203026 205536 203614 205592
rect 203670 205536 203675 205592
rect 583520 205580 584960 205670
rect 74533 205534 203675 205536
rect 74533 205531 74599 205534
rect 202965 205531 203031 205534
rect 203609 205531 203675 205534
rect 125501 205458 125567 205461
rect 226149 205458 226215 205461
rect 125501 205456 226215 205458
rect 125501 205400 125506 205456
rect 125562 205400 226154 205456
rect 226210 205400 226215 205456
rect 125501 205398 226215 205400
rect 125501 205395 125567 205398
rect 226149 205395 226215 205398
rect 232589 205050 232655 205053
rect 323025 205050 323091 205053
rect 232589 205048 323091 205050
rect 232589 204992 232594 205048
rect 232650 204992 323030 205048
rect 323086 204992 323091 205048
rect 232589 204990 323091 204992
rect 232589 204987 232655 204990
rect 323025 204987 323091 204990
rect 86861 204914 86927 204917
rect 250437 204914 250503 204917
rect 86861 204912 250503 204914
rect 86861 204856 86866 204912
rect 86922 204856 250442 204912
rect 250498 204856 250503 204912
rect 86861 204854 250503 204856
rect 86861 204851 86927 204854
rect 250437 204851 250503 204854
rect 69606 204172 69612 204236
rect 69676 204234 69682 204236
rect 212574 204234 212580 204236
rect 69676 204174 212580 204234
rect 69676 204172 69682 204174
rect 212574 204172 212580 204174
rect 212644 204234 212650 204236
rect 213126 204234 213132 204236
rect 212644 204174 213132 204234
rect 212644 204172 212650 204174
rect 213126 204172 213132 204174
rect 213196 204172 213202 204236
rect 114461 204098 114527 204101
rect 215937 204098 216003 204101
rect 114461 204096 216003 204098
rect 114461 204040 114466 204096
rect 114522 204040 215942 204096
rect 215998 204040 216003 204096
rect 114461 204038 216003 204040
rect 114461 204035 114527 204038
rect 215937 204035 216003 204038
rect 195329 203554 195395 203557
rect 318793 203554 318859 203557
rect 195329 203552 318859 203554
rect 195329 203496 195334 203552
rect 195390 203496 318798 203552
rect 318854 203496 318859 203552
rect 195329 203494 318859 203496
rect 195329 203491 195395 203494
rect 318793 203491 318859 203494
rect 213729 203010 213795 203013
rect 583569 203010 583635 203013
rect 213729 203008 583635 203010
rect 213729 202952 213734 203008
rect 213790 202952 583574 203008
rect 583630 202952 583635 203008
rect 213729 202950 583635 202952
rect 213729 202947 213795 202950
rect 583569 202947 583635 202950
rect 66161 202874 66227 202877
rect 233509 202874 233575 202877
rect 66161 202872 233575 202874
rect 66161 202816 66166 202872
rect 66222 202816 233514 202872
rect 233570 202816 233575 202872
rect 66161 202814 233575 202816
rect 66161 202811 66227 202814
rect 233509 202811 233575 202814
rect 129641 202330 129707 202333
rect 195329 202330 195395 202333
rect 129641 202328 195395 202330
rect 129641 202272 129646 202328
rect 129702 202272 195334 202328
rect 195390 202272 195395 202328
rect 129641 202270 195395 202272
rect 129641 202267 129707 202270
rect 195329 202267 195395 202270
rect 304257 202330 304323 202333
rect 309174 202330 309180 202332
rect 304257 202328 309180 202330
rect 304257 202272 304262 202328
rect 304318 202272 309180 202328
rect 304257 202270 309180 202272
rect 304257 202267 304323 202270
rect 309174 202268 309180 202270
rect 309244 202268 309250 202332
rect 118601 202194 118667 202197
rect 193857 202194 193923 202197
rect 118601 202192 193923 202194
rect 118601 202136 118606 202192
rect 118662 202136 193862 202192
rect 193918 202136 193923 202192
rect 118601 202134 193923 202136
rect 118601 202131 118667 202134
rect 193857 202131 193923 202134
rect 199469 202194 199535 202197
rect 307937 202194 308003 202197
rect 199469 202192 308003 202194
rect 199469 202136 199474 202192
rect 199530 202136 307942 202192
rect 307998 202136 308003 202192
rect 199469 202134 308003 202136
rect 199469 202131 199535 202134
rect 307937 202131 308003 202134
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 85481 200970 85547 200973
rect 167821 200970 167887 200973
rect 85481 200968 167887 200970
rect 85481 200912 85486 200968
rect 85542 200912 167826 200968
rect 167882 200912 167887 200968
rect 85481 200910 167887 200912
rect 85481 200907 85547 200910
rect 167821 200907 167887 200910
rect 102041 200834 102107 200837
rect 245653 200834 245719 200837
rect 102041 200832 245719 200834
rect 102041 200776 102046 200832
rect 102102 200776 245658 200832
rect 245714 200776 245719 200832
rect 102041 200774 245719 200776
rect 102041 200771 102107 200774
rect 245653 200771 245719 200774
rect 162117 200698 162183 200701
rect 329833 200698 329899 200701
rect 162117 200696 329899 200698
rect 162117 200640 162122 200696
rect 162178 200640 329838 200696
rect 329894 200640 329899 200696
rect 162117 200638 329899 200640
rect 162117 200635 162183 200638
rect 329833 200635 329899 200638
rect 315941 200156 316007 200157
rect 315941 200154 315988 200156
rect 315896 200152 315988 200154
rect 316052 200154 316058 200156
rect 315896 200096 315946 200152
rect 315896 200094 315988 200096
rect 315941 200092 315988 200094
rect 316052 200094 316134 200154
rect 316052 200092 316058 200094
rect 315941 200091 316007 200092
rect 63217 200018 63283 200021
rect 211797 200018 211863 200021
rect 315941 200018 316007 200021
rect 63217 200016 211863 200018
rect 63217 199960 63222 200016
rect 63278 199960 211802 200016
rect 211858 199960 211863 200016
rect 63217 199958 211863 199960
rect 315896 200016 316050 200018
rect 315896 199960 315946 200016
rect 316002 199960 316050 200016
rect 315896 199958 316050 199960
rect 63217 199955 63283 199958
rect 211797 199955 211863 199958
rect 315941 199955 316050 199958
rect 315990 199884 316050 199955
rect 315982 199820 315988 199884
rect 316052 199820 316058 199884
rect 222929 199474 222995 199477
rect 281758 199474 281764 199476
rect 222929 199472 281764 199474
rect 222929 199416 222934 199472
rect 222990 199416 281764 199472
rect 222929 199414 281764 199416
rect 222929 199411 222995 199414
rect 281758 199412 281764 199414
rect 281828 199412 281834 199476
rect 95141 199338 95207 199341
rect 351913 199338 351979 199341
rect 95141 199336 351979 199338
rect 95141 199280 95146 199336
rect 95202 199280 351918 199336
rect 351974 199280 351979 199336
rect 95141 199278 351979 199280
rect 95141 199275 95207 199278
rect 351913 199275 351979 199278
rect 54937 198658 55003 198661
rect 220077 198658 220143 198661
rect 54937 198656 220143 198658
rect 54937 198600 54942 198656
rect 54998 198600 220082 198656
rect 220138 198600 220143 198656
rect 54937 198598 220143 198600
rect 54937 198595 55003 198598
rect 220077 198595 220143 198598
rect 133689 198114 133755 198117
rect 184289 198114 184355 198117
rect 133689 198112 184355 198114
rect 133689 198056 133694 198112
rect 133750 198056 184294 198112
rect 184350 198056 184355 198112
rect 133689 198054 184355 198056
rect 133689 198051 133755 198054
rect 184289 198051 184355 198054
rect 36537 197978 36603 197981
rect 150382 197978 150388 197980
rect 36537 197976 150388 197978
rect 36537 197920 36542 197976
rect 36598 197920 150388 197976
rect 36537 197918 150388 197920
rect 36537 197915 36603 197918
rect 150382 197916 150388 197918
rect 150452 197916 150458 197980
rect 159214 197916 159220 197980
rect 159284 197978 159290 197980
rect 168414 197978 168420 197980
rect 159284 197918 168420 197978
rect 159284 197916 159290 197918
rect 168414 197916 168420 197918
rect 168484 197916 168490 197980
rect 197261 197978 197327 197981
rect 271965 197978 272031 197981
rect 197261 197976 272031 197978
rect 197261 197920 197266 197976
rect 197322 197920 271970 197976
rect 272026 197920 272031 197976
rect 197261 197918 272031 197920
rect 197261 197915 197327 197918
rect 271965 197915 272031 197918
rect 188429 196754 188495 196757
rect 285806 196754 285812 196756
rect 188429 196752 285812 196754
rect 188429 196696 188434 196752
rect 188490 196696 285812 196752
rect 188429 196694 285812 196696
rect 188429 196691 188495 196694
rect 285806 196692 285812 196694
rect 285876 196692 285882 196756
rect 73061 196618 73127 196621
rect 358813 196618 358879 196621
rect 73061 196616 358879 196618
rect 73061 196560 73066 196616
rect 73122 196560 358818 196616
rect 358874 196560 358879 196616
rect 73061 196558 358879 196560
rect 73061 196555 73127 196558
rect 358813 196555 358879 196558
rect 139209 195938 139275 195941
rect 242934 195938 242940 195940
rect 139209 195936 242940 195938
rect 139209 195880 139214 195936
rect 139270 195880 242940 195936
rect 139209 195878 242940 195880
rect 139209 195875 139275 195878
rect 242934 195876 242940 195878
rect 243004 195876 243010 195940
rect 214649 195394 214715 195397
rect 285622 195394 285628 195396
rect 214649 195392 285628 195394
rect 214649 195336 214654 195392
rect 214710 195336 285628 195392
rect 214649 195334 285628 195336
rect 214649 195331 214715 195334
rect 285622 195332 285628 195334
rect 285692 195332 285698 195396
rect 88241 195258 88307 195261
rect 322197 195258 322263 195261
rect 88241 195256 322263 195258
rect 88241 195200 88246 195256
rect 88302 195200 322202 195256
rect 322258 195200 322263 195256
rect 88241 195198 322263 195200
rect 88241 195195 88307 195198
rect 322197 195195 322263 195198
rect 241278 194108 241284 194172
rect 241348 194170 241354 194172
rect 271873 194170 271939 194173
rect 241348 194168 271939 194170
rect 241348 194112 271878 194168
rect 271934 194112 271939 194168
rect 241348 194110 271939 194112
rect 241348 194108 241354 194110
rect 271873 194107 271939 194110
rect 213821 194034 213887 194037
rect 265750 194034 265756 194036
rect 213821 194032 265756 194034
rect 213821 193976 213826 194032
rect 213882 193976 265756 194032
rect 213821 193974 265756 193976
rect 213821 193971 213887 193974
rect 265750 193972 265756 193974
rect 265820 193972 265826 194036
rect 133781 193898 133847 193901
rect 309726 193898 309732 193900
rect 133781 193896 309732 193898
rect 133781 193840 133786 193896
rect 133842 193840 309732 193896
rect 133781 193838 309732 193840
rect 133781 193835 133847 193838
rect 309726 193836 309732 193838
rect 309796 193836 309802 193900
rect 61837 193218 61903 193221
rect 266353 193220 266419 193221
rect 266302 193218 266308 193220
rect 61837 193216 266308 193218
rect 266372 193216 266419 193220
rect 61837 193160 61842 193216
rect 61898 193160 266308 193216
rect 266414 193160 266419 193216
rect 61837 193158 266308 193160
rect 61837 193155 61903 193158
rect 266302 193156 266308 193158
rect 266372 193156 266419 193160
rect 266353 193155 266419 193156
rect 583661 193082 583727 193085
rect 583526 193080 583727 193082
rect 583526 193024 583666 193080
rect 583722 193024 583727 193080
rect 583526 193022 583727 193024
rect 188286 192612 188292 192676
rect 188356 192674 188362 192676
rect 240777 192674 240843 192677
rect 583526 192674 583586 193022
rect 583661 193019 583727 193022
rect 188356 192672 240843 192674
rect 188356 192616 240782 192672
rect 240838 192616 240843 192672
rect 188356 192614 240843 192616
rect 188356 192612 188362 192614
rect 240777 192611 240843 192614
rect 583342 192628 583586 192674
rect 583342 192614 584960 192628
rect 83958 192476 83964 192540
rect 84028 192538 84034 192540
rect 189717 192538 189783 192541
rect 84028 192536 189783 192538
rect 84028 192480 189722 192536
rect 189778 192480 189783 192536
rect 84028 192478 189783 192480
rect 84028 192476 84034 192478
rect 189717 192475 189783 192478
rect 218697 192538 218763 192541
rect 281574 192538 281580 192540
rect 218697 192536 281580 192538
rect 218697 192480 218702 192536
rect 218758 192480 281580 192536
rect 218697 192478 281580 192480
rect 218697 192475 218763 192478
rect 281574 192476 281580 192478
rect 281644 192476 281650 192540
rect 583342 192538 583402 192614
rect 583520 192538 584960 192614
rect 583342 192478 584960 192538
rect 583520 192388 584960 192478
rect 151721 191042 151787 191045
rect 320173 191042 320239 191045
rect 151721 191040 320239 191042
rect 151721 190984 151726 191040
rect 151782 190984 320178 191040
rect 320234 190984 320239 191040
rect 151721 190982 320239 190984
rect 151721 190979 151787 190982
rect 320173 190979 320239 190982
rect 250713 190634 250779 190637
rect 280286 190634 280292 190636
rect 250713 190632 280292 190634
rect 250713 190576 250718 190632
rect 250774 190576 280292 190632
rect 250713 190574 280292 190576
rect 250713 190571 250779 190574
rect 280286 190572 280292 190574
rect 280356 190572 280362 190636
rect 218421 190498 218487 190501
rect 315941 190500 316007 190501
rect 304942 190498 304948 190500
rect 218421 190496 304948 190498
rect 218421 190440 218426 190496
rect 218482 190440 304948 190496
rect 218421 190438 304948 190440
rect 218421 190435 218487 190438
rect 304942 190436 304948 190438
rect 305012 190436 305018 190500
rect 315941 190498 315988 190500
rect 315896 190496 315988 190498
rect 316052 190498 316058 190500
rect 315896 190440 315946 190496
rect 315896 190438 315988 190440
rect 315941 190436 315988 190438
rect 316052 190438 316134 190498
rect 316052 190436 316058 190438
rect 315941 190435 316007 190436
rect 315941 190364 316007 190365
rect 315941 190362 315988 190364
rect 315896 190360 315988 190362
rect 316052 190362 316058 190364
rect 315896 190304 315946 190360
rect 315896 190302 315988 190304
rect 315941 190300 315988 190302
rect 316052 190302 316134 190362
rect 316052 190300 316058 190302
rect 315941 190299 316007 190300
rect 133086 189892 133092 189956
rect 133156 189954 133162 189956
rect 228357 189954 228423 189957
rect 133156 189952 228423 189954
rect 133156 189896 228362 189952
rect 228418 189896 228423 189952
rect 133156 189894 228423 189896
rect 133156 189892 133162 189894
rect 228357 189891 228423 189894
rect 143390 189756 143396 189820
rect 143460 189818 143466 189820
rect 241513 189818 241579 189821
rect 143460 189816 241579 189818
rect 143460 189760 241518 189816
rect 241574 189760 241579 189816
rect 143460 189758 241579 189760
rect 143460 189756 143466 189758
rect 241513 189755 241579 189758
rect 258717 189818 258783 189821
rect 301681 189818 301747 189821
rect 258717 189816 301747 189818
rect 258717 189760 258722 189816
rect 258778 189760 301686 189816
rect 301742 189760 301747 189816
rect 258717 189758 301747 189760
rect 258717 189755 258783 189758
rect 301681 189755 301747 189758
rect 89621 189682 89687 189685
rect 275134 189682 275140 189684
rect 89621 189680 275140 189682
rect 89621 189624 89626 189680
rect 89682 189624 275140 189680
rect 89621 189622 275140 189624
rect 89621 189619 89687 189622
rect 275134 189620 275140 189622
rect 275204 189620 275210 189684
rect 291837 189682 291903 189685
rect 312302 189682 312308 189684
rect 291837 189680 312308 189682
rect 291837 189624 291842 189680
rect 291898 189624 312308 189680
rect 291837 189622 312308 189624
rect 291837 189619 291903 189622
rect 312302 189620 312308 189622
rect 312372 189620 312378 189684
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 111701 188458 111767 188461
rect 186957 188458 187023 188461
rect 111701 188456 187023 188458
rect 111701 188400 111706 188456
rect 111762 188400 186962 188456
rect 187018 188400 187023 188456
rect 111701 188398 187023 188400
rect 111701 188395 111767 188398
rect 186957 188395 187023 188398
rect 197169 188458 197235 188461
rect 272558 188458 272564 188460
rect 197169 188456 272564 188458
rect 197169 188400 197174 188456
rect 197230 188400 272564 188456
rect 197169 188398 272564 188400
rect 197169 188395 197235 188398
rect 272558 188396 272564 188398
rect 272628 188396 272634 188460
rect 302877 188458 302943 188461
rect 316166 188458 316172 188460
rect 302877 188456 316172 188458
rect 302877 188400 302882 188456
rect 302938 188400 316172 188456
rect 302877 188398 316172 188400
rect 302877 188395 302943 188398
rect 316166 188396 316172 188398
rect 316236 188396 316242 188460
rect 81341 188322 81407 188325
rect 313222 188322 313228 188324
rect 81341 188320 313228 188322
rect 81341 188264 81346 188320
rect 81402 188264 313228 188320
rect 81341 188262 313228 188264
rect 81341 188259 81407 188262
rect 313222 188260 313228 188262
rect 313292 188260 313298 188324
rect 160737 187098 160803 187101
rect 173157 187098 173223 187101
rect 160737 187096 173223 187098
rect 160737 187040 160742 187096
rect 160798 187040 173162 187096
rect 173218 187040 173223 187096
rect 160737 187038 173223 187040
rect 160737 187035 160803 187038
rect 173157 187035 173223 187038
rect 182081 187098 182147 187101
rect 278865 187098 278931 187101
rect 182081 187096 278931 187098
rect 182081 187040 182086 187096
rect 182142 187040 278870 187096
rect 278926 187040 278931 187096
rect 182081 187038 278931 187040
rect 182081 187035 182147 187038
rect 278865 187035 278931 187038
rect 93761 186962 93827 186965
rect 202229 186962 202295 186965
rect 93761 186960 202295 186962
rect 93761 186904 93766 186960
rect 93822 186904 202234 186960
rect 202290 186904 202295 186960
rect 93761 186902 202295 186904
rect 93761 186899 93827 186902
rect 202229 186899 202295 186902
rect 209037 186962 209103 186965
rect 327349 186962 327415 186965
rect 209037 186960 327415 186962
rect 209037 186904 209042 186960
rect 209098 186904 327354 186960
rect 327410 186904 327415 186960
rect 209037 186902 327415 186904
rect 209037 186899 209103 186902
rect 327349 186899 327415 186902
rect 256049 185874 256115 185877
rect 267774 185874 267780 185876
rect 256049 185872 267780 185874
rect 256049 185816 256054 185872
rect 256110 185816 267780 185872
rect 256049 185814 267780 185816
rect 256049 185811 256115 185814
rect 267774 185812 267780 185814
rect 267844 185812 267850 185876
rect 237230 185676 237236 185740
rect 237300 185738 237306 185740
rect 302325 185738 302391 185741
rect 237300 185736 302391 185738
rect 237300 185680 302330 185736
rect 302386 185680 302391 185736
rect 237300 185678 302391 185680
rect 237300 185676 237306 185678
rect 302325 185675 302391 185678
rect 79961 185602 80027 185605
rect 288934 185602 288940 185604
rect 79961 185600 288940 185602
rect 79961 185544 79966 185600
rect 80022 185544 288940 185600
rect 79961 185542 288940 185544
rect 79961 185539 80027 185542
rect 288934 185540 288940 185542
rect 289004 185540 289010 185604
rect 189809 184378 189875 184381
rect 244273 184378 244339 184381
rect 189809 184376 244339 184378
rect 189809 184320 189814 184376
rect 189870 184320 244278 184376
rect 244334 184320 244339 184376
rect 189809 184318 244339 184320
rect 189809 184315 189875 184318
rect 244273 184315 244339 184318
rect 258809 184378 258875 184381
rect 285765 184378 285831 184381
rect 258809 184376 285831 184378
rect 258809 184320 258814 184376
rect 258870 184320 285770 184376
rect 285826 184320 285831 184376
rect 258809 184318 285831 184320
rect 258809 184315 258875 184318
rect 285765 184315 285831 184318
rect 206921 184242 206987 184245
rect 324497 184242 324563 184245
rect 206921 184240 324563 184242
rect 206921 184184 206926 184240
rect 206982 184184 324502 184240
rect 324558 184184 324563 184240
rect 206921 184182 324563 184184
rect 206921 184179 206987 184182
rect 324497 184179 324563 184182
rect 104801 183834 104867 183837
rect 177481 183834 177547 183837
rect 104801 183832 177547 183834
rect 104801 183776 104806 183832
rect 104862 183776 177486 183832
rect 177542 183776 177547 183832
rect 104801 183774 177547 183776
rect 104801 183771 104867 183774
rect 177481 183771 177547 183774
rect 101949 183698 102015 183701
rect 188429 183698 188495 183701
rect 101949 183696 188495 183698
rect 101949 183640 101954 183696
rect 102010 183640 188434 183696
rect 188490 183640 188495 183696
rect 101949 183638 188495 183640
rect 101949 183635 102015 183638
rect 188429 183635 188495 183638
rect 193029 183154 193095 183157
rect 227713 183154 227779 183157
rect 193029 183152 227779 183154
rect 193029 183096 193034 183152
rect 193090 183096 227718 183152
rect 227774 183096 227779 183152
rect 193029 183094 227779 183096
rect 193029 183091 193095 183094
rect 227713 183091 227779 183094
rect 206277 183018 206343 183021
rect 267917 183018 267983 183021
rect 206277 183016 267983 183018
rect 206277 182960 206282 183016
rect 206338 182960 267922 183016
rect 267978 182960 267983 183016
rect 206277 182958 267983 182960
rect 206277 182955 206343 182958
rect 267917 182955 267983 182958
rect 304257 183018 304323 183021
rect 314929 183018 314995 183021
rect 304257 183016 314995 183018
rect 304257 182960 304262 183016
rect 304318 182960 314934 183016
rect 314990 182960 314995 183016
rect 304257 182958 314995 182960
rect 304257 182955 304323 182958
rect 314929 182955 314995 182958
rect 226977 182882 227043 182885
rect 307845 182882 307911 182885
rect 226977 182880 307911 182882
rect 226977 182824 226982 182880
rect 227038 182824 307850 182880
rect 307906 182824 307911 182880
rect 226977 182822 307911 182824
rect 226977 182819 227043 182822
rect 307845 182819 307911 182822
rect 99465 182202 99531 182205
rect 176009 182202 176075 182205
rect 99465 182200 176075 182202
rect 99465 182144 99470 182200
rect 99526 182144 176014 182200
rect 176070 182144 176075 182200
rect 99465 182142 176075 182144
rect 99465 182139 99531 182142
rect 176009 182139 176075 182142
rect 297357 181522 297423 181525
rect 320449 181522 320515 181525
rect 297357 181520 320515 181522
rect 297357 181464 297362 181520
rect 297418 181464 320454 181520
rect 320510 181464 320515 181520
rect 297357 181462 320515 181464
rect 297357 181459 297423 181462
rect 320449 181459 320515 181462
rect 216438 181324 216444 181388
rect 216508 181386 216514 181388
rect 302366 181386 302372 181388
rect 216508 181326 302372 181386
rect 216508 181324 216514 181326
rect 302366 181324 302372 181326
rect 302436 181324 302442 181388
rect 107469 180978 107535 180981
rect 167729 180978 167795 180981
rect 107469 180976 167795 180978
rect 107469 180920 107474 180976
rect 107530 180920 167734 180976
rect 167790 180920 167795 180976
rect 107469 180918 167795 180920
rect 107469 180915 107535 180918
rect 167729 180915 167795 180918
rect 315982 180916 315988 180980
rect 316052 180916 316058 180980
rect 315990 180845 316050 180916
rect 116945 180842 117011 180845
rect 238109 180842 238175 180845
rect 116945 180840 238175 180842
rect 116945 180784 116950 180840
rect 117006 180784 238114 180840
rect 238170 180784 238175 180840
rect 116945 180782 238175 180784
rect 116945 180779 117011 180782
rect 238109 180779 238175 180782
rect 258073 180842 258139 180845
rect 267958 180842 267964 180844
rect 258073 180840 267964 180842
rect 258073 180784 258078 180840
rect 258134 180784 267964 180840
rect 258073 180782 267964 180784
rect 258073 180779 258139 180782
rect 267958 180780 267964 180782
rect 268028 180780 268034 180844
rect 315941 180842 316050 180845
rect 315896 180840 316050 180842
rect 315896 180784 315946 180840
rect 316002 180784 316050 180840
rect 315896 180782 316050 180784
rect 315941 180779 316007 180782
rect 315941 180708 316007 180709
rect 315941 180706 315988 180708
rect 315896 180704 315988 180706
rect 316052 180706 316058 180708
rect 315896 180648 315946 180704
rect 315896 180646 315988 180648
rect 315941 180644 315988 180646
rect 316052 180646 316134 180706
rect 316052 180644 316058 180646
rect 315941 180643 316007 180644
rect 232589 180162 232655 180165
rect 305126 180162 305132 180164
rect 232589 180160 305132 180162
rect 232589 180104 232594 180160
rect 232650 180104 305132 180160
rect 232589 180102 305132 180104
rect 232589 180099 232655 180102
rect 305126 180100 305132 180102
rect 305196 180100 305202 180164
rect 191741 180026 191807 180029
rect 280286 180026 280292 180028
rect 191741 180024 280292 180026
rect 191741 179968 191746 180024
rect 191802 179968 280292 180024
rect 191741 179966 280292 179968
rect 191741 179963 191807 179966
rect 280286 179964 280292 179966
rect 280356 179964 280362 180028
rect 295977 180026 296043 180029
rect 301814 180026 301820 180028
rect 295977 180024 301820 180026
rect 295977 179968 295982 180024
rect 296038 179968 301820 180024
rect 295977 179966 301820 179968
rect 295977 179963 296043 179966
rect 301814 179964 301820 179966
rect 301884 179964 301890 180028
rect 304441 180026 304507 180029
rect 323209 180026 323275 180029
rect 304441 180024 323275 180026
rect 304441 179968 304446 180024
rect 304502 179968 323214 180024
rect 323270 179968 323275 180024
rect 304441 179966 323275 179968
rect 304441 179963 304507 179966
rect 323209 179963 323275 179966
rect 112253 179618 112319 179621
rect 182909 179618 182975 179621
rect 112253 179616 182975 179618
rect 112253 179560 112258 179616
rect 112314 179560 182914 179616
rect 182970 179560 182975 179616
rect 112253 179558 182975 179560
rect 112253 179555 112319 179558
rect 182909 179555 182975 179558
rect 105445 179482 105511 179485
rect 249057 179482 249123 179485
rect 105445 179480 249123 179482
rect 105445 179424 105450 179480
rect 105506 179424 249062 179480
rect 249118 179424 249123 179480
rect 105445 179422 249123 179424
rect 105445 179419 105511 179422
rect 249057 179419 249123 179422
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 204897 178666 204963 178669
rect 308622 178666 308628 178668
rect 204897 178664 308628 178666
rect 204897 178608 204902 178664
rect 204958 178608 308628 178664
rect 204897 178606 308628 178608
rect 204897 178603 204963 178606
rect 308622 178604 308628 178606
rect 308692 178604 308698 178668
rect 110638 178196 110644 178260
rect 110708 178258 110714 178260
rect 171869 178258 171935 178261
rect 110708 178256 171935 178258
rect 110708 178200 171874 178256
rect 171930 178200 171935 178256
rect 110708 178198 171935 178200
rect 110708 178196 110714 178198
rect 171869 178195 171935 178198
rect 259361 178258 259427 178261
rect 263910 178258 263916 178260
rect 259361 178256 263916 178258
rect 259361 178200 259366 178256
rect 259422 178200 263916 178256
rect 259361 178198 263916 178200
rect 259361 178195 259427 178198
rect 263910 178196 263916 178198
rect 263980 178196 263986 178260
rect 220077 178122 220143 178125
rect 97030 178120 220143 178122
rect 97030 178064 220082 178120
rect 220138 178064 220143 178120
rect 97030 178062 220143 178064
rect 97030 177988 97090 178062
rect 220077 178059 220143 178062
rect 250529 178122 250595 178125
rect 290590 178122 290596 178124
rect 250529 178120 290596 178122
rect 250529 178064 250534 178120
rect 250590 178064 290596 178120
rect 250529 178062 290596 178064
rect 250529 178059 250595 178062
rect 290590 178060 290596 178062
rect 290660 178060 290666 178124
rect 297449 178122 297515 178125
rect 302509 178122 302575 178125
rect 297449 178120 302575 178122
rect 297449 178064 297454 178120
rect 297510 178064 302514 178120
rect 302570 178064 302575 178120
rect 297449 178062 302575 178064
rect 297449 178059 297515 178062
rect 302509 178059 302575 178062
rect 97022 177924 97028 177988
rect 97092 177924 97098 177988
rect 216029 177986 216095 177989
rect 259361 177986 259427 177989
rect 216029 177984 259427 177986
rect 216029 177928 216034 177984
rect 216090 177928 259366 177984
rect 259422 177928 259427 177984
rect 216029 177926 259427 177928
rect 216029 177923 216095 177926
rect 259361 177923 259427 177926
rect 100702 177516 100708 177580
rect 100772 177578 100778 177580
rect 101949 177578 102015 177581
rect 100772 177576 102015 177578
rect 100772 177520 101954 177576
rect 102010 177520 102015 177576
rect 100772 177518 102015 177520
rect 100772 177516 100778 177518
rect 101949 177515 102015 177518
rect 104566 177516 104572 177580
rect 104636 177578 104642 177580
rect 104801 177578 104867 177581
rect 104636 177576 104867 177578
rect 104636 177520 104806 177576
rect 104862 177520 104867 177576
rect 104636 177518 104867 177520
rect 104636 177516 104642 177518
rect 104801 177515 104867 177518
rect 105670 177516 105676 177580
rect 105740 177578 105746 177580
rect 106181 177578 106247 177581
rect 105740 177576 106247 177578
rect 105740 177520 106186 177576
rect 106242 177520 106247 177576
rect 105740 177518 106247 177520
rect 105740 177516 105746 177518
rect 106181 177515 106247 177518
rect 106958 177516 106964 177580
rect 107028 177578 107034 177580
rect 107469 177578 107535 177581
rect 107028 177576 107535 177578
rect 107028 177520 107474 177576
rect 107530 177520 107535 177576
rect 107028 177518 107535 177520
rect 107028 177516 107034 177518
rect 107469 177515 107535 177518
rect 113214 177516 113220 177580
rect 113284 177578 113290 177580
rect 113725 177578 113791 177581
rect 116945 177580 117011 177581
rect 116894 177578 116900 177580
rect 113284 177576 113791 177578
rect 113284 177520 113730 177576
rect 113786 177520 113791 177576
rect 113284 177518 113791 177520
rect 116854 177518 116900 177578
rect 116964 177576 117011 177580
rect 117006 177520 117011 177576
rect 113284 177516 113290 177518
rect 113725 177515 113791 177518
rect 116894 177516 116900 177518
rect 116964 177516 117011 177520
rect 119470 177516 119476 177580
rect 119540 177578 119546 177580
rect 119981 177578 120047 177581
rect 119540 177576 120047 177578
rect 119540 177520 119986 177576
rect 120042 177520 120047 177576
rect 119540 177518 120047 177520
rect 119540 177516 119546 177518
rect 116945 177515 117011 177516
rect 119981 177515 120047 177518
rect 120758 177516 120764 177580
rect 120828 177578 120834 177580
rect 121361 177578 121427 177581
rect 120828 177576 121427 177578
rect 120828 177520 121366 177576
rect 121422 177520 121427 177576
rect 120828 177518 121427 177520
rect 120828 177516 120834 177518
rect 121361 177515 121427 177518
rect 125726 177516 125732 177580
rect 125796 177578 125802 177580
rect 126053 177578 126119 177581
rect 125796 177576 126119 177578
rect 125796 177520 126058 177576
rect 126114 177520 126119 177576
rect 125796 177518 126119 177520
rect 125796 177516 125802 177518
rect 126053 177515 126119 177518
rect 129406 177516 129412 177580
rect 129476 177578 129482 177580
rect 129641 177578 129707 177581
rect 129476 177576 129707 177578
rect 129476 177520 129646 177576
rect 129702 177520 129707 177576
rect 129476 177518 129707 177520
rect 129476 177516 129482 177518
rect 129641 177515 129707 177518
rect 148174 177516 148180 177580
rect 148244 177578 148250 177580
rect 148961 177578 149027 177581
rect 148244 177576 149027 177578
rect 148244 177520 148966 177576
rect 149022 177520 149027 177576
rect 148244 177518 149027 177520
rect 148244 177516 148250 177518
rect 148961 177515 149027 177518
rect 258206 177516 258212 177580
rect 258276 177578 258282 177580
rect 264145 177578 264211 177581
rect 258276 177576 264211 177578
rect 258276 177520 264150 177576
rect 264206 177520 264211 177576
rect 258276 177518 264211 177520
rect 258276 177516 258282 177518
rect 264145 177515 264211 177518
rect 260097 177442 260163 177445
rect 270677 177442 270743 177445
rect 260097 177440 270743 177442
rect 260097 177384 260102 177440
rect 260158 177384 270682 177440
rect 270738 177384 270743 177440
rect 260097 177382 270743 177384
rect 260097 177379 260163 177382
rect 270677 177379 270743 177382
rect 294597 177442 294663 177445
rect 301262 177442 301268 177444
rect 294597 177440 301268 177442
rect 294597 177384 294602 177440
rect 294658 177384 301268 177440
rect 294597 177382 301268 177384
rect 294597 177379 294663 177382
rect 301262 177380 301268 177382
rect 301332 177380 301338 177444
rect 191189 177306 191255 177309
rect 264881 177306 264947 177309
rect 191189 177304 264947 177306
rect 191189 177248 191194 177304
rect 191250 177248 264886 177304
rect 264942 177248 264947 177304
rect 191189 177246 264947 177248
rect 191189 177243 191255 177246
rect 264881 177243 264947 177246
rect 291929 177306 291995 177309
rect 309317 177306 309383 177309
rect 291929 177304 309383 177306
rect 291929 177248 291934 177304
rect 291990 177248 309322 177304
rect 309378 177248 309383 177304
rect 291929 177246 309383 177248
rect 291929 177243 291995 177246
rect 309317 177243 309383 177246
rect 112110 177108 112116 177172
rect 112180 177170 112186 177172
rect 112253 177170 112319 177173
rect 112180 177168 112319 177170
rect 112180 177112 112258 177168
rect 112314 177112 112319 177168
rect 112180 177110 112319 177112
rect 112180 177108 112186 177110
rect 112253 177107 112319 177110
rect 118366 177108 118372 177172
rect 118436 177170 118442 177172
rect 118509 177170 118575 177173
rect 118436 177168 118575 177170
rect 118436 177112 118514 177168
rect 118570 177112 118575 177168
rect 118436 177110 118575 177112
rect 118436 177108 118442 177110
rect 118509 177107 118575 177110
rect 108062 176972 108068 177036
rect 108132 177034 108138 177036
rect 238017 177034 238083 177037
rect 108132 177032 238083 177034
rect 108132 176976 238022 177032
rect 238078 176976 238083 177032
rect 108132 176974 238083 176976
rect 108132 176972 108138 176974
rect 238017 176971 238083 176974
rect 98310 176836 98316 176900
rect 98380 176898 98386 176900
rect 166349 176898 166415 176901
rect 98380 176896 166415 176898
rect 98380 176840 166354 176896
rect 166410 176840 166415 176896
rect 98380 176838 166415 176840
rect 98380 176836 98386 176838
rect 166349 176835 166415 176838
rect 264329 176898 264395 176901
rect 274817 176898 274883 176901
rect 264329 176896 274883 176898
rect 264329 176840 264334 176896
rect 264390 176840 274822 176896
rect 274878 176840 274883 176896
rect 264329 176838 274883 176840
rect 264329 176835 264395 176838
rect 274817 176835 274883 176838
rect 99465 176762 99531 176765
rect 102041 176764 102107 176765
rect 101990 176762 101996 176764
rect 99422 176760 99531 176762
rect 99422 176704 99470 176760
rect 99526 176704 99531 176760
rect 99422 176699 99531 176704
rect 101950 176702 101996 176762
rect 102060 176760 102107 176764
rect 103329 176762 103395 176765
rect 115841 176764 115907 176765
rect 124489 176764 124555 176765
rect 115790 176762 115796 176764
rect 102102 176704 102107 176760
rect 101990 176700 101996 176702
rect 102060 176700 102107 176704
rect 102041 176699 102107 176700
rect 103286 176760 103395 176762
rect 103286 176704 103334 176760
rect 103390 176704 103395 176760
rect 103286 176699 103395 176704
rect 115750 176702 115796 176762
rect 115860 176760 115907 176764
rect 124438 176762 124444 176764
rect 115902 176704 115907 176760
rect 115790 176700 115796 176702
rect 115860 176700 115907 176704
rect 124398 176702 124444 176762
rect 124508 176760 124555 176764
rect 124550 176704 124555 176760
rect 124438 176700 124444 176702
rect 124508 176700 124555 176704
rect 127014 176700 127020 176764
rect 127084 176762 127090 176764
rect 127617 176762 127683 176765
rect 132401 176764 132467 176765
rect 134425 176764 134491 176765
rect 136081 176764 136147 176765
rect 132350 176762 132356 176764
rect 127084 176760 127683 176762
rect 127084 176704 127622 176760
rect 127678 176704 127683 176760
rect 127084 176702 127683 176704
rect 132310 176702 132356 176762
rect 132420 176760 132467 176764
rect 134374 176762 134380 176764
rect 132462 176704 132467 176760
rect 127084 176700 127090 176702
rect 115841 176699 115907 176700
rect 124489 176699 124555 176700
rect 127617 176699 127683 176702
rect 132350 176700 132356 176702
rect 132420 176700 132467 176704
rect 134334 176702 134380 176762
rect 134444 176760 134491 176764
rect 136030 176762 136036 176764
rect 134486 176704 134491 176760
rect 134374 176700 134380 176702
rect 134444 176700 134491 176704
rect 135990 176702 136036 176762
rect 136100 176760 136147 176764
rect 136142 176704 136147 176760
rect 136030 176700 136036 176702
rect 136100 176700 136147 176704
rect 158846 176700 158852 176764
rect 158916 176762 158922 176764
rect 158989 176762 159055 176765
rect 158916 176760 159055 176762
rect 158916 176704 158994 176760
rect 159050 176704 159055 176760
rect 158916 176702 159055 176704
rect 158916 176700 158922 176702
rect 132401 176699 132467 176700
rect 134425 176699 134491 176700
rect 136081 176699 136147 176700
rect 158989 176699 159055 176702
rect 237373 176762 237439 176765
rect 265014 176762 265020 176764
rect 237373 176760 265020 176762
rect 237373 176704 237378 176760
rect 237434 176704 265020 176760
rect 237373 176702 265020 176704
rect 237373 176699 237439 176702
rect 265014 176700 265020 176702
rect 265084 176700 265090 176764
rect 276606 176700 276612 176764
rect 276676 176762 276682 176764
rect 300853 176762 300919 176765
rect 276676 176760 300919 176762
rect 276676 176704 300858 176760
rect 300914 176704 300919 176760
rect 276676 176702 300919 176704
rect 276676 176700 276682 176702
rect 300853 176699 300919 176702
rect 99422 176492 99482 176699
rect 103286 176492 103346 176699
rect 193121 176626 193187 176629
rect 259729 176626 259795 176629
rect 193121 176624 259795 176626
rect 193121 176568 193126 176624
rect 193182 176568 259734 176624
rect 259790 176568 259795 176624
rect 193121 176566 259795 176568
rect 193121 176563 193187 176566
rect 259729 176563 259795 176566
rect 265617 176626 265683 176629
rect 268009 176626 268075 176629
rect 265617 176624 268075 176626
rect 265617 176568 265622 176624
rect 265678 176568 268014 176624
rect 268070 176568 268075 176624
rect 265617 176566 268075 176568
rect 265617 176563 265683 176566
rect 268009 176563 268075 176566
rect 301681 176626 301747 176629
rect 306598 176626 306604 176628
rect 301681 176624 306604 176626
rect 301681 176568 301686 176624
rect 301742 176568 306604 176624
rect 301681 176566 306604 176568
rect 301681 176563 301747 176566
rect 306598 176564 306604 176566
rect 306668 176564 306674 176628
rect 99414 176428 99420 176492
rect 99484 176428 99490 176492
rect 103278 176428 103284 176492
rect 103348 176428 103354 176492
rect 244917 176490 244983 176493
rect 249701 176490 249767 176493
rect 244917 176488 249767 176490
rect 244917 176432 244922 176488
rect 244978 176432 249706 176488
rect 249762 176432 249767 176488
rect 244917 176430 249767 176432
rect 244917 176427 244983 176430
rect 249701 176427 249767 176430
rect 300853 176082 300919 176085
rect 300853 176080 301330 176082
rect -960 175796 480 176036
rect 300853 176024 300858 176080
rect 300914 176024 301330 176080
rect 300853 176022 301330 176024
rect 300853 176019 300919 176022
rect 261477 175946 261543 175949
rect 265157 175946 265223 175949
rect 298185 175948 298251 175949
rect 298134 175946 298140 175948
rect 261477 175944 265223 175946
rect 261477 175888 261482 175944
rect 261538 175888 265162 175944
rect 265218 175888 265223 175944
rect 261477 175886 265223 175888
rect 298094 175886 298140 175946
rect 298204 175944 298251 175948
rect 298246 175888 298251 175944
rect 261477 175883 261543 175886
rect 265157 175883 265223 175886
rect 298134 175884 298140 175886
rect 298204 175884 298251 175888
rect 298185 175883 298251 175884
rect 130745 175812 130811 175813
rect 130694 175810 130700 175812
rect 130654 175750 130700 175810
rect 130764 175808 130811 175812
rect 130806 175752 130811 175808
rect 130694 175748 130700 175750
rect 130764 175748 130811 175752
rect 130745 175747 130811 175748
rect 262213 175810 262279 175813
rect 262213 175808 263242 175810
rect 262213 175752 262218 175808
rect 262274 175752 263242 175808
rect 262213 175750 263242 175752
rect 262213 175747 262279 175750
rect 114318 175612 114324 175676
rect 114388 175674 114394 175676
rect 164734 175674 164740 175676
rect 114388 175614 164740 175674
rect 114388 175612 114394 175614
rect 164734 175612 164740 175614
rect 164804 175612 164810 175676
rect 249517 175674 249583 175677
rect 249517 175672 252172 175674
rect 249517 175616 249522 175672
rect 249578 175616 252172 175672
rect 263182 175644 263242 175750
rect 287973 175674 288039 175677
rect 287973 175672 290076 175674
rect 249517 175614 252172 175616
rect 287973 175616 287978 175672
rect 288034 175616 290076 175672
rect 287973 175614 290076 175616
rect 249517 175611 249583 175614
rect 287973 175611 288039 175614
rect 121862 175476 121868 175540
rect 121932 175538 121938 175540
rect 185761 175538 185827 175541
rect 121932 175536 185827 175538
rect 121932 175480 185766 175536
rect 185822 175480 185827 175536
rect 301270 175508 301330 176022
rect 121932 175478 185827 175480
rect 121932 175476 121938 175478
rect 185761 175475 185827 175478
rect 109534 175340 109540 175404
rect 109604 175402 109610 175404
rect 181437 175402 181503 175405
rect 109604 175400 181503 175402
rect 109604 175344 181442 175400
rect 181498 175344 181503 175400
rect 109604 175342 181503 175344
rect 109604 175340 109610 175342
rect 181437 175339 181503 175342
rect 264973 175266 265039 175269
rect 263948 175264 265039 175266
rect 263948 175208 264978 175264
rect 265034 175208 265039 175264
rect 263948 175206 265039 175208
rect 264973 175203 265039 175206
rect 287789 175266 287855 175269
rect 301405 175266 301471 175269
rect 287789 175264 290076 175266
rect 287789 175208 287794 175264
rect 287850 175208 290076 175264
rect 287789 175206 290076 175208
rect 301405 175264 301514 175266
rect 301405 175208 301410 175264
rect 301466 175208 301514 175264
rect 287789 175203 287855 175206
rect 301405 175203 301514 175208
rect 123109 174996 123175 174997
rect 123064 174994 123070 174996
rect 123018 174934 123070 174994
rect 123134 174992 123175 174996
rect 123170 174936 123175 174992
rect 123064 174932 123070 174934
rect 123134 174932 123175 174936
rect 123109 174931 123175 174932
rect 249701 174994 249767 174997
rect 249701 174992 252172 174994
rect 249701 174936 249706 174992
rect 249762 174936 252172 174992
rect 249701 174934 252172 174936
rect 249701 174931 249767 174934
rect 128096 174796 128102 174860
rect 128166 174858 128172 174860
rect 168465 174858 168531 174861
rect 128166 174856 168531 174858
rect 128166 174800 168470 174856
rect 168526 174800 168531 174856
rect 128166 174798 168531 174800
rect 128166 174796 128172 174798
rect 168465 174795 168531 174798
rect 287881 174858 287947 174861
rect 287881 174856 290076 174858
rect 287881 174800 287886 174856
rect 287942 174800 290076 174856
rect 287881 174798 290076 174800
rect 287881 174795 287947 174798
rect 133270 174660 133276 174724
rect 133340 174722 133346 174724
rect 264237 174722 264303 174725
rect 133340 174662 252202 174722
rect 263948 174720 264303 174722
rect 263948 174664 264242 174720
rect 264298 174664 264303 174720
rect 301454 174692 301514 175203
rect 263948 174662 264303 174664
rect 133340 174660 133346 174662
rect 252142 174284 252202 174662
rect 264237 174659 264303 174662
rect 285213 174450 285279 174453
rect 301405 174450 301471 174453
rect 285213 174448 290076 174450
rect 285213 174392 285218 174448
rect 285274 174392 290076 174448
rect 285213 174390 290076 174392
rect 301405 174448 301514 174450
rect 301405 174392 301410 174448
rect 301466 174392 301514 174448
rect 285213 174387 285279 174390
rect 301405 174387 301514 174392
rect 264145 174314 264211 174317
rect 263948 174312 264211 174314
rect 263948 174256 264150 174312
rect 264206 174256 264211 174312
rect 263948 174254 264211 174256
rect 264145 174251 264211 174254
rect 288341 174042 288407 174045
rect 288341 174040 290076 174042
rect 288341 173984 288346 174040
rect 288402 173984 290076 174040
rect 301454 174012 301514 174387
rect 288341 173982 290076 173984
rect 288341 173979 288407 173982
rect 173341 173906 173407 173909
rect 251817 173906 251883 173909
rect 173341 173904 251883 173906
rect 173341 173848 173346 173904
rect 173402 173848 251822 173904
rect 251878 173848 251883 173904
rect 173341 173846 251883 173848
rect 173341 173843 173407 173846
rect 251817 173843 251883 173846
rect 266353 173770 266419 173773
rect 263948 173768 266419 173770
rect 263948 173712 266358 173768
rect 266414 173712 266419 173768
rect 263948 173710 266419 173712
rect 266353 173707 266419 173710
rect 301262 173708 301268 173772
rect 301332 173708 301338 173772
rect 249701 173634 249767 173637
rect 287605 173634 287671 173637
rect 249701 173632 252172 173634
rect 249701 173576 249706 173632
rect 249762 173576 252172 173632
rect 249701 173574 252172 173576
rect 287605 173632 290076 173634
rect 287605 173576 287610 173632
rect 287666 173576 290076 173632
rect 287605 173574 290076 173576
rect 249701 173571 249767 173574
rect 287605 173571 287671 173574
rect 269757 173362 269823 173365
rect 263948 173360 269823 173362
rect 263948 173304 269762 173360
rect 269818 173304 269823 173360
rect 263948 173302 269823 173304
rect 269757 173299 269823 173302
rect 301270 173196 301330 173708
rect 248597 172954 248663 172957
rect 248597 172952 252172 172954
rect 248597 172896 248602 172952
rect 248658 172896 252172 172952
rect 248597 172894 252172 172896
rect 248597 172891 248663 172894
rect 266629 172818 266695 172821
rect 263948 172816 266695 172818
rect 263948 172760 266634 172816
rect 266690 172760 266695 172816
rect 263948 172758 266695 172760
rect 266629 172755 266695 172758
rect 279509 172818 279575 172821
rect 290046 172818 290106 173060
rect 279509 172816 290106 172818
rect 279509 172760 279514 172816
rect 279570 172760 290106 172816
rect 279509 172758 290106 172760
rect 279509 172755 279575 172758
rect 288341 172682 288407 172685
rect 288341 172680 290076 172682
rect 288341 172624 288346 172680
rect 288402 172624 290076 172680
rect 288341 172622 290076 172624
rect 288341 172619 288407 172622
rect 266854 172484 266860 172548
rect 266924 172546 266930 172548
rect 267958 172546 267964 172548
rect 266924 172486 267964 172546
rect 266924 172484 266930 172486
rect 267958 172484 267964 172486
rect 268028 172484 268034 172548
rect 303613 172546 303679 172549
rect 301852 172544 303679 172546
rect 301852 172488 303618 172544
rect 303674 172488 303679 172544
rect 301852 172486 303679 172488
rect 303613 172483 303679 172486
rect 198089 172410 198155 172413
rect 250713 172410 250779 172413
rect 266353 172410 266419 172413
rect 198089 172408 250779 172410
rect 198089 172352 198094 172408
rect 198150 172352 250718 172408
rect 250774 172352 250779 172408
rect 198089 172350 250779 172352
rect 263948 172408 266419 172410
rect 263948 172352 266358 172408
rect 266414 172352 266419 172408
rect 263948 172350 266419 172352
rect 198089 172347 198155 172350
rect 250713 172347 250779 172350
rect 266353 172347 266419 172350
rect 249333 172274 249399 172277
rect 287237 172274 287303 172277
rect 249333 172272 252172 172274
rect 249333 172216 249338 172272
rect 249394 172216 252172 172272
rect 249333 172214 252172 172216
rect 287237 172272 290076 172274
rect 287237 172216 287242 172272
rect 287298 172216 290076 172272
rect 287237 172214 290076 172216
rect 249333 172211 249399 172214
rect 287237 172211 287303 172214
rect 266629 171866 266695 171869
rect 263948 171864 266695 171866
rect 263948 171808 266634 171864
rect 266690 171808 266695 171864
rect 263948 171806 266695 171808
rect 266629 171803 266695 171806
rect 288249 171866 288315 171869
rect 288249 171864 290076 171866
rect 288249 171808 288254 171864
rect 288310 171808 290076 171864
rect 288249 171806 290076 171808
rect 288249 171803 288315 171806
rect 303889 171730 303955 171733
rect 301852 171728 303955 171730
rect 301852 171672 303894 171728
rect 303950 171672 303955 171728
rect 301852 171670 303955 171672
rect 303889 171667 303955 171670
rect 248597 171594 248663 171597
rect 248597 171592 252172 171594
rect 164694 171322 164754 171570
rect 248597 171536 248602 171592
rect 248658 171536 252172 171592
rect 248597 171534 252172 171536
rect 248597 171531 248663 171534
rect 264421 171458 264487 171461
rect 263948 171456 264487 171458
rect 263948 171400 264426 171456
rect 264482 171400 264487 171456
rect 263948 171398 264487 171400
rect 264421 171395 264487 171398
rect 288341 171458 288407 171461
rect 288341 171456 290076 171458
rect 288341 171400 288346 171456
rect 288402 171400 290076 171456
rect 288341 171398 290076 171400
rect 288341 171395 288407 171398
rect 169017 171322 169083 171325
rect 164694 171320 169083 171322
rect 164694 171264 169022 171320
rect 169078 171264 169083 171320
rect 164694 171262 169083 171264
rect 169017 171259 169083 171262
rect 315982 171260 315988 171324
rect 316052 171260 316058 171324
rect 315990 171189 316050 171260
rect 315941 171186 316050 171189
rect 315896 171184 316050 171186
rect 315896 171128 315946 171184
rect 316002 171128 316050 171184
rect 315896 171126 316050 171128
rect 315941 171123 316007 171126
rect 249701 171050 249767 171053
rect 288341 171050 288407 171053
rect 315941 171052 316007 171053
rect 315941 171050 315988 171052
rect 249701 171048 252172 171050
rect 249701 170992 249706 171048
rect 249762 170992 252172 171048
rect 249701 170990 252172 170992
rect 288341 171048 290076 171050
rect 288341 170992 288346 171048
rect 288402 170992 290076 171048
rect 288341 170990 290076 170992
rect 315896 171048 315988 171050
rect 316052 171050 316058 171052
rect 315896 170992 315946 171048
rect 315896 170990 315988 170992
rect 249701 170987 249767 170990
rect 288341 170987 288407 170990
rect 315941 170988 315988 170990
rect 316052 170990 316134 171050
rect 316052 170988 316058 170990
rect 315941 170987 316007 170988
rect 304901 170914 304967 170917
rect 263948 170854 267750 170914
rect 301852 170912 304967 170914
rect 301852 170856 304906 170912
rect 304962 170856 304967 170912
rect 301852 170854 304967 170856
rect 266353 170506 266419 170509
rect 263948 170504 266419 170506
rect 263948 170448 266358 170504
rect 266414 170448 266419 170504
rect 263948 170446 266419 170448
rect 266353 170443 266419 170446
rect 249609 170370 249675 170373
rect 249609 170368 252172 170370
rect 249609 170312 249614 170368
rect 249670 170312 252172 170368
rect 249609 170310 252172 170312
rect 249609 170307 249675 170310
rect 267690 170234 267750 170854
rect 304901 170851 304967 170854
rect 301313 170642 301379 170645
rect 301270 170640 301379 170642
rect 301270 170584 301318 170640
rect 301374 170584 301379 170640
rect 301270 170579 301379 170584
rect 270033 170370 270099 170373
rect 277577 170370 277643 170373
rect 270033 170368 277643 170370
rect 270033 170312 270038 170368
rect 270094 170312 277582 170368
rect 277638 170312 277643 170368
rect 270033 170310 277643 170312
rect 270033 170307 270099 170310
rect 277577 170307 277643 170310
rect 276197 170234 276263 170237
rect 290046 170234 290106 170476
rect 267690 170232 276263 170234
rect 267690 170176 276202 170232
rect 276258 170176 276263 170232
rect 267690 170174 276263 170176
rect 276197 170171 276263 170174
rect 277350 170174 290106 170234
rect 301270 170204 301330 170579
rect 272701 170098 272767 170101
rect 277350 170098 277410 170174
rect 272701 170096 277410 170098
rect 272701 170040 272706 170096
rect 272762 170040 277410 170096
rect 272701 170038 277410 170040
rect 286409 170098 286475 170101
rect 286409 170096 290076 170098
rect 286409 170040 286414 170096
rect 286470 170040 290076 170096
rect 286409 170038 290076 170040
rect 272701 170035 272767 170038
rect 286409 170035 286475 170038
rect 266721 169962 266787 169965
rect 263948 169960 266787 169962
rect 263948 169904 266726 169960
rect 266782 169904 266787 169960
rect 263948 169902 266787 169904
rect 266721 169899 266787 169902
rect 166257 169690 166323 169693
rect 247769 169690 247835 169693
rect 166257 169688 247835 169690
rect 166257 169632 166262 169688
rect 166318 169632 247774 169688
rect 247830 169632 247835 169688
rect 166257 169630 247835 169632
rect 166257 169627 166323 169630
rect 247769 169627 247835 169630
rect 249701 169690 249767 169693
rect 288157 169690 288223 169693
rect 249701 169688 252172 169690
rect 249701 169632 249706 169688
rect 249762 169632 252172 169688
rect 249701 169630 252172 169632
rect 288157 169688 290076 169690
rect 288157 169632 288162 169688
rect 288218 169632 290076 169688
rect 288157 169630 290076 169632
rect 249701 169627 249767 169630
rect 288157 169627 288223 169630
rect 266353 169554 266419 169557
rect 263948 169552 266419 169554
rect 263948 169496 266358 169552
rect 266414 169496 266419 169552
rect 263948 169494 266419 169496
rect 266353 169491 266419 169494
rect 303889 169418 303955 169421
rect 301852 169416 303955 169418
rect 301852 169360 303894 169416
rect 303950 169360 303955 169416
rect 301852 169358 303955 169360
rect 303889 169355 303955 169358
rect 288249 169282 288315 169285
rect 288249 169280 290076 169282
rect 288249 169224 288254 169280
rect 288310 169224 290076 169280
rect 288249 169222 290076 169224
rect 288249 169219 288315 169222
rect 266997 169146 267063 169149
rect 269246 169146 269252 169148
rect 266997 169144 269252 169146
rect 266997 169088 267002 169144
rect 267058 169088 269252 169144
rect 266997 169086 269252 169088
rect 266997 169083 267063 169086
rect 269246 169084 269252 169086
rect 269316 169084 269322 169148
rect 249241 169010 249307 169013
rect 266353 169010 266419 169013
rect 249241 169008 252172 169010
rect 249241 168952 249246 169008
rect 249302 168952 252172 169008
rect 249241 168950 252172 168952
rect 263948 169008 266419 169010
rect 263948 168952 266358 169008
rect 266414 168952 266419 169008
rect 263948 168950 266419 168952
rect 249241 168947 249307 168950
rect 266353 168947 266419 168950
rect 272149 168602 272215 168605
rect 263948 168600 272215 168602
rect 263948 168544 272154 168600
rect 272210 168544 272215 168600
rect 263948 168542 272215 168544
rect 272149 168539 272215 168542
rect 284937 168602 285003 168605
rect 290046 168602 290106 168844
rect 302509 168738 302575 168741
rect 301852 168736 302575 168738
rect 301852 168680 302514 168736
rect 302570 168680 302575 168736
rect 301852 168678 302575 168680
rect 302509 168675 302575 168678
rect 284937 168600 290106 168602
rect 284937 168544 284942 168600
rect 284998 168544 290106 168600
rect 284937 168542 290106 168544
rect 284937 168539 285003 168542
rect 282177 168466 282243 168469
rect 282177 168464 290076 168466
rect 282177 168408 282182 168464
rect 282238 168408 290076 168464
rect 282177 168406 290076 168408
rect 282177 168403 282243 168406
rect 249701 168330 249767 168333
rect 249701 168328 252172 168330
rect 249701 168272 249706 168328
rect 249762 168272 252172 168328
rect 249701 168270 252172 168272
rect 249701 168267 249767 168270
rect 267641 168058 267707 168061
rect 263948 168056 267707 168058
rect 263948 168000 267646 168056
rect 267702 168000 267707 168056
rect 263948 167998 267707 168000
rect 267641 167995 267707 167998
rect 287973 167922 288039 167925
rect 305126 167922 305132 167924
rect 287973 167920 290076 167922
rect 287973 167864 287978 167920
rect 288034 167864 290076 167920
rect 287973 167862 290076 167864
rect 301852 167862 305132 167922
rect 287973 167859 288039 167862
rect 305126 167860 305132 167862
rect 305196 167860 305202 167924
rect 249609 167650 249675 167653
rect 266353 167650 266419 167653
rect 249609 167648 252172 167650
rect 249609 167592 249614 167648
rect 249670 167592 252172 167648
rect 249609 167590 252172 167592
rect 263948 167648 266419 167650
rect 263948 167592 266358 167648
rect 266414 167592 266419 167648
rect 263948 167590 266419 167592
rect 249609 167587 249675 167590
rect 266353 167587 266419 167590
rect 266721 167650 266787 167653
rect 281533 167650 281599 167653
rect 266721 167648 281599 167650
rect 266721 167592 266726 167648
rect 266782 167592 281538 167648
rect 281594 167592 281599 167648
rect 266721 167590 281599 167592
rect 266721 167587 266787 167590
rect 281533 167587 281599 167590
rect 289169 167514 289235 167517
rect 289169 167512 290076 167514
rect 289169 167456 289174 167512
rect 289230 167456 290076 167512
rect 289169 167454 290076 167456
rect 289169 167451 289235 167454
rect 278773 167378 278839 167381
rect 267690 167376 278839 167378
rect 267690 167320 278778 167376
rect 278834 167320 278839 167376
rect 267690 167318 278839 167320
rect 267690 167106 267750 167318
rect 278773 167315 278839 167318
rect 263948 167046 267750 167106
rect 288341 167106 288407 167109
rect 303889 167106 303955 167109
rect 288341 167104 290076 167106
rect 288341 167048 288346 167104
rect 288402 167048 290076 167104
rect 288341 167046 290076 167048
rect 301852 167104 303955 167106
rect 301852 167048 303894 167104
rect 303950 167048 303955 167104
rect 301852 167046 303955 167048
rect 288341 167043 288407 167046
rect 303889 167043 303955 167046
rect 248413 166970 248479 166973
rect 248413 166968 252172 166970
rect 248413 166912 248418 166968
rect 248474 166912 252172 166968
rect 248413 166910 252172 166912
rect 248413 166907 248479 166910
rect 267641 166698 267707 166701
rect 263948 166696 267707 166698
rect 263948 166640 267646 166696
rect 267702 166640 267707 166696
rect 263948 166638 267707 166640
rect 267641 166635 267707 166638
rect 288341 166698 288407 166701
rect 288341 166696 290076 166698
rect 288341 166640 288346 166696
rect 288402 166640 290076 166696
rect 288341 166638 290076 166640
rect 288341 166635 288407 166638
rect 270350 166500 270356 166564
rect 270420 166562 270426 166564
rect 277485 166562 277551 166565
rect 270420 166560 277551 166562
rect 270420 166504 277490 166560
rect 277546 166504 277551 166560
rect 270420 166502 277551 166504
rect 270420 166500 270426 166502
rect 277485 166499 277551 166502
rect 248505 166426 248571 166429
rect 276841 166426 276907 166429
rect 288249 166426 288315 166429
rect 303889 166426 303955 166429
rect 248505 166424 252172 166426
rect 248505 166368 248510 166424
rect 248566 166368 252172 166424
rect 248505 166366 252172 166368
rect 276841 166424 288315 166426
rect 276841 166368 276846 166424
rect 276902 166368 288254 166424
rect 288310 166368 288315 166424
rect 276841 166366 288315 166368
rect 301852 166424 303955 166426
rect 301852 166368 303894 166424
rect 303950 166368 303955 166424
rect 301852 166366 303955 166368
rect 248505 166363 248571 166366
rect 276841 166363 276907 166366
rect 288249 166363 288315 166366
rect 303889 166363 303955 166366
rect 268326 166228 268332 166292
rect 268396 166290 268402 166292
rect 282913 166290 282979 166293
rect 268396 166288 282979 166290
rect 268396 166232 282918 166288
rect 282974 166232 282979 166288
rect 268396 166230 282979 166232
rect 268396 166228 268402 166230
rect 282913 166227 282979 166230
rect 288249 166290 288315 166293
rect 288249 166288 290076 166290
rect 288249 166232 288254 166288
rect 288310 166232 290076 166288
rect 288249 166230 290076 166232
rect 288249 166227 288315 166230
rect 266353 166154 266419 166157
rect 263948 166152 266419 166154
rect 263948 166096 266358 166152
rect 266414 166096 266419 166152
rect 263948 166094 266419 166096
rect 266353 166091 266419 166094
rect 238109 166018 238175 166021
rect 238109 166016 252202 166018
rect 238109 165960 238114 166016
rect 238170 165960 252202 166016
rect 238109 165958 252202 165960
rect 238109 165955 238175 165958
rect 252142 165716 252202 165958
rect 288065 165882 288131 165885
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 288065 165880 290076 165882
rect 288065 165824 288070 165880
rect 288126 165824 290076 165880
rect 288065 165822 290076 165824
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 288065 165819 288131 165822
rect 580165 165819 580231 165822
rect 270677 165746 270743 165749
rect 263948 165744 270743 165746
rect 263948 165688 270682 165744
rect 270738 165688 270743 165744
rect 583520 165732 584960 165822
rect 263948 165686 270743 165688
rect 270677 165683 270743 165686
rect 265014 165548 265020 165612
rect 265084 165610 265090 165612
rect 265341 165610 265407 165613
rect 265084 165608 265407 165610
rect 265084 165552 265346 165608
rect 265402 165552 265407 165608
rect 265084 165550 265407 165552
rect 265084 165548 265090 165550
rect 265341 165547 265407 165550
rect 271965 165610 272031 165613
rect 272558 165610 272564 165612
rect 271965 165608 272564 165610
rect 271965 165552 271970 165608
rect 272026 165552 272564 165608
rect 271965 165550 272564 165552
rect 271965 165547 272031 165550
rect 272558 165548 272564 165550
rect 272628 165548 272634 165612
rect 266353 165202 266419 165205
rect 263948 165200 266419 165202
rect 263948 165144 266358 165200
rect 266414 165144 266419 165200
rect 263948 165142 266419 165144
rect 266353 165139 266419 165142
rect 248413 165066 248479 165069
rect 290046 165066 290106 165308
rect 248413 165064 252172 165066
rect 248413 165008 248418 165064
rect 248474 165008 252172 165064
rect 248413 165006 252172 165008
rect 288574 165006 290106 165066
rect 301822 165066 301882 165580
rect 301822 165006 306390 165066
rect 248413 165003 248479 165006
rect 265566 164868 265572 164932
rect 265636 164930 265642 164932
rect 287789 164930 287855 164933
rect 265636 164928 287855 164930
rect 265636 164872 287794 164928
rect 287850 164872 287855 164928
rect 265636 164870 287855 164872
rect 265636 164868 265642 164870
rect 287789 164867 287855 164870
rect 265157 164794 265223 164797
rect 263948 164792 265223 164794
rect 263948 164736 265162 164792
rect 265218 164736 265223 164792
rect 263948 164734 265223 164736
rect 265157 164731 265223 164734
rect 273989 164658 274055 164661
rect 288574 164658 288634 165006
rect 303889 164930 303955 164933
rect 301852 164928 303955 164930
rect 273989 164656 288634 164658
rect 273989 164600 273994 164656
rect 274050 164600 288634 164656
rect 273989 164598 288634 164600
rect 288709 164658 288775 164661
rect 290046 164658 290106 164900
rect 301852 164872 303894 164928
rect 303950 164872 303955 164928
rect 301852 164870 303955 164872
rect 303889 164867 303955 164870
rect 288709 164656 290106 164658
rect 288709 164600 288714 164656
rect 288770 164600 290106 164656
rect 288709 164598 290106 164600
rect 273989 164595 274055 164598
rect 288709 164595 288775 164598
rect 264053 164522 264119 164525
rect 287421 164522 287487 164525
rect 264053 164520 264162 164522
rect 264053 164464 264058 164520
rect 264114 164464 264162 164520
rect 264053 164459 264162 164464
rect 287421 164520 290076 164522
rect 287421 164464 287426 164520
rect 287482 164464 290076 164520
rect 287421 164462 290076 164464
rect 287421 164459 287487 164462
rect 164734 164324 164740 164388
rect 164804 164386 164810 164388
rect 264102 164386 264162 164459
rect 164804 164326 238770 164386
rect 164804 164324 164810 164326
rect 238710 164250 238770 164326
rect 244230 164326 252172 164386
rect 263948 164326 264162 164386
rect 306330 164386 306390 165006
rect 306598 164386 306604 164388
rect 306330 164326 306604 164386
rect 244230 164250 244290 164326
rect 306598 164324 306604 164326
rect 306668 164324 306674 164388
rect 273437 164252 273503 164253
rect 273437 164250 273484 164252
rect 238710 164190 244290 164250
rect 273392 164248 273484 164250
rect 273392 164192 273442 164248
rect 273392 164190 273484 164192
rect 273437 164188 273484 164190
rect 273548 164188 273554 164252
rect 273437 164187 273503 164188
rect 288157 164114 288223 164117
rect 303889 164114 303955 164117
rect 288157 164112 290076 164114
rect 288157 164056 288162 164112
rect 288218 164056 290076 164112
rect 288157 164054 290076 164056
rect 301852 164112 303955 164114
rect 301852 164056 303894 164112
rect 303950 164056 303955 164112
rect 301852 164054 303955 164056
rect 288157 164051 288223 164054
rect 303889 164051 303955 164054
rect 269062 163842 269068 163844
rect 263948 163782 269068 163842
rect 269062 163780 269068 163782
rect 269132 163780 269138 163844
rect 248413 163706 248479 163709
rect 287881 163706 287947 163709
rect 248413 163704 252172 163706
rect 248413 163648 248418 163704
rect 248474 163648 252172 163704
rect 248413 163646 252172 163648
rect 287881 163704 290076 163706
rect 287881 163648 287886 163704
rect 287942 163648 290076 163704
rect 287881 163646 290076 163648
rect 248413 163643 248479 163646
rect 287881 163643 287947 163646
rect 266353 163434 266419 163437
rect 263948 163432 266419 163434
rect 263948 163376 266358 163432
rect 266414 163376 266419 163432
rect 263948 163374 266419 163376
rect 266353 163371 266419 163374
rect 269614 163372 269620 163436
rect 269684 163434 269690 163436
rect 287421 163434 287487 163437
rect 269684 163432 287487 163434
rect 269684 163376 287426 163432
rect 287482 163376 287487 163432
rect 269684 163374 287487 163376
rect 269684 163372 269690 163374
rect 287421 163371 287487 163374
rect 288249 163298 288315 163301
rect 303889 163298 303955 163301
rect 288249 163296 290076 163298
rect 288249 163240 288254 163296
rect 288310 163240 290076 163296
rect 288249 163238 290076 163240
rect 301852 163296 303955 163298
rect 301852 163240 303894 163296
rect 303950 163240 303955 163296
rect 301852 163238 303955 163240
rect 288249 163235 288315 163238
rect 303889 163235 303955 163238
rect 248505 163026 248571 163029
rect 248505 163024 252172 163026
rect -960 162890 480 162980
rect 248505 162968 248510 163024
rect 248566 162968 252172 163024
rect 248505 162966 252172 162968
rect 248505 162963 248571 162966
rect 3233 162890 3299 162893
rect 266721 162890 266787 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect 263948 162888 266787 162890
rect 263948 162832 266726 162888
rect 266782 162832 266787 162888
rect 263948 162830 266787 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 266721 162827 266787 162830
rect 286317 162890 286383 162893
rect 286317 162888 290076 162890
rect 286317 162832 286322 162888
rect 286378 162832 290076 162888
rect 286317 162830 290076 162832
rect 286317 162827 286383 162830
rect 270585 162754 270651 162757
rect 270718 162754 270724 162756
rect 270585 162752 270724 162754
rect 270585 162696 270590 162752
rect 270646 162696 270724 162752
rect 270585 162694 270724 162696
rect 270585 162691 270651 162694
rect 270718 162692 270724 162694
rect 270788 162692 270794 162756
rect 283782 162692 283788 162756
rect 283852 162754 283858 162756
rect 285673 162754 285739 162757
rect 283852 162752 285739 162754
rect 283852 162696 285678 162752
rect 285734 162696 285739 162752
rect 283852 162694 285739 162696
rect 283852 162692 283858 162694
rect 285673 162691 285739 162694
rect 303889 162618 303955 162621
rect 301852 162616 303955 162618
rect 301852 162560 303894 162616
rect 303950 162560 303955 162616
rect 301852 162558 303955 162560
rect 303889 162555 303955 162558
rect 276238 162482 276244 162484
rect 263948 162422 276244 162482
rect 276238 162420 276244 162422
rect 276308 162420 276314 162484
rect 248413 162346 248479 162349
rect 288341 162346 288407 162349
rect 248413 162344 252172 162346
rect 248413 162288 248418 162344
rect 248474 162288 252172 162344
rect 248413 162286 252172 162288
rect 288341 162344 290076 162346
rect 288341 162288 288346 162344
rect 288402 162288 290076 162344
rect 288341 162286 290076 162288
rect 248413 162283 248479 162286
rect 288341 162283 288407 162286
rect 275277 162074 275343 162077
rect 288065 162074 288131 162077
rect 275277 162072 288131 162074
rect 275277 162016 275282 162072
rect 275338 162016 288070 162072
rect 288126 162016 288131 162072
rect 275277 162014 288131 162016
rect 275277 162011 275343 162014
rect 288065 162011 288131 162014
rect 266353 161938 266419 161941
rect 263948 161936 266419 161938
rect 263948 161880 266358 161936
rect 266414 161880 266419 161936
rect 263948 161878 266419 161880
rect 266353 161875 266419 161878
rect 287145 161938 287211 161941
rect 287145 161936 290076 161938
rect 287145 161880 287150 161936
rect 287206 161880 290076 161936
rect 287145 161878 290076 161880
rect 287145 161875 287211 161878
rect 248505 161802 248571 161805
rect 302325 161802 302391 161805
rect 248505 161800 252172 161802
rect 248505 161744 248510 161800
rect 248566 161744 252172 161800
rect 248505 161742 252172 161744
rect 301852 161800 302391 161802
rect 301852 161744 302330 161800
rect 302386 161744 302391 161800
rect 301852 161742 302391 161744
rect 248505 161739 248571 161742
rect 302325 161739 302391 161742
rect 315982 161604 315988 161668
rect 316052 161604 316058 161668
rect 315990 161533 316050 161604
rect 266537 161530 266603 161533
rect 263948 161528 266603 161530
rect 263948 161472 266542 161528
rect 266598 161472 266603 161528
rect 263948 161470 266603 161472
rect 266537 161467 266603 161470
rect 274030 161468 274036 161532
rect 274100 161530 274106 161532
rect 315941 161530 316050 161533
rect 274100 161470 290076 161530
rect 315896 161528 316050 161530
rect 315896 161472 315946 161528
rect 316002 161472 316050 161528
rect 315896 161470 316050 161472
rect 274100 161468 274106 161470
rect 315941 161467 316007 161470
rect 315941 161394 316007 161397
rect 315896 161392 316050 161394
rect 315896 161336 315946 161392
rect 316002 161336 316050 161392
rect 315896 161334 316050 161336
rect 315941 161331 316050 161334
rect 315990 161260 316050 161331
rect 315982 161196 315988 161260
rect 316052 161196 316058 161260
rect 248413 161122 248479 161125
rect 287513 161122 287579 161125
rect 303889 161122 303955 161125
rect 248413 161120 252172 161122
rect 248413 161064 248418 161120
rect 248474 161064 252172 161120
rect 248413 161062 252172 161064
rect 287513 161120 290076 161122
rect 287513 161064 287518 161120
rect 287574 161064 290076 161120
rect 287513 161062 290076 161064
rect 301852 161120 303955 161122
rect 301852 161064 303894 161120
rect 303950 161064 303955 161120
rect 301852 161062 303955 161064
rect 248413 161059 248479 161062
rect 287513 161059 287579 161062
rect 303889 161059 303955 161062
rect 266353 160986 266419 160989
rect 263948 160984 266419 160986
rect 263948 160928 266358 160984
rect 266414 160928 266419 160984
rect 263948 160926 266419 160928
rect 266353 160923 266419 160926
rect 301313 160850 301379 160853
rect 301270 160848 301379 160850
rect 301270 160792 301318 160848
rect 301374 160792 301379 160848
rect 301270 160787 301379 160792
rect 175917 160714 175983 160717
rect 240133 160714 240199 160717
rect 175917 160712 240199 160714
rect 175917 160656 175922 160712
rect 175978 160656 240138 160712
rect 240194 160656 240199 160712
rect 175917 160654 240199 160656
rect 175917 160651 175983 160654
rect 240133 160651 240199 160654
rect 267733 160714 267799 160717
rect 284293 160714 284359 160717
rect 267733 160712 284359 160714
rect 267733 160656 267738 160712
rect 267794 160656 284298 160712
rect 284354 160656 284359 160712
rect 267733 160654 284359 160656
rect 267733 160651 267799 160654
rect 284293 160651 284359 160654
rect 265065 160578 265131 160581
rect 263948 160576 265131 160578
rect 263948 160520 265070 160576
rect 265126 160520 265131 160576
rect 263948 160518 265131 160520
rect 265065 160515 265131 160518
rect 248505 160442 248571 160445
rect 278037 160442 278103 160445
rect 290046 160442 290106 160684
rect 248505 160440 252172 160442
rect 248505 160384 248510 160440
rect 248566 160384 252172 160440
rect 248505 160382 252172 160384
rect 278037 160440 290106 160442
rect 278037 160384 278042 160440
rect 278098 160384 290106 160440
rect 278037 160382 290106 160384
rect 248505 160379 248571 160382
rect 278037 160379 278103 160382
rect 286501 160306 286567 160309
rect 286501 160304 290076 160306
rect 286501 160248 286506 160304
rect 286562 160248 290076 160304
rect 301270 160276 301330 160787
rect 286501 160246 290076 160248
rect 286501 160243 286567 160246
rect 266537 160170 266603 160173
rect 267774 160170 267780 160172
rect 266537 160168 267780 160170
rect 266537 160112 266542 160168
rect 266598 160112 267780 160168
rect 266537 160110 267780 160112
rect 266537 160107 266603 160110
rect 267774 160108 267780 160110
rect 267844 160108 267850 160172
rect 266445 160034 266511 160037
rect 263948 160032 266511 160034
rect 263948 159976 266450 160032
rect 266506 159976 266511 160032
rect 263948 159974 266511 159976
rect 266445 159971 266511 159974
rect 249149 159762 249215 159765
rect 288341 159762 288407 159765
rect 249149 159760 252172 159762
rect 249149 159704 249154 159760
rect 249210 159704 252172 159760
rect 249149 159702 252172 159704
rect 288341 159760 290076 159762
rect 288341 159704 288346 159760
rect 288402 159704 290076 159760
rect 288341 159702 290076 159704
rect 249149 159699 249215 159702
rect 288341 159699 288407 159702
rect 267641 159626 267707 159629
rect 263948 159624 267707 159626
rect 263948 159568 267646 159624
rect 267702 159568 267707 159624
rect 263948 159566 267707 159568
rect 267641 159563 267707 159566
rect 302417 159490 302483 159493
rect 301852 159488 302483 159490
rect 301852 159432 302422 159488
rect 302478 159432 302483 159488
rect 301852 159430 302483 159432
rect 302417 159427 302483 159430
rect 266813 159354 266879 159357
rect 274725 159354 274791 159357
rect 266813 159352 274791 159354
rect 266813 159296 266818 159352
rect 266874 159296 274730 159352
rect 274786 159296 274791 159352
rect 266813 159294 274791 159296
rect 266813 159291 266879 159294
rect 274725 159291 274791 159294
rect 248413 159082 248479 159085
rect 266302 159082 266308 159084
rect 248413 159080 252172 159082
rect 248413 159024 248418 159080
rect 248474 159024 252172 159080
rect 248413 159022 252172 159024
rect 263948 159022 266308 159082
rect 248413 159019 248479 159022
rect 266302 159020 266308 159022
rect 266372 159020 266378 159084
rect 268377 159082 268443 159085
rect 290046 159082 290106 159324
rect 268377 159080 290106 159082
rect 268377 159024 268382 159080
rect 268438 159024 290106 159080
rect 268377 159022 290106 159024
rect 268377 159019 268443 159022
rect 287421 158946 287487 158949
rect 287421 158944 290076 158946
rect 287421 158888 287426 158944
rect 287482 158888 290076 158944
rect 287421 158886 290076 158888
rect 287421 158883 287487 158886
rect 303797 158810 303863 158813
rect 301852 158808 303863 158810
rect 301852 158752 303802 158808
rect 303858 158752 303863 158808
rect 301852 158750 303863 158752
rect 303797 158747 303863 158750
rect 263948 158614 267750 158674
rect 267690 158538 267750 158614
rect 269205 158538 269271 158541
rect 267690 158536 269271 158538
rect 267690 158480 269210 158536
rect 269266 158480 269271 158536
rect 267690 158478 269271 158480
rect 269205 158475 269271 158478
rect 288249 158538 288315 158541
rect 288249 158536 290076 158538
rect 288249 158480 288254 158536
rect 288310 158480 290076 158536
rect 288249 158478 290076 158480
rect 288249 158475 288315 158478
rect 248413 158402 248479 158405
rect 248413 158400 252172 158402
rect 248413 158344 248418 158400
rect 248474 158344 252172 158400
rect 248413 158342 252172 158344
rect 248413 158339 248479 158342
rect 266353 158130 266419 158133
rect 263948 158128 266419 158130
rect 263948 158072 266358 158128
rect 266414 158072 266419 158128
rect 263948 158070 266419 158072
rect 266353 158067 266419 158070
rect 288341 158130 288407 158133
rect 288341 158128 290076 158130
rect 288341 158072 288346 158128
rect 288402 158072 290076 158128
rect 288341 158070 290076 158072
rect 288341 158067 288407 158070
rect 275553 157994 275619 157997
rect 283005 157994 283071 157997
rect 303613 157994 303679 157997
rect 275553 157992 283071 157994
rect 275553 157936 275558 157992
rect 275614 157936 283010 157992
rect 283066 157936 283071 157992
rect 275553 157934 283071 157936
rect 301852 157992 303679 157994
rect 301852 157936 303618 157992
rect 303674 157936 303679 157992
rect 301852 157934 303679 157936
rect 275553 157931 275619 157934
rect 283005 157931 283071 157934
rect 303613 157931 303679 157934
rect 249057 157722 249123 157725
rect 266629 157722 266695 157725
rect 249057 157720 252172 157722
rect 249057 157664 249062 157720
rect 249118 157664 252172 157720
rect 249057 157662 252172 157664
rect 263948 157720 266695 157722
rect 263948 157664 266634 157720
rect 266690 157664 266695 157720
rect 263948 157662 266695 157664
rect 249057 157659 249123 157662
rect 266629 157659 266695 157662
rect 277350 157662 290076 157722
rect 272517 157586 272583 157589
rect 277350 157586 277410 157662
rect 272517 157584 277410 157586
rect 272517 157528 272522 157584
rect 272578 157528 277410 157584
rect 272517 157526 277410 157528
rect 272517 157523 272583 157526
rect 269113 157450 269179 157453
rect 278773 157452 278839 157453
rect 270350 157450 270356 157452
rect 269113 157448 270356 157450
rect 269113 157392 269118 157448
rect 269174 157392 270356 157448
rect 269113 157390 270356 157392
rect 269113 157387 269179 157390
rect 270350 157388 270356 157390
rect 270420 157388 270426 157452
rect 278773 157450 278820 157452
rect 278728 157448 278820 157450
rect 278728 157392 278778 157448
rect 278728 157390 278820 157392
rect 278773 157388 278820 157390
rect 278884 157388 278890 157452
rect 287697 157450 287763 157453
rect 288382 157450 288388 157452
rect 287697 157448 288388 157450
rect 287697 157392 287702 157448
rect 287758 157392 288388 157448
rect 287697 157390 288388 157392
rect 278773 157387 278839 157388
rect 287697 157387 287763 157390
rect 288382 157388 288388 157390
rect 288452 157388 288458 157452
rect 303797 157314 303863 157317
rect 301852 157312 303863 157314
rect 301852 157256 303802 157312
rect 303858 157256 303863 157312
rect 301852 157254 303863 157256
rect 303797 157251 303863 157254
rect 249701 157178 249767 157181
rect 266353 157178 266419 157181
rect 249701 157176 252172 157178
rect 249701 157120 249706 157176
rect 249762 157120 252172 157176
rect 249701 157118 252172 157120
rect 263948 157176 266419 157178
rect 263948 157120 266358 157176
rect 266414 157120 266419 157176
rect 263948 157118 266419 157120
rect 249701 157115 249767 157118
rect 266353 157115 266419 157118
rect 288157 157178 288223 157181
rect 288157 157176 290076 157178
rect 288157 157120 288162 157176
rect 288218 157120 290076 157176
rect 288157 157118 290076 157120
rect 288157 157115 288223 157118
rect 266537 156906 266603 156909
rect 265390 156904 266603 156906
rect 265390 156848 266542 156904
rect 266598 156848 266603 156904
rect 265390 156846 266603 156848
rect 265390 156770 265450 156846
rect 266537 156843 266603 156846
rect 268510 156844 268516 156908
rect 268580 156906 268586 156908
rect 278865 156906 278931 156909
rect 268580 156904 278931 156906
rect 268580 156848 278870 156904
rect 278926 156848 278931 156904
rect 268580 156846 278931 156848
rect 268580 156844 268586 156846
rect 278865 156843 278931 156846
rect 263948 156710 265450 156770
rect 266445 156770 266511 156773
rect 285765 156770 285831 156773
rect 266445 156768 285831 156770
rect 266445 156712 266450 156768
rect 266506 156712 285770 156768
rect 285826 156712 285831 156768
rect 266445 156710 285831 156712
rect 266445 156707 266511 156710
rect 285765 156707 285831 156710
rect 288065 156770 288131 156773
rect 288065 156768 290076 156770
rect 288065 156712 288070 156768
rect 288126 156712 290076 156768
rect 288065 156710 290076 156712
rect 288065 156707 288131 156710
rect 267038 156572 267044 156636
rect 267108 156634 267114 156636
rect 288433 156634 288499 156637
rect 267108 156632 288499 156634
rect 267108 156576 288438 156632
rect 288494 156576 288499 156632
rect 267108 156574 288499 156576
rect 267108 156572 267114 156574
rect 288433 156571 288499 156574
rect 249609 156498 249675 156501
rect 303889 156498 303955 156501
rect 249609 156496 252172 156498
rect 249609 156440 249614 156496
rect 249670 156440 252172 156496
rect 249609 156438 252172 156440
rect 301852 156496 303955 156498
rect 301852 156440 303894 156496
rect 303950 156440 303955 156496
rect 301852 156438 303955 156440
rect 249609 156435 249675 156438
rect 303889 156435 303955 156438
rect 287010 156302 290076 156362
rect 266854 156226 266860 156228
rect 263948 156166 266860 156226
rect 266854 156164 266860 156166
rect 266924 156164 266930 156228
rect 273437 155956 273503 155957
rect 273437 155954 273484 155956
rect 273392 155952 273484 155954
rect 273392 155896 273442 155952
rect 273392 155894 273484 155896
rect 273437 155892 273484 155894
rect 273548 155892 273554 155956
rect 285029 155954 285095 155957
rect 287010 155954 287070 156302
rect 285029 155952 287070 155954
rect 285029 155896 285034 155952
rect 285090 155896 287070 155952
rect 285029 155894 287070 155896
rect 287973 155954 288039 155957
rect 287973 155952 290076 155954
rect 287973 155896 287978 155952
rect 288034 155896 290076 155952
rect 287973 155894 290076 155896
rect 273437 155891 273503 155892
rect 285029 155891 285095 155894
rect 287973 155891 288039 155894
rect 249701 155818 249767 155821
rect 266353 155818 266419 155821
rect 249701 155816 252172 155818
rect 249701 155760 249706 155816
rect 249762 155760 252172 155816
rect 249701 155758 252172 155760
rect 263948 155816 266419 155818
rect 263948 155760 266358 155816
rect 266414 155760 266419 155816
rect 263948 155758 266419 155760
rect 249701 155755 249767 155758
rect 266353 155755 266419 155758
rect 303797 155682 303863 155685
rect 301852 155680 303863 155682
rect 301852 155624 303802 155680
rect 303858 155624 303863 155680
rect 301852 155622 303863 155624
rect 303797 155619 303863 155622
rect 266445 155274 266511 155277
rect 263948 155272 266511 155274
rect 263948 155216 266450 155272
rect 266506 155216 266511 155272
rect 263948 155214 266511 155216
rect 266445 155211 266511 155214
rect 271137 155274 271203 155277
rect 288065 155274 288131 155277
rect 290046 155274 290106 155516
rect 271137 155272 288131 155274
rect 271137 155216 271142 155272
rect 271198 155216 288070 155272
rect 288126 155216 288131 155272
rect 271137 155214 288131 155216
rect 271137 155211 271203 155214
rect 288065 155211 288131 155214
rect 288206 155214 290106 155274
rect 249609 155138 249675 155141
rect 249609 155136 252172 155138
rect 249609 155080 249614 155136
rect 249670 155080 252172 155136
rect 249609 155078 252172 155080
rect 249609 155075 249675 155078
rect 273294 154866 273300 154868
rect 263948 154806 273300 154866
rect 273294 154804 273300 154806
rect 273364 154804 273370 154868
rect 286593 154866 286659 154869
rect 288206 154866 288266 155214
rect 288341 155138 288407 155141
rect 288341 155136 290076 155138
rect 288341 155080 288346 155136
rect 288402 155080 290076 155136
rect 288341 155078 290076 155080
rect 288341 155075 288407 155078
rect 303613 155002 303679 155005
rect 301852 155000 303679 155002
rect 301852 154944 303618 155000
rect 303674 154944 303679 155000
rect 301852 154942 303679 154944
rect 303613 154939 303679 154942
rect 286593 154864 288266 154866
rect 286593 154808 286598 154864
rect 286654 154808 288266 154864
rect 286593 154806 288266 154808
rect 286593 154803 286659 154806
rect 287789 154594 287855 154597
rect 287789 154592 290076 154594
rect 287789 154536 287794 154592
rect 287850 154536 290076 154592
rect 287789 154534 290076 154536
rect 287789 154531 287855 154534
rect 249149 154458 249215 154461
rect 265065 154460 265131 154461
rect 265014 154458 265020 154460
rect 249149 154456 252172 154458
rect 249149 154400 249154 154456
rect 249210 154400 252172 154456
rect 249149 154398 252172 154400
rect 264974 154398 265020 154458
rect 265084 154456 265131 154460
rect 265126 154400 265131 154456
rect 249149 154395 249215 154398
rect 265014 154396 265020 154398
rect 265084 154396 265131 154400
rect 265065 154395 265131 154396
rect 265750 154322 265756 154324
rect 263948 154262 265756 154322
rect 265750 154260 265756 154262
rect 265820 154260 265826 154324
rect 303613 154186 303679 154189
rect 301852 154184 303679 154186
rect 266353 153914 266419 153917
rect 263948 153912 266419 153914
rect 263948 153856 266358 153912
rect 266414 153856 266419 153912
rect 263948 153854 266419 153856
rect 266353 153851 266419 153854
rect 278221 153914 278287 153917
rect 290046 153914 290106 154156
rect 301852 154128 303618 154184
rect 303674 154128 303679 154184
rect 301852 154126 303679 154128
rect 303613 154123 303679 154126
rect 278221 153912 290106 153914
rect 278221 153856 278226 153912
rect 278282 153856 290106 153912
rect 278221 153854 290106 153856
rect 278221 153851 278287 153854
rect 249701 153778 249767 153781
rect 264881 153778 264947 153781
rect 280102 153778 280108 153780
rect 249701 153776 252172 153778
rect 249701 153720 249706 153776
rect 249762 153720 252172 153776
rect 249701 153718 252172 153720
rect 264881 153776 280108 153778
rect 264881 153720 264886 153776
rect 264942 153720 280108 153776
rect 264881 153718 280108 153720
rect 249701 153715 249767 153718
rect 264881 153715 264947 153718
rect 280102 153716 280108 153718
rect 280172 153716 280178 153780
rect 289077 153778 289143 153781
rect 289077 153776 290076 153778
rect 289077 153720 289082 153776
rect 289138 153720 290076 153776
rect 289077 153718 290076 153720
rect 289077 153715 289143 153718
rect 303797 153506 303863 153509
rect 301852 153504 303863 153506
rect 301852 153448 303802 153504
rect 303858 153448 303863 153504
rect 301852 153446 303863 153448
rect 303797 153443 303863 153446
rect 266353 153370 266419 153373
rect 263948 153368 266419 153370
rect 263948 153312 266358 153368
rect 266414 153312 266419 153368
rect 263948 153310 266419 153312
rect 266353 153307 266419 153310
rect 280654 153308 280660 153372
rect 280724 153370 280730 153372
rect 280724 153310 290076 153370
rect 280724 153308 280730 153310
rect 248965 153098 249031 153101
rect 248965 153096 252172 153098
rect 248965 153040 248970 153096
rect 249026 153040 252172 153096
rect 248965 153038 252172 153040
rect 248965 153035 249031 153038
rect 266721 152962 266787 152965
rect 263948 152960 266787 152962
rect 263948 152904 266726 152960
rect 266782 152904 266787 152960
rect 263948 152902 266787 152904
rect 266721 152899 266787 152902
rect 290046 152690 290106 152932
rect 303797 152690 303863 152693
rect 287010 152630 290106 152690
rect 301852 152688 303863 152690
rect 301852 152632 303802 152688
rect 303858 152632 303863 152688
rect 301852 152630 303863 152632
rect 249333 152554 249399 152557
rect 265341 152554 265407 152557
rect 249333 152552 252172 152554
rect 249333 152496 249338 152552
rect 249394 152496 252172 152552
rect 249333 152494 252172 152496
rect 263948 152552 265407 152554
rect 263948 152496 265346 152552
rect 265402 152496 265407 152552
rect 263948 152494 265407 152496
rect 249333 152491 249399 152494
rect 265341 152491 265407 152494
rect 266721 152418 266787 152421
rect 278129 152418 278195 152421
rect 266721 152416 278195 152418
rect 266721 152360 266726 152416
rect 266782 152360 278134 152416
rect 278190 152360 278195 152416
rect 266721 152358 278195 152360
rect 266721 152355 266787 152358
rect 278129 152355 278195 152358
rect 276790 152084 276796 152148
rect 276860 152146 276866 152148
rect 287010 152146 287070 152630
rect 303797 152627 303863 152630
rect 583385 152690 583451 152693
rect 583520 152690 584960 152780
rect 583385 152688 584960 152690
rect 583385 152632 583390 152688
rect 583446 152632 584960 152688
rect 583385 152630 584960 152632
rect 583385 152627 583451 152630
rect 288249 152554 288315 152557
rect 288249 152552 290076 152554
rect 288249 152496 288254 152552
rect 288310 152496 290076 152552
rect 583520 152540 584960 152630
rect 288249 152494 290076 152496
rect 288249 152491 288315 152494
rect 276860 152086 287070 152146
rect 276860 152084 276866 152086
rect 266813 152010 266879 152013
rect 263948 152008 266879 152010
rect 263948 151952 266818 152008
rect 266874 151952 266879 152008
rect 263948 151950 266879 151952
rect 266813 151947 266879 151950
rect 288341 152010 288407 152013
rect 288341 152008 290076 152010
rect 288341 151952 288346 152008
rect 288402 151952 290076 152008
rect 288341 151950 290076 151952
rect 288341 151947 288407 151950
rect 249701 151874 249767 151877
rect 303889 151874 303955 151877
rect 315941 151876 316007 151877
rect 315941 151874 315988 151876
rect 249701 151872 252172 151874
rect 249701 151816 249706 151872
rect 249762 151816 252172 151872
rect 249701 151814 252172 151816
rect 301852 151872 303955 151874
rect 301852 151816 303894 151872
rect 303950 151816 303955 151872
rect 301852 151814 303955 151816
rect 315896 151872 315988 151874
rect 316052 151874 316058 151876
rect 315896 151816 315946 151872
rect 315896 151814 315988 151816
rect 249701 151811 249767 151814
rect 303889 151811 303955 151814
rect 315941 151812 315988 151814
rect 316052 151814 316134 151874
rect 316052 151812 316058 151814
rect 315941 151811 316007 151812
rect 315941 151738 316007 151741
rect 315896 151736 316050 151738
rect 315896 151680 315946 151736
rect 316002 151680 316050 151736
rect 315896 151678 316050 151680
rect 315941 151675 316050 151678
rect 266353 151602 266419 151605
rect 263948 151600 266419 151602
rect 263948 151544 266358 151600
rect 266414 151544 266419 151600
rect 263948 151542 266419 151544
rect 266353 151539 266419 151542
rect 288341 151602 288407 151605
rect 315990 151604 316050 151675
rect 288341 151600 290076 151602
rect 288341 151544 288346 151600
rect 288402 151544 290076 151600
rect 288341 151542 290076 151544
rect 288341 151539 288407 151542
rect 315982 151540 315988 151604
rect 316052 151540 316058 151604
rect 266445 151330 266511 151333
rect 268326 151330 268332 151332
rect 266445 151328 268332 151330
rect 266445 151272 266450 151328
rect 266506 151272 268332 151328
rect 266445 151270 268332 151272
rect 266445 151267 266511 151270
rect 268326 151268 268332 151270
rect 268396 151268 268402 151332
rect 249241 151194 249307 151197
rect 249241 151192 252172 151194
rect 249241 151136 249246 151192
rect 249302 151136 252172 151192
rect 249241 151134 252172 151136
rect 249241 151131 249307 151134
rect 266854 151132 266860 151196
rect 266924 151194 266930 151196
rect 276749 151194 276815 151197
rect 266924 151192 276815 151194
rect 266924 151136 276754 151192
rect 276810 151136 276815 151192
rect 266924 151134 276815 151136
rect 266924 151132 266930 151134
rect 276749 151131 276815 151134
rect 287973 151194 288039 151197
rect 303705 151194 303771 151197
rect 287973 151192 290076 151194
rect 287973 151136 287978 151192
rect 288034 151136 290076 151192
rect 287973 151134 290076 151136
rect 301852 151192 303771 151194
rect 301852 151136 303710 151192
rect 303766 151136 303771 151192
rect 301852 151134 303771 151136
rect 287973 151131 288039 151134
rect 303705 151131 303771 151134
rect 264094 151058 264100 151060
rect 263948 150998 264100 151058
rect 264094 150996 264100 150998
rect 264164 150996 264170 151060
rect 269798 150996 269804 151060
rect 269868 151058 269874 151060
rect 285806 151058 285812 151060
rect 269868 150998 285812 151058
rect 269868 150996 269874 150998
rect 285806 150996 285812 150998
rect 285876 150996 285882 151060
rect 288249 150786 288315 150789
rect 288249 150784 290076 150786
rect 288249 150728 288254 150784
rect 288310 150728 290076 150784
rect 288249 150726 290076 150728
rect 288249 150723 288315 150726
rect 301313 150650 301379 150653
rect 263948 150590 267750 150650
rect 249701 150514 249767 150517
rect 249701 150512 252172 150514
rect 249701 150456 249706 150512
rect 249762 150456 252172 150512
rect 249701 150454 252172 150456
rect 249701 150451 249767 150454
rect 264094 150452 264100 150516
rect 264164 150514 264170 150516
rect 264881 150514 264947 150517
rect 264164 150512 264947 150514
rect 264164 150456 264886 150512
rect 264942 150456 264947 150512
rect 264164 150454 264947 150456
rect 267690 150514 267750 150590
rect 301270 150648 301379 150650
rect 301270 150592 301318 150648
rect 301374 150592 301379 150648
rect 301270 150587 301379 150592
rect 284518 150514 284524 150516
rect 267690 150454 284524 150514
rect 264164 150452 264170 150454
rect 264881 150451 264947 150454
rect 284518 150452 284524 150454
rect 284588 150452 284594 150516
rect 288341 150378 288407 150381
rect 288341 150376 290076 150378
rect 288341 150320 288346 150376
rect 288402 150320 290076 150376
rect 301270 150348 301330 150587
rect 288341 150318 290076 150320
rect 288341 150315 288407 150318
rect 266721 150106 266787 150109
rect 263948 150104 266787 150106
rect 263948 150048 266726 150104
rect 266782 150048 266787 150104
rect 263948 150046 266787 150048
rect 266721 150043 266787 150046
rect -960 149834 480 149924
rect 268694 149908 268700 149972
rect 268764 149970 268770 149972
rect 268764 149910 290076 149970
rect 268764 149908 268770 149910
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 249609 149834 249675 149837
rect 249609 149832 252172 149834
rect 249609 149776 249614 149832
rect 249670 149776 252172 149832
rect 249609 149774 252172 149776
rect 249609 149771 249675 149774
rect 272558 149772 272564 149836
rect 272628 149834 272634 149836
rect 288249 149834 288315 149837
rect 272628 149832 288315 149834
rect 272628 149776 288254 149832
rect 288310 149776 288315 149832
rect 272628 149774 288315 149776
rect 272628 149772 272634 149774
rect 288249 149771 288315 149774
rect 266353 149698 266419 149701
rect 263948 149696 266419 149698
rect 263948 149640 266358 149696
rect 266414 149640 266419 149696
rect 263948 149638 266419 149640
rect 266353 149635 266419 149638
rect 266537 149698 266603 149701
rect 283782 149698 283788 149700
rect 266537 149696 283788 149698
rect 266537 149640 266542 149696
rect 266598 149640 283788 149696
rect 266537 149638 283788 149640
rect 266537 149635 266603 149638
rect 283782 149636 283788 149638
rect 283852 149636 283858 149700
rect 303797 149698 303863 149701
rect 301852 149696 303863 149698
rect 301852 149640 303802 149696
rect 303858 149640 303863 149696
rect 301852 149638 303863 149640
rect 303797 149635 303863 149638
rect 285070 149228 285076 149292
rect 285140 149290 285146 149292
rect 290046 149290 290106 149532
rect 285140 149230 290106 149290
rect 285140 149228 285146 149230
rect 248965 149154 249031 149157
rect 265249 149154 265315 149157
rect 248965 149152 252172 149154
rect 248965 149096 248970 149152
rect 249026 149096 252172 149152
rect 248965 149094 252172 149096
rect 263948 149152 265315 149154
rect 263948 149096 265254 149152
rect 265310 149096 265315 149152
rect 263948 149094 265315 149096
rect 248965 149091 249031 149094
rect 265249 149091 265315 149094
rect 288341 149018 288407 149021
rect 288341 149016 290076 149018
rect 288341 148960 288346 149016
rect 288402 148960 290076 149016
rect 288341 148958 290076 148960
rect 288341 148955 288407 148958
rect 303797 148882 303863 148885
rect 301852 148880 303863 148882
rect 301852 148824 303802 148880
rect 303858 148824 303863 148880
rect 301852 148822 303863 148824
rect 303797 148819 303863 148822
rect 266537 148746 266603 148749
rect 263948 148744 266603 148746
rect 263948 148688 266542 148744
rect 266598 148688 266603 148744
rect 263948 148686 266603 148688
rect 266537 148683 266603 148686
rect 282269 148746 282335 148749
rect 288525 148746 288591 148749
rect 282269 148744 288591 148746
rect 282269 148688 282274 148744
rect 282330 148688 288530 148744
rect 288586 148688 288591 148744
rect 282269 148686 288591 148688
rect 282269 148683 282335 148686
rect 288525 148683 288591 148686
rect 287237 148610 287303 148613
rect 287237 148608 290076 148610
rect 287237 148552 287242 148608
rect 287298 148552 290076 148608
rect 287237 148550 290076 148552
rect 287237 148547 287303 148550
rect 249425 148474 249491 148477
rect 249425 148472 252172 148474
rect 249425 148416 249430 148472
rect 249486 148416 252172 148472
rect 249425 148414 252172 148416
rect 249425 148411 249491 148414
rect 266169 148338 266235 148341
rect 266169 148336 290106 148338
rect 266169 148280 266174 148336
rect 266230 148280 290106 148336
rect 266169 148278 290106 148280
rect 266169 148275 266235 148278
rect 266445 148202 266511 148205
rect 263948 148200 266511 148202
rect 263948 148144 266450 148200
rect 266506 148144 266511 148200
rect 290046 148172 290106 148278
rect 263948 148142 266511 148144
rect 266445 148139 266511 148142
rect 304901 148066 304967 148069
rect 301852 148064 304967 148066
rect 301852 148008 304906 148064
rect 304962 148008 304967 148064
rect 301852 148006 304967 148008
rect 304901 148003 304967 148006
rect 249241 147930 249307 147933
rect 288525 147930 288591 147933
rect 249241 147928 252172 147930
rect 249241 147872 249246 147928
rect 249302 147872 252172 147928
rect 249241 147870 252172 147872
rect 288525 147928 290106 147930
rect 288525 147872 288530 147928
rect 288586 147872 290106 147928
rect 288525 147870 290106 147872
rect 249241 147867 249307 147870
rect 288525 147867 288591 147870
rect 267038 147794 267044 147796
rect 263948 147734 267044 147794
rect 267038 147732 267044 147734
rect 267108 147732 267114 147796
rect 290046 147764 290106 147870
rect 288341 147386 288407 147389
rect 303705 147386 303771 147389
rect 288341 147384 290076 147386
rect 288341 147328 288346 147384
rect 288402 147328 290076 147384
rect 288341 147326 290076 147328
rect 301852 147384 303771 147386
rect 301852 147328 303710 147384
rect 303766 147328 303771 147384
rect 301852 147326 303771 147328
rect 288341 147323 288407 147326
rect 303705 147323 303771 147326
rect 249149 147250 249215 147253
rect 266353 147250 266419 147253
rect 249149 147248 252172 147250
rect 249149 147192 249154 147248
rect 249210 147192 252172 147248
rect 249149 147190 252172 147192
rect 263948 147248 266419 147250
rect 263948 147192 266358 147248
rect 266414 147192 266419 147248
rect 263948 147190 266419 147192
rect 249149 147187 249215 147190
rect 266353 147187 266419 147190
rect 280061 147114 280127 147117
rect 287697 147114 287763 147117
rect 280061 147112 287763 147114
rect 280061 147056 280066 147112
rect 280122 147056 287702 147112
rect 287758 147056 287763 147112
rect 280061 147054 287763 147056
rect 280061 147051 280127 147054
rect 287697 147051 287763 147054
rect 301814 147052 301820 147116
rect 301884 147052 301890 147116
rect 287421 146978 287487 146981
rect 287421 146976 290076 146978
rect 287421 146920 287426 146976
rect 287482 146920 290076 146976
rect 287421 146918 290076 146920
rect 287421 146915 287487 146918
rect 263948 146782 267750 146842
rect 249701 146570 249767 146573
rect 249701 146568 252172 146570
rect 249701 146512 249706 146568
rect 249762 146512 252172 146568
rect 249701 146510 252172 146512
rect 249701 146507 249767 146510
rect 267690 146434 267750 146782
rect 301822 146540 301882 147052
rect 281758 146434 281764 146436
rect 267690 146374 281764 146434
rect 281758 146372 281764 146374
rect 281828 146372 281834 146436
rect 287010 146374 290076 146434
rect 264145 146298 264211 146301
rect 263948 146296 264211 146298
rect 263948 146240 264150 146296
rect 264206 146240 264211 146296
rect 263948 146238 264211 146240
rect 264145 146235 264211 146238
rect 249609 145890 249675 145893
rect 268510 145890 268516 145892
rect 249609 145888 252172 145890
rect 249609 145832 249614 145888
rect 249670 145832 252172 145888
rect 249609 145830 252172 145832
rect 263948 145830 268516 145890
rect 249609 145827 249675 145830
rect 268510 145828 268516 145830
rect 268580 145828 268586 145892
rect 271086 145828 271092 145892
rect 271156 145890 271162 145892
rect 287010 145890 287070 146374
rect 288065 146026 288131 146029
rect 288065 146024 290076 146026
rect 288065 145968 288070 146024
rect 288126 145968 290076 146024
rect 288065 145966 290076 145968
rect 288065 145963 288131 145966
rect 303797 145890 303863 145893
rect 271156 145830 287070 145890
rect 301852 145888 303863 145890
rect 301852 145832 303802 145888
rect 303858 145832 303863 145888
rect 301852 145830 303863 145832
rect 271156 145828 271162 145830
rect 303797 145827 303863 145830
rect 268326 145692 268332 145756
rect 268396 145754 268402 145756
rect 287421 145754 287487 145757
rect 268396 145752 287487 145754
rect 268396 145696 287426 145752
rect 287482 145696 287487 145752
rect 268396 145694 287487 145696
rect 268396 145692 268402 145694
rect 287421 145691 287487 145694
rect 264329 145618 264395 145621
rect 284334 145618 284340 145620
rect 264329 145616 284340 145618
rect 264329 145560 264334 145616
rect 264390 145560 284340 145616
rect 264329 145558 284340 145560
rect 264329 145555 264395 145558
rect 284334 145556 284340 145558
rect 284404 145556 284410 145620
rect 288249 145618 288315 145621
rect 288249 145616 290076 145618
rect 288249 145560 288254 145616
rect 288310 145560 290076 145616
rect 288249 145558 290076 145560
rect 288249 145555 288315 145558
rect 264094 145346 264100 145348
rect 263948 145286 264100 145346
rect 264094 145284 264100 145286
rect 264164 145284 264170 145348
rect 249701 145210 249767 145213
rect 287421 145210 287487 145213
rect 249701 145208 252172 145210
rect 249701 145152 249706 145208
rect 249762 145152 252172 145208
rect 249701 145150 252172 145152
rect 287421 145208 290076 145210
rect 287421 145152 287426 145208
rect 287482 145152 290076 145208
rect 287421 145150 290076 145152
rect 249701 145147 249767 145150
rect 287421 145147 287487 145150
rect 303705 145074 303771 145077
rect 301852 145072 303771 145074
rect 301852 145016 303710 145072
rect 303766 145016 303771 145072
rect 301852 145014 303771 145016
rect 303705 145011 303771 145014
rect 267641 144938 267707 144941
rect 263948 144936 267707 144938
rect 263948 144880 267646 144936
rect 267702 144880 267707 144936
rect 263948 144878 267707 144880
rect 267641 144875 267707 144878
rect 267733 144802 267799 144805
rect 271965 144802 272031 144805
rect 267733 144800 272031 144802
rect 267733 144744 267738 144800
rect 267794 144744 271970 144800
rect 272026 144744 272031 144800
rect 267733 144742 272031 144744
rect 267733 144739 267799 144742
rect 271965 144739 272031 144742
rect 278814 144740 278820 144804
rect 278884 144802 278890 144804
rect 280286 144802 280292 144804
rect 278884 144742 280292 144802
rect 278884 144740 278890 144742
rect 280286 144740 280292 144742
rect 280356 144740 280362 144804
rect 288157 144802 288223 144805
rect 288157 144800 290076 144802
rect 288157 144744 288162 144800
rect 288218 144744 290076 144800
rect 288157 144742 290076 144744
rect 288157 144739 288223 144742
rect 249149 144530 249215 144533
rect 249149 144528 252172 144530
rect 249149 144472 249154 144528
rect 249210 144472 252172 144528
rect 249149 144470 252172 144472
rect 249149 144467 249215 144470
rect 287697 144394 287763 144397
rect 263948 144334 267750 144394
rect 266353 143986 266419 143989
rect 263948 143984 266419 143986
rect 263948 143928 266358 143984
rect 266414 143928 266419 143984
rect 263948 143926 266419 143928
rect 266353 143923 266419 143926
rect 249701 143850 249767 143853
rect 249701 143848 252172 143850
rect 249701 143792 249706 143848
rect 249762 143792 252172 143848
rect 249701 143790 252172 143792
rect 249701 143787 249767 143790
rect 267690 143578 267750 144334
rect 287697 144392 290076 144394
rect 287697 144336 287702 144392
rect 287758 144336 290076 144392
rect 287697 144334 290076 144336
rect 287697 144331 287763 144334
rect 303797 144258 303863 144261
rect 301852 144256 303863 144258
rect 301852 144200 303802 144256
rect 303858 144200 303863 144256
rect 301852 144198 303863 144200
rect 303797 144195 303863 144198
rect 279785 143850 279851 143853
rect 279785 143848 290076 143850
rect 279785 143792 279790 143848
rect 279846 143792 290076 143848
rect 279785 143790 290076 143792
rect 279785 143787 279851 143790
rect 280061 143578 280127 143581
rect 309317 143578 309383 143581
rect 267690 143576 280127 143578
rect 267690 143520 280066 143576
rect 280122 143520 280127 143576
rect 267690 143518 280127 143520
rect 301852 143576 309383 143578
rect 301852 143520 309322 143576
rect 309378 143520 309383 143576
rect 301852 143518 309383 143520
rect 280061 143515 280127 143518
rect 309317 143515 309383 143518
rect 266997 143442 267063 143445
rect 263948 143440 267063 143442
rect 263948 143384 267002 143440
rect 267058 143384 267063 143440
rect 263948 143382 267063 143384
rect 266997 143379 267063 143382
rect 184054 142700 184060 142764
rect 184124 142762 184130 142764
rect 243537 142762 243603 142765
rect 252142 142762 252202 143276
rect 280838 143108 280844 143172
rect 280908 143170 280914 143172
rect 290046 143170 290106 143412
rect 280908 143110 290106 143170
rect 280908 143108 280914 143110
rect 266353 143034 266419 143037
rect 263948 143032 266419 143034
rect 263948 142976 266358 143032
rect 266414 142976 266419 143032
rect 263948 142974 266419 142976
rect 266353 142971 266419 142974
rect 287973 143034 288039 143037
rect 287973 143032 290076 143034
rect 287973 142976 287978 143032
rect 288034 142976 290076 143032
rect 287973 142974 290076 142976
rect 287973 142971 288039 142974
rect 184124 142760 243603 142762
rect 184124 142704 243542 142760
rect 243598 142704 243603 142760
rect 184124 142702 243603 142704
rect 184124 142700 184130 142702
rect 243537 142699 243603 142702
rect 248370 142702 252202 142762
rect 188429 142218 188495 142221
rect 248370 142218 248430 142702
rect 267222 142700 267228 142764
rect 267292 142762 267298 142764
rect 282545 142762 282611 142765
rect 306414 142762 306420 142764
rect 267292 142760 282611 142762
rect 267292 142704 282550 142760
rect 282606 142704 282611 142760
rect 267292 142702 282611 142704
rect 301852 142702 306420 142762
rect 267292 142700 267298 142702
rect 282545 142699 282611 142702
rect 306414 142700 306420 142702
rect 306484 142700 306490 142764
rect 249701 142626 249767 142629
rect 287881 142626 287947 142629
rect 249701 142624 252172 142626
rect 249701 142568 249706 142624
rect 249762 142568 252172 142624
rect 249701 142566 252172 142568
rect 287881 142624 290076 142626
rect 287881 142568 287886 142624
rect 287942 142568 290076 142624
rect 287881 142566 290076 142568
rect 249701 142563 249767 142566
rect 287881 142563 287947 142566
rect 265014 142490 265020 142492
rect 263948 142430 265020 142490
rect 265014 142428 265020 142430
rect 265084 142428 265090 142492
rect 315941 142220 316007 142221
rect 188429 142216 248430 142218
rect 188429 142160 188434 142216
rect 188490 142160 248430 142216
rect 188429 142158 248430 142160
rect 188429 142155 188495 142158
rect 286174 142156 286180 142220
rect 286244 142218 286250 142220
rect 315941 142218 315988 142220
rect 286244 142158 290076 142218
rect 315896 142216 315988 142218
rect 316052 142218 316058 142220
rect 315896 142160 315946 142216
rect 315896 142158 315988 142160
rect 286244 142156 286250 142158
rect 315941 142156 315988 142158
rect 316052 142158 316134 142218
rect 316052 142156 316058 142158
rect 315941 142155 316007 142156
rect 265433 142082 265499 142085
rect 303981 142082 304047 142085
rect 315941 142084 316007 142085
rect 315941 142082 315988 142084
rect 263948 142080 265499 142082
rect 263948 142024 265438 142080
rect 265494 142024 265499 142080
rect 263948 142022 265499 142024
rect 301852 142080 304047 142082
rect 301852 142024 303986 142080
rect 304042 142024 304047 142080
rect 301852 142022 304047 142024
rect 315896 142080 315988 142082
rect 316052 142082 316058 142084
rect 315896 142024 315946 142080
rect 315896 142022 315988 142024
rect 265433 142019 265499 142022
rect 303981 142019 304047 142022
rect 315941 142020 315988 142022
rect 316052 142022 316134 142082
rect 316052 142020 316058 142022
rect 315941 142019 316007 142020
rect 249609 141946 249675 141949
rect 249609 141944 252172 141946
rect 249609 141888 249614 141944
rect 249670 141888 252172 141944
rect 249609 141886 252172 141888
rect 249609 141883 249675 141886
rect 264329 141674 264395 141677
rect 263948 141672 264395 141674
rect 263948 141616 264334 141672
rect 264390 141616 264395 141672
rect 263948 141614 264395 141616
rect 264329 141611 264395 141614
rect 213126 141340 213132 141404
rect 213196 141402 213202 141404
rect 222837 141402 222903 141405
rect 213196 141400 222903 141402
rect 213196 141344 222842 141400
rect 222898 141344 222903 141400
rect 213196 141342 222903 141344
rect 213196 141340 213202 141342
rect 222837 141339 222903 141342
rect 273846 141340 273852 141404
rect 273916 141402 273922 141404
rect 290046 141402 290106 141780
rect 273916 141342 290106 141402
rect 273916 141340 273922 141342
rect 249701 141266 249767 141269
rect 287421 141266 287487 141269
rect 303797 141266 303863 141269
rect 249701 141264 252172 141266
rect 249701 141208 249706 141264
rect 249762 141208 252172 141264
rect 249701 141206 252172 141208
rect 287421 141264 290076 141266
rect 287421 141208 287426 141264
rect 287482 141208 290076 141264
rect 287421 141206 290076 141208
rect 301852 141264 303863 141266
rect 301852 141208 303802 141264
rect 303858 141208 303863 141264
rect 301852 141206 303863 141208
rect 249701 141203 249767 141206
rect 287421 141203 287487 141206
rect 303797 141203 303863 141206
rect 263948 141070 267750 141130
rect 267690 140994 267750 141070
rect 277526 140994 277532 140996
rect 267690 140934 277532 140994
rect 277526 140932 277532 140934
rect 277596 140932 277602 140996
rect 283782 140932 283788 140996
rect 283852 140994 283858 140996
rect 283852 140934 290106 140994
rect 283852 140932 283858 140934
rect 265433 140858 265499 140861
rect 273478 140858 273484 140860
rect 265433 140856 273484 140858
rect 265433 140800 265438 140856
rect 265494 140800 273484 140856
rect 265433 140798 273484 140800
rect 265433 140795 265499 140798
rect 273478 140796 273484 140798
rect 273548 140796 273554 140860
rect 290046 140828 290106 140934
rect 269798 140722 269804 140724
rect 263948 140662 269804 140722
rect 269798 140660 269804 140662
rect 269868 140660 269874 140724
rect 249149 140586 249215 140589
rect 249149 140584 252172 140586
rect 249149 140528 249154 140584
rect 249210 140528 252172 140584
rect 249149 140526 252172 140528
rect 249149 140523 249215 140526
rect 288198 140388 288204 140452
rect 288268 140450 288274 140452
rect 302366 140450 302372 140452
rect 288268 140390 290076 140450
rect 301852 140390 302372 140450
rect 288268 140388 288274 140390
rect 302366 140388 302372 140390
rect 302436 140388 302442 140452
rect 263948 140118 267750 140178
rect 248965 139906 249031 139909
rect 248965 139904 252172 139906
rect 248965 139848 248970 139904
rect 249026 139848 252172 139904
rect 248965 139846 252172 139848
rect 248965 139843 249031 139846
rect 264145 139770 264211 139773
rect 263948 139768 264211 139770
rect 263948 139712 264150 139768
rect 264206 139712 264211 139768
rect 263948 139710 264211 139712
rect 264145 139707 264211 139710
rect 267690 139498 267750 140118
rect 270350 139980 270356 140044
rect 270420 140042 270426 140044
rect 288617 140042 288683 140045
rect 270420 140040 288683 140042
rect 270420 139984 288622 140040
rect 288678 139984 288683 140040
rect 270420 139982 288683 139984
rect 270420 139980 270426 139982
rect 288617 139979 288683 139982
rect 282494 139708 282500 139772
rect 282564 139770 282570 139772
rect 290046 139770 290106 140012
rect 303613 139770 303679 139773
rect 282564 139710 290106 139770
rect 301852 139768 303679 139770
rect 301852 139712 303618 139768
rect 303674 139712 303679 139768
rect 301852 139710 303679 139712
rect 282564 139708 282570 139710
rect 303613 139707 303679 139710
rect 287789 139634 287855 139637
rect 287789 139632 290076 139634
rect 287789 139576 287794 139632
rect 287850 139576 290076 139632
rect 287789 139574 290076 139576
rect 287789 139571 287855 139574
rect 285622 139498 285628 139500
rect 267690 139438 285628 139498
rect 285622 139436 285628 139438
rect 285692 139436 285698 139500
rect 583201 139362 583267 139365
rect 583520 139362 584960 139452
rect 583201 139360 584960 139362
rect 583201 139304 583206 139360
rect 583262 139304 584960 139360
rect 583201 139302 584960 139304
rect 583201 139299 583267 139302
rect 249057 139226 249123 139229
rect 288249 139226 288315 139229
rect 249057 139224 252172 139226
rect 249057 139168 249062 139224
rect 249118 139168 252172 139224
rect 249057 139166 252172 139168
rect 263948 139166 267750 139226
rect 249057 139163 249123 139166
rect 266353 138818 266419 138821
rect 263948 138816 266419 138818
rect 263948 138760 266358 138816
rect 266414 138760 266419 138816
rect 263948 138758 266419 138760
rect 266353 138755 266419 138758
rect 249701 138682 249767 138685
rect 249701 138680 252172 138682
rect 249701 138624 249706 138680
rect 249762 138624 252172 138680
rect 249701 138622 252172 138624
rect 249701 138619 249767 138622
rect 267690 138410 267750 139166
rect 288249 139224 290076 139226
rect 288249 139168 288254 139224
rect 288310 139168 290076 139224
rect 583520 139212 584960 139302
rect 288249 139166 290076 139168
rect 288249 139163 288315 139166
rect 304257 138954 304323 138957
rect 301852 138952 304323 138954
rect 301852 138896 304262 138952
rect 304318 138896 304323 138952
rect 301852 138894 304323 138896
rect 304257 138891 304323 138894
rect 269798 138620 269804 138684
rect 269868 138682 269874 138684
rect 283833 138682 283899 138685
rect 269868 138680 283899 138682
rect 269868 138624 283838 138680
rect 283894 138624 283899 138680
rect 269868 138622 283899 138624
rect 269868 138620 269874 138622
rect 283833 138619 283899 138622
rect 289353 138682 289419 138685
rect 289353 138680 290076 138682
rect 289353 138624 289358 138680
rect 289414 138624 290076 138680
rect 289353 138622 290076 138624
rect 289353 138619 289419 138622
rect 288382 138410 288388 138412
rect 267690 138350 288388 138410
rect 288382 138348 288388 138350
rect 288452 138348 288458 138412
rect 270350 138274 270356 138276
rect 263948 138214 270356 138274
rect 270350 138212 270356 138214
rect 270420 138212 270426 138276
rect 288341 138274 288407 138277
rect 303797 138274 303863 138277
rect 288341 138272 290076 138274
rect 288341 138216 288346 138272
rect 288402 138216 290076 138272
rect 288341 138214 290076 138216
rect 301852 138272 303863 138274
rect 301852 138216 303802 138272
rect 303858 138216 303863 138272
rect 301852 138214 303863 138216
rect 288341 138211 288407 138214
rect 303797 138211 303863 138214
rect 249149 138002 249215 138005
rect 249149 138000 252172 138002
rect 249149 137944 249154 138000
rect 249210 137944 252172 138000
rect 249149 137942 252172 137944
rect 249149 137939 249215 137942
rect 290590 137940 290596 138004
rect 290660 137940 290666 138004
rect 270534 137866 270540 137868
rect 263948 137806 270540 137866
rect 270534 137804 270540 137806
rect 270604 137804 270610 137868
rect 290598 137836 290658 137940
rect 288341 137458 288407 137461
rect 303797 137458 303863 137461
rect 288341 137456 290076 137458
rect 288341 137400 288346 137456
rect 288402 137400 290076 137456
rect 288341 137398 290076 137400
rect 301852 137456 303863 137458
rect 301852 137400 303802 137456
rect 303858 137400 303863 137456
rect 301852 137398 303863 137400
rect 288341 137395 288407 137398
rect 303797 137395 303863 137398
rect 249701 137322 249767 137325
rect 265433 137322 265499 137325
rect 249701 137320 252172 137322
rect 249701 137264 249706 137320
rect 249762 137264 252172 137320
rect 249701 137262 252172 137264
rect 263948 137320 265499 137322
rect 263948 137264 265438 137320
rect 265494 137264 265499 137320
rect 263948 137262 265499 137264
rect 249701 137259 249767 137262
rect 265433 137259 265499 137262
rect 287094 137050 287100 137052
rect 282134 136990 287100 137050
rect 281574 136914 281580 136916
rect -960 136778 480 136868
rect 263948 136854 281580 136914
rect 281574 136852 281580 136854
rect 281644 136852 281650 136916
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 265433 136778 265499 136781
rect 282134 136778 282194 136990
rect 287094 136988 287100 136990
rect 287164 136988 287170 137052
rect 288574 136990 290076 137050
rect 282310 136852 282316 136916
rect 282380 136914 282386 136916
rect 288574 136914 288634 136990
rect 282380 136854 288634 136914
rect 282380 136852 282386 136854
rect 265433 136776 282194 136778
rect 265433 136720 265438 136776
rect 265494 136720 282194 136776
rect 265433 136718 282194 136720
rect 265433 136715 265499 136718
rect 249149 136642 249215 136645
rect 289445 136642 289511 136645
rect 302182 136642 302188 136644
rect 249149 136640 252172 136642
rect 249149 136584 249154 136640
rect 249210 136584 252172 136640
rect 249149 136582 252172 136584
rect 289445 136640 290076 136642
rect 289445 136584 289450 136640
rect 289506 136584 290076 136640
rect 289445 136582 290076 136584
rect 301852 136582 302188 136642
rect 249149 136579 249215 136582
rect 289445 136579 289511 136582
rect 302182 136580 302188 136582
rect 302252 136580 302258 136644
rect 263948 136310 267750 136370
rect 249701 135962 249767 135965
rect 266353 135962 266419 135965
rect 249701 135960 252172 135962
rect 249701 135904 249706 135960
rect 249762 135904 252172 135960
rect 249701 135902 252172 135904
rect 263948 135960 266419 135962
rect 263948 135904 266358 135960
rect 266414 135904 266419 135960
rect 263948 135902 266419 135904
rect 249701 135899 249767 135902
rect 266353 135899 266419 135902
rect 231301 135554 231367 135557
rect 231301 135552 252202 135554
rect 231301 135496 231306 135552
rect 231362 135496 252202 135552
rect 231301 135494 252202 135496
rect 231301 135491 231367 135494
rect 252142 135252 252202 135494
rect 266353 135418 266419 135421
rect 263948 135416 266419 135418
rect 263948 135360 266358 135416
rect 266414 135360 266419 135416
rect 263948 135358 266419 135360
rect 266353 135355 266419 135358
rect 267690 135282 267750 136310
rect 289261 136234 289327 136237
rect 289261 136232 290076 136234
rect 289261 136176 289266 136232
rect 289322 136176 290076 136232
rect 289261 136174 290076 136176
rect 289261 136171 289327 136174
rect 303613 135962 303679 135965
rect 301852 135960 303679 135962
rect 301852 135904 303618 135960
rect 303674 135904 303679 135960
rect 301852 135902 303679 135904
rect 303613 135899 303679 135902
rect 278630 135628 278636 135692
rect 278700 135690 278706 135692
rect 278700 135630 290076 135690
rect 278700 135628 278706 135630
rect 284886 135356 284892 135420
rect 284956 135418 284962 135420
rect 284956 135358 290106 135418
rect 284956 135356 284962 135358
rect 278814 135282 278820 135284
rect 267690 135222 278820 135282
rect 278814 135220 278820 135222
rect 278884 135220 278890 135284
rect 290046 135252 290106 135358
rect 266445 135010 266511 135013
rect 263948 135008 266511 135010
rect 263948 134952 266450 135008
rect 266506 134952 266511 135008
rect 263948 134950 266511 134952
rect 266445 134947 266511 134950
rect 287830 134812 287836 134876
rect 287900 134874 287906 134876
rect 287900 134814 290076 134874
rect 287900 134812 287906 134814
rect 249701 134602 249767 134605
rect 266997 134602 267063 134605
rect 278630 134602 278636 134604
rect 249701 134600 252172 134602
rect 249701 134544 249706 134600
rect 249762 134544 252172 134600
rect 249701 134542 252172 134544
rect 266997 134600 278636 134602
rect 266997 134544 267002 134600
rect 267058 134544 278636 134600
rect 266997 134542 278636 134544
rect 249701 134539 249767 134542
rect 266997 134539 267063 134542
rect 278630 134540 278636 134542
rect 278700 134540 278706 134604
rect 301822 134602 301882 135116
rect 313457 134602 313523 134605
rect 301822 134600 313523 134602
rect 301822 134544 313462 134600
rect 313518 134544 313523 134600
rect 301822 134542 313523 134544
rect 313457 134539 313523 134542
rect 266353 134466 266419 134469
rect 263948 134464 266419 134466
rect 263948 134408 266358 134464
rect 266414 134408 266419 134464
rect 263948 134406 266419 134408
rect 266353 134403 266419 134406
rect 271638 134404 271644 134468
rect 271708 134466 271714 134468
rect 288198 134466 288204 134468
rect 271708 134406 288204 134466
rect 271708 134404 271714 134406
rect 288198 134404 288204 134406
rect 288268 134404 288274 134468
rect 303705 134466 303771 134469
rect 301852 134464 303771 134466
rect 277894 134132 277900 134196
rect 277964 134194 277970 134196
rect 290046 134194 290106 134436
rect 301852 134408 303710 134464
rect 303766 134408 303771 134464
rect 301852 134406 303771 134408
rect 303705 134403 303771 134406
rect 277964 134134 290106 134194
rect 277964 134132 277970 134134
rect 267089 134058 267155 134061
rect 263948 134056 267155 134058
rect 263948 134000 267094 134056
rect 267150 134000 267155 134056
rect 263948 133998 267155 134000
rect 267089 133995 267155 133998
rect 240869 133922 240935 133925
rect 240869 133920 252172 133922
rect 240869 133864 240874 133920
rect 240930 133864 252172 133920
rect 240869 133862 252172 133864
rect 240869 133859 240935 133862
rect 290230 133788 290290 134028
rect 290222 133724 290228 133788
rect 290292 133724 290298 133788
rect 287145 133650 287211 133653
rect 303797 133650 303863 133653
rect 287145 133648 290076 133650
rect 287145 133592 287150 133648
rect 287206 133592 290076 133648
rect 287145 133590 290076 133592
rect 301852 133648 303863 133650
rect 301852 133592 303802 133648
rect 303858 133592 303863 133648
rect 301852 133590 303863 133592
rect 287145 133587 287211 133590
rect 303797 133587 303863 133590
rect 267181 133514 267247 133517
rect 263948 133512 267247 133514
rect 263948 133456 267186 133512
rect 267242 133456 267247 133512
rect 263948 133454 267247 133456
rect 267181 133451 267247 133454
rect 212390 133044 212396 133108
rect 212460 133106 212466 133108
rect 234061 133106 234127 133109
rect 212460 133104 234127 133106
rect 212460 133048 234066 133104
rect 234122 133048 234127 133104
rect 212460 133046 234127 133048
rect 212460 133044 212466 133046
rect 234061 133043 234127 133046
rect 247769 132834 247835 132837
rect 252142 132834 252202 133348
rect 266353 133106 266419 133109
rect 263948 133104 266419 133106
rect 263948 133048 266358 133104
rect 266414 133048 266419 133104
rect 263948 133046 266419 133048
rect 266353 133043 266419 133046
rect 288341 133106 288407 133109
rect 288341 133104 290076 133106
rect 288341 133048 288346 133104
rect 288402 133048 290076 133104
rect 288341 133046 290076 133048
rect 288341 133043 288407 133046
rect 247769 132832 252202 132834
rect 247769 132776 247774 132832
rect 247830 132776 252202 132832
rect 247769 132774 252202 132776
rect 247769 132771 247835 132774
rect 265750 132772 265756 132836
rect 265820 132834 265826 132836
rect 303889 132834 303955 132837
rect 265820 132774 290106 132834
rect 301852 132832 303955 132834
rect 301852 132776 303894 132832
rect 303950 132776 303955 132832
rect 301852 132774 303955 132776
rect 265820 132772 265826 132774
rect 250302 132638 252172 132698
rect 290046 132668 290106 132774
rect 303889 132771 303955 132774
rect 206277 132562 206343 132565
rect 250302 132562 250362 132638
rect 315982 132636 315988 132700
rect 316052 132636 316058 132700
rect 315990 132565 316050 132636
rect 266353 132562 266419 132565
rect 315941 132562 316050 132565
rect 206277 132560 250362 132562
rect 206277 132504 206282 132560
rect 206338 132504 250362 132560
rect 206277 132502 250362 132504
rect 263948 132560 266419 132562
rect 263948 132504 266358 132560
rect 266414 132504 266419 132560
rect 263948 132502 266419 132504
rect 315896 132560 316050 132562
rect 315896 132504 315946 132560
rect 316002 132504 316050 132560
rect 315896 132502 316050 132504
rect 206277 132499 206343 132502
rect 266353 132499 266419 132502
rect 315941 132499 316007 132502
rect 278313 132426 278379 132429
rect 315941 132428 316007 132429
rect 315941 132426 315988 132428
rect 267690 132424 278379 132426
rect 267690 132368 278318 132424
rect 278374 132368 278379 132424
rect 267690 132366 278379 132368
rect 315896 132424 315988 132426
rect 316052 132426 316058 132428
rect 315896 132368 315946 132424
rect 315896 132366 315988 132368
rect 267690 132154 267750 132366
rect 278313 132363 278379 132366
rect 315941 132364 315988 132366
rect 316052 132366 316134 132426
rect 316052 132364 316058 132366
rect 315941 132363 316007 132364
rect 288341 132290 288407 132293
rect 288341 132288 290076 132290
rect 288341 132232 288346 132288
rect 288402 132232 290076 132288
rect 288341 132230 290076 132232
rect 288341 132227 288407 132230
rect 303797 132154 303863 132157
rect 263948 132094 267750 132154
rect 301852 132152 303863 132154
rect 301852 132096 303802 132152
rect 303858 132096 303863 132152
rect 301852 132094 303863 132096
rect 303797 132091 303863 132094
rect 249701 132018 249767 132021
rect 249701 132016 252172 132018
rect 249701 131960 249706 132016
rect 249762 131960 252172 132016
rect 249701 131958 252172 131960
rect 249701 131955 249767 131958
rect 275645 131746 275711 131749
rect 282494 131746 282500 131748
rect 275645 131744 282500 131746
rect 275645 131688 275650 131744
rect 275706 131688 282500 131744
rect 275645 131686 282500 131688
rect 275645 131683 275711 131686
rect 282494 131684 282500 131686
rect 282564 131684 282570 131748
rect 266353 131610 266419 131613
rect 290046 131610 290106 131852
rect 263948 131608 266419 131610
rect 263948 131552 266358 131608
rect 266414 131552 266419 131608
rect 263948 131550 266419 131552
rect 266353 131547 266419 131550
rect 267690 131550 290106 131610
rect 264881 131474 264947 131477
rect 267690 131474 267750 131550
rect 264881 131472 267750 131474
rect 264881 131416 264886 131472
rect 264942 131416 267750 131472
rect 264881 131414 267750 131416
rect 264881 131411 264947 131414
rect 289118 131412 289124 131476
rect 289188 131474 289194 131476
rect 289188 131414 290076 131474
rect 289188 131412 289194 131414
rect 249241 131338 249307 131341
rect 303889 131338 303955 131341
rect 249241 131336 252172 131338
rect 249241 131280 249246 131336
rect 249302 131280 252172 131336
rect 249241 131278 252172 131280
rect 301852 131336 303955 131338
rect 301852 131280 303894 131336
rect 303950 131280 303955 131336
rect 301852 131278 303955 131280
rect 249241 131275 249307 131278
rect 303889 131275 303955 131278
rect 266445 131202 266511 131205
rect 263948 131200 266511 131202
rect 263948 131144 266450 131200
rect 266506 131144 266511 131200
rect 263948 131142 266511 131144
rect 266445 131139 266511 131142
rect 266353 131066 266419 131069
rect 286409 131066 286475 131069
rect 266353 131064 286475 131066
rect 266353 131008 266358 131064
rect 266414 131008 286414 131064
rect 286470 131008 286475 131064
rect 266353 131006 286475 131008
rect 266353 131003 266419 131006
rect 286409 131003 286475 131006
rect 289169 131066 289235 131069
rect 289169 131064 290076 131066
rect 289169 131008 289174 131064
rect 289230 131008 290076 131064
rect 289169 131006 290076 131008
rect 289169 131003 289235 131006
rect 249609 130658 249675 130661
rect 272701 130658 272767 130661
rect 303797 130658 303863 130661
rect 249609 130656 252172 130658
rect 249609 130600 249614 130656
rect 249670 130600 252172 130656
rect 249609 130598 252172 130600
rect 263948 130656 272767 130658
rect 263948 130600 272706 130656
rect 272762 130600 272767 130656
rect 263948 130598 272767 130600
rect 301852 130656 303863 130658
rect 301852 130600 303802 130656
rect 303858 130600 303863 130656
rect 301852 130598 303863 130600
rect 249609 130595 249675 130598
rect 272701 130595 272767 130598
rect 303797 130595 303863 130598
rect 288341 130522 288407 130525
rect 288341 130520 290076 130522
rect 288341 130464 288346 130520
rect 288402 130464 290076 130520
rect 288341 130462 290076 130464
rect 288341 130459 288407 130462
rect 286542 130324 286548 130388
rect 286612 130386 286618 130388
rect 289353 130386 289419 130389
rect 286612 130384 289419 130386
rect 286612 130328 289358 130384
rect 289414 130328 289419 130384
rect 286612 130326 289419 130328
rect 286612 130324 286618 130326
rect 289353 130323 289419 130326
rect 266353 130250 266419 130253
rect 263948 130248 266419 130250
rect 263948 130192 266358 130248
rect 266414 130192 266419 130248
rect 263948 130190 266419 130192
rect 266353 130187 266419 130190
rect 277350 130054 290076 130114
rect 249701 129978 249767 129981
rect 271781 129978 271847 129981
rect 277350 129978 277410 130054
rect 249701 129976 252172 129978
rect 249701 129920 249706 129976
rect 249762 129920 252172 129976
rect 249701 129918 252172 129920
rect 271781 129976 277410 129978
rect 271781 129920 271786 129976
rect 271842 129920 277410 129976
rect 271781 129918 277410 129920
rect 249701 129915 249767 129918
rect 271781 129915 271847 129918
rect 266445 129842 266511 129845
rect 305177 129842 305243 129845
rect 263948 129840 266511 129842
rect 263948 129784 266450 129840
rect 266506 129784 266511 129840
rect 263948 129782 266511 129784
rect 301852 129840 305243 129842
rect 301852 129784 305182 129840
rect 305238 129784 305243 129840
rect 301852 129782 305243 129784
rect 266445 129779 266511 129782
rect 305177 129779 305243 129782
rect 288065 129706 288131 129709
rect 288065 129704 290076 129706
rect 288065 129648 288070 129704
rect 288126 129648 290076 129704
rect 288065 129646 290076 129648
rect 288065 129643 288131 129646
rect 67357 129298 67423 129301
rect 68142 129298 68816 129304
rect 67357 129296 68816 129298
rect 67357 129240 67362 129296
rect 67418 129244 68816 129296
rect 249701 129298 249767 129301
rect 266353 129298 266419 129301
rect 249701 129296 252172 129298
rect 67418 129240 68202 129244
rect 67357 129238 68202 129240
rect 249701 129240 249706 129296
rect 249762 129240 252172 129296
rect 249701 129238 252172 129240
rect 263948 129296 266419 129298
rect 263948 129240 266358 129296
rect 266414 129240 266419 129296
rect 263948 129238 266419 129240
rect 67357 129235 67423 129238
rect 249701 129235 249767 129238
rect 266353 129235 266419 129238
rect 287973 129298 288039 129301
rect 287973 129296 290076 129298
rect 287973 129240 287978 129296
rect 288034 129240 290076 129296
rect 287973 129238 290076 129240
rect 287973 129235 288039 129238
rect 303797 129026 303863 129029
rect 301852 129024 303863 129026
rect 301852 128968 303802 129024
rect 303858 128968 303863 129024
rect 301852 128966 303863 128968
rect 303797 128963 303863 128966
rect 266537 128890 266603 128893
rect 263948 128888 266603 128890
rect 263948 128832 266542 128888
rect 266598 128832 266603 128888
rect 263948 128830 266603 128832
rect 266537 128827 266603 128830
rect 289854 128828 289860 128892
rect 289924 128890 289930 128892
rect 289924 128830 290076 128890
rect 289924 128828 289930 128830
rect 250621 128754 250687 128757
rect 250621 128752 252172 128754
rect 250621 128696 250626 128752
rect 250682 128696 252172 128752
rect 250621 128694 252172 128696
rect 250621 128691 250687 128694
rect 287646 128420 287652 128484
rect 287716 128482 287722 128484
rect 287716 128422 290076 128482
rect 287716 128420 287722 128422
rect 282177 128346 282243 128349
rect 263948 128344 282243 128346
rect 263948 128288 282182 128344
rect 282238 128288 282243 128344
rect 263948 128286 282243 128288
rect 282177 128283 282243 128286
rect 282310 128284 282316 128348
rect 282380 128346 282386 128348
rect 287145 128346 287211 128349
rect 303797 128346 303863 128349
rect 282380 128344 287211 128346
rect 282380 128288 287150 128344
rect 287206 128288 287211 128344
rect 282380 128286 287211 128288
rect 301852 128344 303863 128346
rect 301852 128288 303802 128344
rect 303858 128288 303863 128344
rect 301852 128286 303863 128288
rect 282380 128284 282386 128286
rect 287145 128283 287211 128286
rect 303797 128283 303863 128286
rect 266537 128210 266603 128213
rect 269614 128210 269620 128212
rect 266537 128208 269620 128210
rect 266537 128152 266542 128208
rect 266598 128152 269620 128208
rect 266537 128150 269620 128152
rect 266537 128147 266603 128150
rect 269614 128148 269620 128150
rect 269684 128148 269690 128212
rect 67725 128074 67791 128077
rect 68142 128074 68816 128080
rect 67725 128072 68816 128074
rect 67725 128016 67730 128072
rect 67786 128020 68816 128072
rect 249609 128074 249675 128077
rect 249609 128072 252172 128074
rect 67786 128016 68202 128020
rect 67725 128014 68202 128016
rect 249609 128016 249614 128072
rect 249670 128016 252172 128072
rect 249609 128014 252172 128016
rect 67725 128011 67791 128014
rect 249609 128011 249675 128014
rect 264145 127938 264211 127941
rect 263948 127936 264211 127938
rect 263948 127880 264150 127936
rect 264206 127880 264211 127936
rect 263948 127878 264211 127880
rect 264145 127875 264211 127878
rect 287973 127938 288039 127941
rect 287973 127936 290076 127938
rect 287973 127880 287978 127936
rect 288034 127880 290076 127936
rect 287973 127878 290076 127880
rect 287973 127875 288039 127878
rect 288157 127530 288223 127533
rect 303613 127530 303679 127533
rect 288157 127528 290076 127530
rect 288157 127472 288162 127528
rect 288218 127472 290076 127528
rect 288157 127470 290076 127472
rect 301852 127528 303679 127530
rect 301852 127472 303618 127528
rect 303674 127472 303679 127528
rect 301852 127470 303679 127472
rect 288157 127467 288223 127470
rect 303613 127467 303679 127470
rect 249701 127394 249767 127397
rect 266353 127394 266419 127397
rect 249701 127392 252172 127394
rect 249701 127336 249706 127392
rect 249762 127336 252172 127392
rect 249701 127334 252172 127336
rect 263948 127392 266419 127394
rect 263948 127336 266358 127392
rect 266414 127336 266419 127392
rect 263948 127334 266419 127336
rect 249701 127331 249767 127334
rect 266353 127331 266419 127334
rect 270350 127060 270356 127124
rect 270420 127122 270426 127124
rect 270420 127062 290076 127122
rect 270420 127060 270426 127062
rect 272609 126986 272675 126989
rect 263948 126984 272675 126986
rect 263948 126928 272614 126984
rect 272670 126928 272675 126984
rect 263948 126926 272675 126928
rect 272609 126923 272675 126926
rect 308622 126850 308628 126852
rect 301852 126790 308628 126850
rect 308622 126788 308628 126790
rect 308692 126788 308698 126852
rect 249609 126714 249675 126717
rect 249609 126712 252172 126714
rect 249609 126656 249614 126712
rect 249670 126656 252172 126712
rect 249609 126654 252172 126656
rect 249609 126651 249675 126654
rect 265709 126442 265775 126445
rect 290046 126442 290106 126684
rect 263948 126440 265775 126442
rect 263948 126384 265714 126440
rect 265770 126384 265775 126440
rect 263948 126382 265775 126384
rect 265709 126379 265775 126382
rect 277350 126382 290106 126442
rect 66161 126306 66227 126309
rect 68142 126306 68816 126312
rect 66161 126304 68816 126306
rect 66161 126248 66166 126304
rect 66222 126252 68816 126304
rect 66222 126248 68202 126252
rect 66161 126246 68202 126248
rect 66161 126243 66227 126246
rect 277350 126037 277410 126382
rect 288249 126306 288315 126309
rect 288249 126304 290076 126306
rect 288249 126248 288254 126304
rect 288310 126248 290076 126304
rect 288249 126246 290076 126248
rect 288249 126243 288315 126246
rect 249701 126034 249767 126037
rect 266353 126034 266419 126037
rect 249701 126032 252172 126034
rect 249701 125976 249706 126032
rect 249762 125976 252172 126032
rect 249701 125974 252172 125976
rect 263948 126032 266419 126034
rect 263948 125976 266358 126032
rect 266414 125976 266419 126032
rect 263948 125974 266419 125976
rect 249701 125971 249767 125974
rect 266353 125971 266419 125974
rect 277301 126032 277410 126037
rect 304717 126034 304783 126037
rect 277301 125976 277306 126032
rect 277362 125976 277410 126032
rect 277301 125974 277410 125976
rect 301852 126032 304783 126034
rect 301852 125976 304722 126032
rect 304778 125976 304783 126032
rect 301852 125974 304783 125976
rect 277301 125971 277367 125974
rect 304717 125971 304783 125974
rect 580901 126034 580967 126037
rect 583520 126034 584960 126124
rect 580901 126032 584960 126034
rect 580901 125976 580906 126032
rect 580962 125976 584960 126032
rect 580901 125974 584960 125976
rect 580901 125971 580967 125974
rect 288341 125898 288407 125901
rect 288341 125896 290076 125898
rect 288341 125840 288346 125896
rect 288402 125840 290076 125896
rect 583520 125884 584960 125974
rect 288341 125838 290076 125840
rect 288341 125835 288407 125838
rect 266353 125490 266419 125493
rect 263948 125488 266419 125490
rect 263948 125432 266358 125488
rect 266414 125432 266419 125488
rect 263948 125430 266419 125432
rect 266353 125427 266419 125430
rect 249609 125354 249675 125357
rect 288341 125354 288407 125357
rect 249609 125352 252172 125354
rect 249609 125296 249614 125352
rect 249670 125296 252172 125352
rect 249609 125294 252172 125296
rect 288341 125352 290076 125354
rect 288341 125296 288346 125352
rect 288402 125296 290076 125352
rect 288341 125294 290076 125296
rect 249609 125291 249675 125294
rect 288341 125291 288407 125294
rect 67449 125218 67515 125221
rect 68142 125218 68816 125224
rect 302233 125218 302299 125221
rect 67449 125216 68816 125218
rect 67449 125160 67454 125216
rect 67510 125164 68816 125216
rect 301852 125216 302299 125218
rect 67510 125160 68202 125164
rect 67449 125158 68202 125160
rect 301852 125160 302238 125216
rect 302294 125160 302299 125216
rect 301852 125158 302299 125160
rect 67449 125155 67515 125158
rect 302233 125155 302299 125158
rect 266445 125082 266511 125085
rect 263948 125080 266511 125082
rect 263948 125024 266450 125080
rect 266506 125024 266511 125080
rect 263948 125022 266511 125024
rect 266445 125019 266511 125022
rect 268929 124810 268995 124813
rect 288065 124810 288131 124813
rect 268929 124808 288131 124810
rect 268929 124752 268934 124808
rect 268990 124752 288070 124808
rect 288126 124752 288131 124808
rect 268929 124750 288131 124752
rect 268929 124747 268995 124750
rect 288065 124747 288131 124750
rect 249701 124674 249767 124677
rect 274081 124674 274147 124677
rect 290046 124674 290106 124916
rect 249701 124672 252172 124674
rect 249701 124616 249706 124672
rect 249762 124616 252172 124672
rect 249701 124614 252172 124616
rect 274081 124672 290106 124674
rect 274081 124616 274086 124672
rect 274142 124616 290106 124672
rect 274081 124614 290106 124616
rect 249701 124611 249767 124614
rect 274081 124611 274147 124614
rect 267222 124538 267228 124540
rect 263948 124478 267228 124538
rect 267222 124476 267228 124478
rect 267292 124476 267298 124540
rect 287145 124538 287211 124541
rect 303705 124538 303771 124541
rect 287145 124536 290076 124538
rect 287145 124480 287150 124536
rect 287206 124480 290076 124536
rect 287145 124478 290076 124480
rect 301852 124536 303771 124538
rect 301852 124480 303710 124536
rect 303766 124480 303771 124536
rect 301852 124478 303771 124480
rect 287145 124475 287211 124478
rect 303705 124475 303771 124478
rect 248965 124130 249031 124133
rect 266537 124130 266603 124133
rect 248965 124128 252172 124130
rect 248965 124072 248970 124128
rect 249026 124072 252172 124128
rect 248965 124070 252172 124072
rect 263948 124128 266603 124130
rect 263948 124072 266542 124128
rect 266598 124072 266603 124128
rect 263948 124070 266603 124072
rect 248965 124067 249031 124070
rect 266537 124067 266603 124070
rect 287973 124130 288039 124133
rect 287973 124128 290076 124130
rect 287973 124072 287978 124128
rect 288034 124072 290076 124128
rect 287973 124070 290076 124072
rect 287973 124067 288039 124070
rect 265709 123858 265775 123861
rect 288525 123858 288591 123861
rect 265709 123856 288591 123858
rect -960 123572 480 123812
rect 265709 123800 265714 123856
rect 265770 123800 288530 123856
rect 288586 123800 288591 123856
rect 265709 123798 288591 123800
rect 265709 123795 265775 123798
rect 288525 123795 288591 123798
rect 287697 123722 287763 123725
rect 303797 123722 303863 123725
rect 287697 123720 290076 123722
rect 287697 123664 287702 123720
rect 287758 123664 290076 123720
rect 287697 123662 290076 123664
rect 301852 123720 303863 123722
rect 301852 123664 303802 123720
rect 303858 123664 303863 123720
rect 301852 123662 303863 123664
rect 287697 123659 287763 123662
rect 303797 123659 303863 123662
rect 66069 123586 66135 123589
rect 68142 123586 68816 123592
rect 266854 123586 266860 123588
rect 66069 123584 68816 123586
rect 66069 123528 66074 123584
rect 66130 123532 68816 123584
rect 66130 123528 68202 123532
rect 66069 123526 68202 123528
rect 263948 123526 266860 123586
rect 66069 123523 66135 123526
rect 266854 123524 266860 123526
rect 266924 123524 266930 123588
rect 249517 123450 249583 123453
rect 266629 123450 266695 123453
rect 274030 123450 274036 123452
rect 249517 123448 252172 123450
rect 249517 123392 249522 123448
rect 249578 123392 252172 123448
rect 249517 123390 252172 123392
rect 266629 123448 274036 123450
rect 266629 123392 266634 123448
rect 266690 123392 274036 123448
rect 266629 123390 274036 123392
rect 249517 123387 249583 123390
rect 266629 123387 266695 123390
rect 274030 123388 274036 123390
rect 274100 123388 274106 123452
rect 304349 123450 304415 123453
rect 309225 123450 309291 123453
rect 304349 123448 309291 123450
rect 304349 123392 304354 123448
rect 304410 123392 309230 123448
rect 309286 123392 309291 123448
rect 304349 123390 309291 123392
rect 304349 123387 304415 123390
rect 309225 123387 309291 123390
rect 286409 123314 286475 123317
rect 286409 123312 290076 123314
rect 286409 123256 286414 123312
rect 286470 123256 290076 123312
rect 286409 123254 290076 123256
rect 286409 123251 286475 123254
rect 266353 123178 266419 123181
rect 263948 123176 266419 123178
rect 263948 123120 266358 123176
rect 266414 123120 266419 123176
rect 263948 123118 266419 123120
rect 266353 123115 266419 123118
rect 288525 123042 288591 123045
rect 303705 123042 303771 123045
rect 288525 123040 290106 123042
rect 288525 122984 288530 123040
rect 288586 122984 290106 123040
rect 288525 122982 290106 122984
rect 301852 123040 303771 123042
rect 301852 122984 303710 123040
rect 303766 122984 303771 123040
rect 301852 122982 303771 122984
rect 288525 122979 288591 122982
rect 290046 122876 290106 122982
rect 303705 122979 303771 122982
rect 315982 122980 315988 123044
rect 316052 122980 316058 123044
rect 315990 122909 316050 122980
rect 315941 122906 316050 122909
rect 315896 122904 316050 122906
rect 315896 122848 315946 122904
rect 316002 122848 316050 122904
rect 315896 122846 316050 122848
rect 315941 122843 316007 122846
rect 249701 122770 249767 122773
rect 315941 122772 316007 122773
rect 315941 122770 315988 122772
rect 249701 122768 252172 122770
rect 249701 122712 249706 122768
rect 249762 122712 252172 122768
rect 249701 122710 252172 122712
rect 315896 122768 315988 122770
rect 316052 122770 316058 122772
rect 315896 122712 315946 122768
rect 315896 122710 315988 122712
rect 249701 122707 249767 122710
rect 315941 122708 315988 122710
rect 316052 122710 316134 122770
rect 316052 122708 316058 122710
rect 315941 122707 316007 122708
rect 67541 122634 67607 122637
rect 68142 122634 68816 122640
rect 266353 122634 266419 122637
rect 67541 122632 68816 122634
rect 67541 122576 67546 122632
rect 67602 122580 68816 122632
rect 263948 122632 266419 122634
rect 67602 122576 68202 122580
rect 67541 122574 68202 122576
rect 263948 122576 266358 122632
rect 266414 122576 266419 122632
rect 263948 122574 266419 122576
rect 67541 122571 67607 122574
rect 266353 122571 266419 122574
rect 266537 122226 266603 122229
rect 263948 122224 266603 122226
rect 263948 122168 266542 122224
rect 266598 122168 266603 122224
rect 263948 122166 266603 122168
rect 266537 122163 266603 122166
rect 268653 122226 268719 122229
rect 282310 122226 282316 122228
rect 268653 122224 282316 122226
rect 268653 122168 268658 122224
rect 268714 122168 282316 122224
rect 268653 122166 282316 122168
rect 268653 122163 268719 122166
rect 282310 122164 282316 122166
rect 282380 122164 282386 122228
rect 282453 122226 282519 122229
rect 289445 122226 289511 122229
rect 282453 122224 289511 122226
rect 282453 122168 282458 122224
rect 282514 122168 289450 122224
rect 289506 122168 289511 122224
rect 282453 122166 289511 122168
rect 282453 122163 282519 122166
rect 289445 122163 289511 122166
rect 248781 122090 248847 122093
rect 248781 122088 252172 122090
rect 248781 122032 248786 122088
rect 248842 122032 252172 122088
rect 248781 122030 252172 122032
rect 248781 122027 248847 122030
rect 266854 122028 266860 122092
rect 266924 122090 266930 122092
rect 283833 122090 283899 122093
rect 290046 122090 290106 122332
rect 303613 122226 303679 122229
rect 301852 122224 303679 122226
rect 301852 122168 303618 122224
rect 303674 122168 303679 122224
rect 301852 122166 303679 122168
rect 303613 122163 303679 122166
rect 266924 122088 283899 122090
rect 266924 122032 283838 122088
rect 283894 122032 283899 122088
rect 266924 122030 283899 122032
rect 266924 122028 266930 122030
rect 283833 122027 283899 122030
rect 288574 122030 290106 122090
rect 266905 121682 266971 121685
rect 263948 121680 266971 121682
rect 263948 121624 266910 121680
rect 266966 121624 266971 121680
rect 263948 121622 266971 121624
rect 266905 121619 266971 121622
rect 273294 121620 273300 121684
rect 273364 121682 273370 121684
rect 274541 121682 274607 121685
rect 273364 121680 274607 121682
rect 273364 121624 274546 121680
rect 274602 121624 274607 121680
rect 273364 121622 274607 121624
rect 273364 121620 273370 121622
rect 274541 121619 274607 121622
rect 286685 121682 286751 121685
rect 288574 121682 288634 122030
rect 289261 121954 289327 121957
rect 289261 121952 290076 121954
rect 289261 121896 289266 121952
rect 289322 121896 290076 121952
rect 289261 121894 290076 121896
rect 289261 121891 289327 121894
rect 286685 121680 288634 121682
rect 286685 121624 286690 121680
rect 286746 121624 288634 121680
rect 286685 121622 288634 121624
rect 286685 121619 286751 121622
rect 274541 121546 274607 121549
rect 275645 121546 275711 121549
rect 274541 121544 275711 121546
rect 274541 121488 274546 121544
rect 274602 121488 275650 121544
rect 275706 121488 275711 121544
rect 274541 121486 275711 121488
rect 274541 121483 274607 121486
rect 275645 121483 275711 121486
rect 288249 121546 288315 121549
rect 288249 121544 290076 121546
rect 288249 121488 288254 121544
rect 288310 121488 290076 121544
rect 288249 121486 290076 121488
rect 288249 121483 288315 121486
rect 249609 121410 249675 121413
rect 303797 121410 303863 121413
rect 249609 121408 252172 121410
rect 249609 121352 249614 121408
rect 249670 121352 252172 121408
rect 249609 121350 252172 121352
rect 301852 121408 303863 121410
rect 301852 121352 303802 121408
rect 303858 121352 303863 121408
rect 301852 121350 303863 121352
rect 249609 121347 249675 121350
rect 303797 121347 303863 121350
rect 269798 121274 269804 121276
rect 263948 121214 269804 121274
rect 269798 121212 269804 121214
rect 269868 121212 269874 121276
rect 288249 121138 288315 121141
rect 288249 121136 290076 121138
rect 288249 121080 288254 121136
rect 288310 121080 290076 121136
rect 288249 121078 290076 121080
rect 288249 121075 288315 121078
rect 65977 120866 66043 120869
rect 68142 120866 68816 120872
rect 65977 120864 68816 120866
rect 65977 120808 65982 120864
rect 66038 120812 68816 120864
rect 66038 120808 68202 120812
rect 65977 120806 68202 120808
rect 65977 120803 66043 120806
rect 209221 120730 209287 120733
rect 249241 120730 249307 120733
rect 209221 120728 249307 120730
rect 209221 120672 209226 120728
rect 209282 120672 249246 120728
rect 249302 120672 249307 120728
rect 209221 120670 249307 120672
rect 209221 120667 209287 120670
rect 249241 120667 249307 120670
rect 249701 120730 249767 120733
rect 266629 120730 266695 120733
rect 304942 120730 304948 120732
rect 249701 120728 252172 120730
rect 249701 120672 249706 120728
rect 249762 120672 252172 120728
rect 249701 120670 252172 120672
rect 263948 120728 266695 120730
rect 263948 120672 266634 120728
rect 266690 120672 266695 120728
rect 263948 120670 266695 120672
rect 249701 120667 249767 120670
rect 266629 120667 266695 120670
rect 277350 120670 290076 120730
rect 301852 120670 304948 120730
rect 265893 120594 265959 120597
rect 277350 120594 277410 120670
rect 304942 120668 304948 120670
rect 305012 120668 305018 120732
rect 265893 120592 277410 120594
rect 265893 120536 265898 120592
rect 265954 120536 277410 120592
rect 265893 120534 277410 120536
rect 265893 120531 265959 120534
rect 267089 120322 267155 120325
rect 263948 120320 267155 120322
rect 263948 120264 267094 120320
rect 267150 120264 267155 120320
rect 263948 120262 267155 120264
rect 267089 120259 267155 120262
rect 278998 120260 279004 120324
rect 279068 120322 279074 120324
rect 279068 120262 290076 120322
rect 279068 120260 279074 120262
rect 249701 120050 249767 120053
rect 278037 120050 278103 120053
rect 249701 120048 252172 120050
rect 249701 119992 249706 120048
rect 249762 119992 252172 120048
rect 249701 119990 252172 119992
rect 267690 120048 278103 120050
rect 267690 119992 278042 120048
rect 278098 119992 278103 120048
rect 267690 119990 278103 119992
rect 249701 119987 249767 119990
rect 267690 119778 267750 119990
rect 278037 119987 278103 119990
rect 263948 119718 267750 119778
rect 248781 119506 248847 119509
rect 248781 119504 252172 119506
rect 248781 119448 248786 119504
rect 248842 119448 252172 119504
rect 248781 119446 252172 119448
rect 248781 119443 248847 119446
rect 282310 119444 282316 119508
rect 282380 119506 282386 119508
rect 290046 119506 290106 119748
rect 282380 119446 290106 119506
rect 282380 119444 282386 119446
rect 224769 119370 224835 119373
rect 246389 119370 246455 119373
rect 266537 119370 266603 119373
rect 224769 119368 246455 119370
rect 224769 119312 224774 119368
rect 224830 119312 246394 119368
rect 246450 119312 246455 119368
rect 224769 119310 246455 119312
rect 263948 119368 266603 119370
rect 263948 119312 266542 119368
rect 266598 119312 266603 119368
rect 263948 119310 266603 119312
rect 224769 119307 224835 119310
rect 246389 119307 246455 119310
rect 266537 119307 266603 119310
rect 287605 119370 287671 119373
rect 301822 119370 301882 119884
rect 315941 119370 316007 119373
rect 287605 119368 290076 119370
rect 287605 119312 287610 119368
rect 287666 119312 290076 119368
rect 287605 119310 290076 119312
rect 301822 119368 316007 119370
rect 301822 119312 315946 119368
rect 316002 119312 316007 119368
rect 301822 119310 316007 119312
rect 287605 119307 287671 119310
rect 315941 119307 316007 119310
rect 303797 119234 303863 119237
rect 301852 119232 303863 119234
rect 301852 119176 303802 119232
rect 303858 119176 303863 119232
rect 301852 119174 303863 119176
rect 303797 119171 303863 119174
rect 266353 118962 266419 118965
rect 263948 118960 266419 118962
rect 263948 118904 266358 118960
rect 266414 118904 266419 118960
rect 263948 118902 266419 118904
rect 266353 118899 266419 118902
rect 286961 118962 287027 118965
rect 286961 118960 290076 118962
rect 286961 118904 286966 118960
rect 287022 118904 290076 118960
rect 286961 118902 290076 118904
rect 286961 118899 287027 118902
rect 249609 118826 249675 118829
rect 249609 118824 252172 118826
rect 249609 118768 249614 118824
rect 249670 118768 252172 118824
rect 249609 118766 252172 118768
rect 249609 118763 249675 118766
rect 268377 118418 268443 118421
rect 263948 118416 268443 118418
rect 263948 118360 268382 118416
rect 268438 118360 268443 118416
rect 263948 118358 268443 118360
rect 268377 118355 268443 118358
rect 290046 118282 290106 118524
rect 303797 118418 303863 118421
rect 301852 118416 303863 118418
rect 301852 118360 303802 118416
rect 303858 118360 303863 118416
rect 301852 118358 303863 118360
rect 303797 118355 303863 118358
rect 287010 118222 290106 118282
rect 248781 118146 248847 118149
rect 266353 118146 266419 118149
rect 248781 118144 252172 118146
rect 248781 118088 248786 118144
rect 248842 118088 252172 118144
rect 248781 118086 252172 118088
rect 265390 118144 266419 118146
rect 265390 118088 266358 118144
rect 266414 118088 266419 118144
rect 265390 118086 266419 118088
rect 248781 118083 248847 118086
rect 265390 118010 265450 118086
rect 266353 118083 266419 118086
rect 267181 118146 267247 118149
rect 276790 118146 276796 118148
rect 267181 118144 276796 118146
rect 267181 118088 267186 118144
rect 267242 118088 276796 118144
rect 267181 118086 276796 118088
rect 267181 118083 267247 118086
rect 276790 118084 276796 118086
rect 276860 118084 276866 118148
rect 263948 117950 265450 118010
rect 266169 118010 266235 118013
rect 266302 118010 266308 118012
rect 266169 118008 266308 118010
rect 266169 117952 266174 118008
rect 266230 117952 266308 118008
rect 266169 117950 266308 117952
rect 266169 117947 266235 117950
rect 266302 117948 266308 117950
rect 266372 117948 266378 118012
rect 276238 117948 276244 118012
rect 276308 118010 276314 118012
rect 277301 118010 277367 118013
rect 276308 118008 277367 118010
rect 276308 117952 277306 118008
rect 277362 117952 277367 118008
rect 276308 117950 277367 117952
rect 276308 117948 276314 117950
rect 277301 117947 277367 117950
rect 273253 117876 273319 117877
rect 273253 117874 273300 117876
rect 273208 117872 273300 117874
rect 273208 117816 273258 117872
rect 273208 117814 273300 117816
rect 273253 117812 273300 117814
rect 273364 117812 273370 117876
rect 274030 117812 274036 117876
rect 274100 117874 274106 117876
rect 287010 117874 287070 118222
rect 290046 117874 290106 118116
rect 274100 117814 287070 117874
rect 288022 117814 290106 117874
rect 274100 117812 274106 117814
rect 273253 117811 273319 117812
rect 266537 117466 266603 117469
rect 238710 117406 252172 117466
rect 263948 117464 266603 117466
rect 263948 117408 266542 117464
rect 266598 117408 266603 117464
rect 263948 117406 266603 117408
rect 170489 117330 170555 117333
rect 238710 117330 238770 117406
rect 266537 117403 266603 117406
rect 276657 117466 276723 117469
rect 288022 117466 288082 117814
rect 288249 117738 288315 117741
rect 288249 117736 290076 117738
rect 288249 117680 288254 117736
rect 288310 117680 290076 117736
rect 288249 117678 290076 117680
rect 288249 117675 288315 117678
rect 303889 117602 303955 117605
rect 301852 117600 303955 117602
rect 301852 117544 303894 117600
rect 303950 117544 303955 117600
rect 301852 117542 303955 117544
rect 303889 117539 303955 117542
rect 276657 117464 288082 117466
rect 276657 117408 276662 117464
rect 276718 117408 288082 117464
rect 276657 117406 288082 117408
rect 276657 117403 276723 117406
rect 170489 117328 238770 117330
rect 170489 117272 170494 117328
rect 170550 117272 238770 117328
rect 170489 117270 238770 117272
rect 170489 117267 170555 117270
rect 283557 117194 283623 117197
rect 267690 117192 283623 117194
rect 267690 117136 283562 117192
rect 283618 117136 283623 117192
rect 267690 117134 283623 117136
rect 267690 117058 267750 117134
rect 283557 117131 283623 117134
rect 288157 117194 288223 117197
rect 288157 117192 290076 117194
rect 288157 117136 288162 117192
rect 288218 117136 290076 117192
rect 288157 117134 290076 117136
rect 288157 117131 288223 117134
rect 263948 116998 267750 117058
rect 248781 116786 248847 116789
rect 289721 116786 289787 116789
rect 248781 116784 252172 116786
rect 248781 116728 248786 116784
rect 248842 116728 252172 116784
rect 248781 116726 252172 116728
rect 289721 116784 290076 116786
rect 289721 116728 289726 116784
rect 289782 116728 290076 116784
rect 289721 116726 290076 116728
rect 248781 116723 248847 116726
rect 289721 116723 289787 116726
rect 266353 116514 266419 116517
rect 263948 116512 266419 116514
rect 263948 116456 266358 116512
rect 266414 116456 266419 116512
rect 263948 116454 266419 116456
rect 266353 116451 266419 116454
rect 267089 116514 267155 116517
rect 279785 116514 279851 116517
rect 267089 116512 279851 116514
rect 267089 116456 267094 116512
rect 267150 116456 279790 116512
rect 279846 116456 279851 116512
rect 267089 116454 279851 116456
rect 267089 116451 267155 116454
rect 279785 116451 279851 116454
rect 287421 116378 287487 116381
rect 287421 116376 290076 116378
rect 287421 116320 287426 116376
rect 287482 116320 290076 116376
rect 287421 116318 290076 116320
rect 287421 116315 287487 116318
rect 301822 116242 301882 116892
rect 310462 116242 310468 116244
rect 301822 116182 310468 116242
rect 310462 116180 310468 116182
rect 310532 116180 310538 116244
rect 266353 116106 266419 116109
rect 303797 116106 303863 116109
rect 238710 116046 252172 116106
rect 263948 116104 266419 116106
rect 263948 116048 266358 116104
rect 266414 116048 266419 116104
rect 263948 116046 266419 116048
rect 301852 116104 303863 116106
rect 301852 116048 303802 116104
rect 303858 116048 303863 116104
rect 301852 116046 303863 116048
rect 206369 115970 206435 115973
rect 238710 115970 238770 116046
rect 266353 116043 266419 116046
rect 303797 116043 303863 116046
rect 206369 115968 238770 115970
rect 206369 115912 206374 115968
rect 206430 115912 238770 115968
rect 206369 115910 238770 115912
rect 282177 115970 282243 115973
rect 282177 115968 290076 115970
rect 282177 115912 282182 115968
rect 282238 115912 290076 115968
rect 282177 115910 290076 115912
rect 206369 115907 206435 115910
rect 282177 115907 282243 115910
rect 271413 115834 271479 115837
rect 271638 115834 271644 115836
rect 271413 115832 271644 115834
rect 271413 115776 271418 115832
rect 271474 115776 271644 115832
rect 271413 115774 271644 115776
rect 271413 115771 271479 115774
rect 271638 115772 271644 115774
rect 271708 115772 271714 115836
rect 279417 115834 279483 115837
rect 286542 115834 286548 115836
rect 279417 115832 286548 115834
rect 279417 115776 279422 115832
rect 279478 115776 286548 115832
rect 279417 115774 286548 115776
rect 279417 115771 279483 115774
rect 286542 115772 286548 115774
rect 286612 115772 286618 115836
rect 266353 115562 266419 115565
rect 263948 115560 266419 115562
rect 263948 115504 266358 115560
rect 266414 115504 266419 115560
rect 263948 115502 266419 115504
rect 266353 115499 266419 115502
rect 247861 115018 247927 115021
rect 252142 115018 252202 115396
rect 290046 115290 290106 115532
rect 303613 115426 303679 115429
rect 301852 115424 303679 115426
rect 301852 115368 303618 115424
rect 303674 115368 303679 115424
rect 301852 115366 303679 115368
rect 303613 115363 303679 115366
rect 277350 115230 290106 115290
rect 266537 115154 266603 115157
rect 263948 115152 266603 115154
rect 263948 115096 266542 115152
rect 266598 115096 266603 115152
rect 263948 115094 266603 115096
rect 266537 115091 266603 115094
rect 247861 115016 252202 115018
rect 247861 114960 247866 115016
rect 247922 114960 252202 115016
rect 247861 114958 252202 114960
rect 266169 115018 266235 115021
rect 277025 115018 277091 115021
rect 266169 115016 277091 115018
rect 266169 114960 266174 115016
rect 266230 114960 277030 115016
rect 277086 114960 277091 115016
rect 266169 114958 277091 114960
rect 247861 114955 247927 114958
rect 266169 114955 266235 114958
rect 277025 114955 277091 114958
rect 249701 114882 249767 114885
rect 249701 114880 252172 114882
rect 249701 114824 249706 114880
rect 249762 114824 252172 114880
rect 249701 114822 252172 114824
rect 249701 114819 249767 114822
rect 271270 114820 271276 114884
rect 271340 114882 271346 114884
rect 277350 114882 277410 115230
rect 288065 115154 288131 115157
rect 288065 115152 290076 115154
rect 288065 115096 288070 115152
rect 288126 115096 290076 115152
rect 288065 115094 290076 115096
rect 288065 115091 288131 115094
rect 271340 114822 277410 114882
rect 271340 114820 271346 114822
rect 266261 114746 266327 114749
rect 269062 114746 269068 114748
rect 266261 114744 269068 114746
rect 266261 114688 266266 114744
rect 266322 114688 269068 114744
rect 266261 114686 269068 114688
rect 266261 114683 266327 114686
rect 269062 114684 269068 114686
rect 269132 114684 269138 114748
rect 266997 114610 267063 114613
rect 263948 114608 267063 114610
rect 263948 114552 267002 114608
rect 267058 114552 267063 114608
rect 263948 114550 267063 114552
rect 266997 114547 267063 114550
rect 288249 114610 288315 114613
rect 303797 114610 303863 114613
rect 288249 114608 290076 114610
rect 288249 114552 288254 114608
rect 288310 114552 290076 114608
rect 288249 114550 290076 114552
rect 301852 114608 303863 114610
rect 301852 114552 303802 114608
rect 303858 114552 303863 114608
rect 301852 114550 303863 114552
rect 288249 114547 288315 114550
rect 303797 114547 303863 114550
rect 286593 114474 286659 114477
rect 267690 114472 286659 114474
rect 267690 114416 286598 114472
rect 286654 114416 286659 114472
rect 267690 114414 286659 114416
rect 249609 114202 249675 114205
rect 267690 114202 267750 114414
rect 286593 114411 286659 114414
rect 249609 114200 252172 114202
rect 249609 114144 249614 114200
rect 249670 114144 252172 114200
rect 249609 114142 252172 114144
rect 263948 114142 267750 114202
rect 287973 114202 288039 114205
rect 287973 114200 290076 114202
rect 287973 114144 287978 114200
rect 288034 114144 290076 114200
rect 287973 114142 290076 114144
rect 249609 114139 249675 114142
rect 287973 114139 288039 114142
rect 264094 113732 264100 113796
rect 264164 113794 264170 113796
rect 273253 113794 273319 113797
rect 264164 113792 273319 113794
rect 264164 113736 273258 113792
rect 273314 113736 273319 113792
rect 264164 113734 273319 113736
rect 264164 113732 264170 113734
rect 273253 113731 273319 113734
rect 277025 113794 277091 113797
rect 283925 113794 283991 113797
rect 277025 113792 283991 113794
rect 277025 113736 277030 113792
rect 277086 113736 283930 113792
rect 283986 113736 283991 113792
rect 277025 113734 283991 113736
rect 277025 113731 277091 113734
rect 283925 113731 283991 113734
rect 287605 113794 287671 113797
rect 303797 113794 303863 113797
rect 287605 113792 290076 113794
rect 287605 113736 287610 113792
rect 287666 113736 290076 113792
rect 287605 113734 290076 113736
rect 301852 113792 303863 113794
rect 301852 113736 303802 113792
rect 303858 113736 303863 113792
rect 301852 113734 303863 113736
rect 287605 113731 287671 113734
rect 303797 113731 303863 113734
rect 266353 113658 266419 113661
rect 263948 113656 266419 113658
rect 263948 113600 266358 113656
rect 266414 113600 266419 113656
rect 263948 113598 266419 113600
rect 266353 113595 266419 113598
rect 249701 113522 249767 113525
rect 249701 113520 252172 113522
rect 249701 113464 249706 113520
rect 249762 113464 252172 113520
rect 249701 113462 252172 113464
rect 249701 113459 249767 113462
rect 281441 113386 281507 113389
rect 281441 113384 290076 113386
rect 281441 113328 281446 113384
rect 281502 113328 290076 113384
rect 281441 113326 290076 113328
rect 281441 113323 281507 113326
rect 266537 113250 266603 113253
rect 263948 113248 266603 113250
rect 263948 113192 266542 113248
rect 266598 113192 266603 113248
rect 263948 113190 266603 113192
rect 266537 113187 266603 113190
rect 286777 113250 286843 113253
rect 287830 113250 287836 113252
rect 286777 113248 287836 113250
rect 286777 113192 286782 113248
rect 286838 113192 287836 113248
rect 286777 113190 287836 113192
rect 286777 113187 286843 113190
rect 287830 113188 287836 113190
rect 287900 113188 287906 113252
rect 287881 113114 287947 113117
rect 290038 113114 290044 113116
rect 287881 113112 290044 113114
rect 287881 113056 287886 113112
rect 287942 113056 290044 113112
rect 287881 113054 290044 113056
rect 287881 113051 287947 113054
rect 290038 113052 290044 113054
rect 290108 113052 290114 113116
rect 303797 113114 303863 113117
rect 301852 113112 303863 113114
rect 301852 113056 303802 113112
rect 303858 113056 303863 113112
rect 301852 113054 303863 113056
rect 303797 113051 303863 113054
rect 249241 112842 249307 112845
rect 249241 112840 252172 112842
rect 249241 112784 249246 112840
rect 249302 112784 252172 112840
rect 249241 112782 252172 112784
rect 249241 112779 249307 112782
rect 266353 112706 266419 112709
rect 263948 112704 266419 112706
rect 263948 112648 266358 112704
rect 266414 112648 266419 112704
rect 263948 112646 266419 112648
rect 266353 112643 266419 112646
rect 284293 112706 284359 112709
rect 290046 112706 290106 112948
rect 582925 112842 582991 112845
rect 583520 112842 584960 112932
rect 582925 112840 584960 112842
rect 582925 112784 582930 112840
rect 582986 112784 584960 112840
rect 582925 112782 584960 112784
rect 582925 112779 582991 112782
rect 284293 112704 290106 112706
rect 284293 112648 284298 112704
rect 284354 112648 290106 112704
rect 583520 112692 584960 112782
rect 284293 112646 290106 112648
rect 284293 112643 284359 112646
rect 202321 112434 202387 112437
rect 247769 112434 247835 112437
rect 202321 112432 247835 112434
rect 202321 112376 202326 112432
rect 202382 112376 247774 112432
rect 247830 112376 247835 112432
rect 202321 112374 247835 112376
rect 202321 112371 202387 112374
rect 247769 112371 247835 112374
rect 266537 112298 266603 112301
rect 263948 112296 266603 112298
rect 263948 112240 266542 112296
rect 266598 112240 266603 112296
rect 263948 112238 266603 112240
rect 266537 112235 266603 112238
rect 248965 112162 249031 112165
rect 286501 112162 286567 112165
rect 290046 112162 290106 112540
rect 303705 112298 303771 112301
rect 301852 112296 303771 112298
rect 301852 112240 303710 112296
rect 303766 112240 303771 112296
rect 301852 112238 303771 112240
rect 303705 112235 303771 112238
rect 248965 112160 252172 112162
rect 248965 112104 248970 112160
rect 249026 112104 252172 112160
rect 248965 112102 252172 112104
rect 286501 112160 290106 112162
rect 286501 112104 286506 112160
rect 286562 112104 290106 112160
rect 286501 112102 290106 112104
rect 248965 112099 249031 112102
rect 286501 112099 286567 112102
rect 266537 112026 266603 112029
rect 268694 112026 268700 112028
rect 266537 112024 268700 112026
rect 266537 111968 266542 112024
rect 266598 111968 268700 112024
rect 266537 111966 268700 111968
rect 266537 111963 266603 111966
rect 268694 111964 268700 111966
rect 268764 111964 268770 112028
rect 285622 111964 285628 112028
rect 285692 112026 285698 112028
rect 286961 112026 287027 112029
rect 285692 112024 287027 112026
rect 285692 111968 286966 112024
rect 287022 111968 287027 112024
rect 285692 111966 287027 111968
rect 285692 111964 285698 111966
rect 286961 111963 287027 111966
rect 287094 111964 287100 112028
rect 287164 112026 287170 112028
rect 288341 112026 288407 112029
rect 287164 112024 288407 112026
rect 287164 111968 288346 112024
rect 288402 111968 288407 112024
rect 287164 111966 288407 111968
rect 287164 111964 287170 111966
rect 288341 111963 288407 111966
rect 288574 111966 290076 112026
rect 268561 111890 268627 111893
rect 288574 111890 288634 111966
rect 268561 111888 288634 111890
rect 268561 111832 268566 111888
rect 268622 111832 288634 111888
rect 268561 111830 288634 111832
rect 268561 111827 268627 111830
rect 168281 111754 168347 111757
rect 280654 111754 280660 111756
rect 164694 111752 168347 111754
rect 164694 111696 168286 111752
rect 168342 111696 168347 111752
rect 164694 111694 168347 111696
rect 263948 111694 280660 111754
rect 168281 111691 168347 111694
rect 280654 111692 280660 111694
rect 280724 111692 280730 111756
rect 287973 111618 288039 111621
rect 303797 111618 303863 111621
rect 287973 111616 290076 111618
rect 287973 111560 287978 111616
rect 288034 111560 290076 111616
rect 287973 111558 290076 111560
rect 301852 111616 303863 111618
rect 301852 111560 303802 111616
rect 303858 111560 303863 111616
rect 301852 111558 303863 111560
rect 287973 111555 288039 111558
rect 303797 111555 303863 111558
rect 249241 111482 249307 111485
rect 249241 111480 252172 111482
rect 249241 111424 249246 111480
rect 249302 111424 252172 111480
rect 249241 111422 252172 111424
rect 249241 111419 249307 111422
rect 267181 111346 267247 111349
rect 263948 111344 267247 111346
rect 263948 111288 267186 111344
rect 267242 111288 267247 111344
rect 263948 111286 267247 111288
rect 267181 111283 267247 111286
rect 288249 111210 288315 111213
rect 288249 111208 290076 111210
rect 288249 111152 288254 111208
rect 288310 111152 290076 111208
rect 288249 111150 290076 111152
rect 288249 111147 288315 111150
rect 168005 111074 168071 111077
rect 177389 111074 177455 111077
rect 168005 111072 177455 111074
rect 168005 111016 168010 111072
rect 168066 111016 177394 111072
rect 177450 111016 177455 111072
rect 168005 111014 177455 111016
rect 168005 111011 168071 111014
rect 177389 111011 177455 111014
rect 177573 111074 177639 111077
rect 240869 111074 240935 111077
rect 177573 111072 240935 111074
rect 177573 111016 177578 111072
rect 177634 111016 240874 111072
rect 240930 111016 240935 111072
rect 177573 111014 240935 111016
rect 177573 111011 177639 111014
rect 240869 111011 240935 111014
rect 272517 111074 272583 111077
rect 286685 111074 286751 111077
rect 272517 111072 286751 111074
rect 272517 111016 272522 111072
rect 272578 111016 286690 111072
rect 286746 111016 286751 111072
rect 272517 111014 286751 111016
rect 272517 111011 272583 111014
rect 286685 111011 286751 111014
rect 248965 110802 249031 110805
rect 266445 110802 266511 110805
rect 248965 110800 252172 110802
rect -960 110666 480 110756
rect 248965 110744 248970 110800
rect 249026 110744 252172 110800
rect 248965 110742 252172 110744
rect 263948 110800 266511 110802
rect 263948 110744 266450 110800
rect 266506 110744 266511 110800
rect 263948 110742 266511 110744
rect 248965 110739 249031 110742
rect 266445 110739 266511 110742
rect 275553 110802 275619 110805
rect 303705 110802 303771 110805
rect 275553 110800 290076 110802
rect 275553 110744 275558 110800
rect 275614 110744 290076 110800
rect 275553 110742 290076 110744
rect 301852 110800 303771 110802
rect 301852 110744 303710 110800
rect 303766 110744 303771 110800
rect 301852 110742 303771 110744
rect 275553 110739 275619 110742
rect 303705 110739 303771 110742
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 267774 110468 267780 110532
rect 267844 110530 267850 110532
rect 268929 110530 268995 110533
rect 267844 110528 268995 110530
rect 267844 110472 268934 110528
rect 268990 110472 268995 110528
rect 267844 110470 268995 110472
rect 267844 110468 267850 110470
rect 268929 110467 268995 110470
rect 167913 110394 167979 110397
rect 283649 110394 283715 110397
rect 164694 110392 167979 110394
rect 164694 110336 167918 110392
rect 167974 110336 167979 110392
rect 164694 110334 167979 110336
rect 263948 110392 283715 110394
rect 263948 110336 283654 110392
rect 283710 110336 283715 110392
rect 263948 110334 283715 110336
rect 164694 110098 164754 110334
rect 167913 110331 167979 110334
rect 283649 110331 283715 110334
rect 288249 110394 288315 110397
rect 288249 110392 290076 110394
rect 288249 110336 288254 110392
rect 288310 110336 290076 110392
rect 288249 110334 290076 110336
rect 288249 110331 288315 110334
rect 249609 110258 249675 110261
rect 267273 110258 267339 110261
rect 268653 110258 268719 110261
rect 249609 110256 252172 110258
rect 249609 110200 249614 110256
rect 249670 110200 252172 110256
rect 249609 110198 252172 110200
rect 267273 110256 268719 110258
rect 267273 110200 267278 110256
rect 267334 110200 268658 110256
rect 268714 110200 268719 110256
rect 267273 110198 268719 110200
rect 249609 110195 249675 110198
rect 267273 110195 267339 110198
rect 268653 110195 268719 110198
rect 277350 109926 290076 109986
rect 266445 109850 266511 109853
rect 263948 109848 266511 109850
rect 263948 109792 266450 109848
rect 266506 109792 266511 109848
rect 263948 109790 266511 109792
rect 266445 109787 266511 109790
rect 273989 109850 274055 109853
rect 277350 109850 277410 109926
rect 273989 109848 277410 109850
rect 273989 109792 273994 109848
rect 274050 109792 277410 109848
rect 273989 109790 277410 109792
rect 273989 109787 274055 109790
rect 269614 109652 269620 109716
rect 269684 109714 269690 109716
rect 284293 109714 284359 109717
rect 269684 109712 284359 109714
rect 269684 109656 284298 109712
rect 284354 109656 284359 109712
rect 269684 109654 284359 109656
rect 269684 109652 269690 109654
rect 284293 109651 284359 109654
rect 249701 109578 249767 109581
rect 288341 109578 288407 109581
rect 249701 109576 252172 109578
rect 249701 109520 249706 109576
rect 249762 109520 252172 109576
rect 249701 109518 252172 109520
rect 288341 109576 290076 109578
rect 288341 109520 288346 109576
rect 288402 109520 290076 109576
rect 288341 109518 290076 109520
rect 249701 109515 249767 109518
rect 288341 109515 288407 109518
rect 266353 109442 266419 109445
rect 263948 109440 266419 109442
rect 263948 109384 266358 109440
rect 266414 109384 266419 109440
rect 263948 109382 266419 109384
rect 301822 109442 301882 109956
rect 309174 109442 309180 109444
rect 301822 109382 309180 109442
rect 266353 109379 266419 109382
rect 309174 109380 309180 109382
rect 309244 109380 309250 109444
rect 301852 109246 306390 109306
rect 270217 109170 270283 109173
rect 270350 109170 270356 109172
rect 270217 109168 270356 109170
rect 270217 109112 270222 109168
rect 270278 109112 270356 109168
rect 270217 109110 270356 109112
rect 270217 109107 270283 109110
rect 270350 109108 270356 109110
rect 270420 109108 270426 109172
rect 306330 109170 306390 109246
rect 312302 109170 312308 109172
rect 306330 109110 312308 109170
rect 312302 109108 312308 109110
rect 312372 109108 312378 109172
rect 167729 109034 167795 109037
rect 164694 109032 167795 109034
rect 164694 108976 167734 109032
rect 167790 108976 167795 109032
rect 164694 108974 167795 108976
rect 164694 108738 164754 108974
rect 167729 108971 167795 108974
rect 282453 109034 282519 109037
rect 287789 109034 287855 109037
rect 282453 109032 287855 109034
rect 282453 108976 282458 109032
rect 282514 108976 287794 109032
rect 287850 108976 287855 109032
rect 282453 108974 287855 108976
rect 282453 108971 282519 108974
rect 287789 108971 287855 108974
rect 249701 108898 249767 108901
rect 272558 108898 272564 108900
rect 249701 108896 252172 108898
rect 249701 108840 249706 108896
rect 249762 108840 252172 108896
rect 249701 108838 252172 108840
rect 263948 108838 272564 108898
rect 249701 108835 249767 108838
rect 272558 108836 272564 108838
rect 272628 108836 272634 108900
rect 286317 108762 286383 108765
rect 290046 108762 290106 109004
rect 286317 108760 290106 108762
rect 286317 108704 286322 108760
rect 286378 108704 290106 108760
rect 286317 108702 290106 108704
rect 286317 108699 286383 108702
rect 288341 108626 288407 108629
rect 288341 108624 290076 108626
rect 288341 108568 288346 108624
rect 288402 108568 290076 108624
rect 288341 108566 290076 108568
rect 288341 108563 288407 108566
rect 266353 108490 266419 108493
rect 304257 108490 304323 108493
rect 263948 108488 266419 108490
rect 263948 108432 266358 108488
rect 266414 108432 266419 108488
rect 263948 108430 266419 108432
rect 301852 108488 304323 108490
rect 301852 108432 304262 108488
rect 304318 108432 304323 108488
rect 301852 108430 304323 108432
rect 266353 108427 266419 108430
rect 304257 108427 304323 108430
rect 177389 108354 177455 108357
rect 249149 108354 249215 108357
rect 177389 108352 249215 108354
rect 177389 108296 177394 108352
rect 177450 108296 249154 108352
rect 249210 108296 249215 108352
rect 177389 108294 249215 108296
rect 177389 108291 177455 108294
rect 249149 108291 249215 108294
rect 249517 108218 249583 108221
rect 289077 108218 289143 108221
rect 249517 108216 252172 108218
rect 249517 108160 249522 108216
rect 249578 108160 252172 108216
rect 249517 108158 252172 108160
rect 289077 108216 290076 108218
rect 289077 108160 289082 108216
rect 289138 108160 290076 108216
rect 289077 108158 290076 108160
rect 249517 108155 249583 108158
rect 289077 108155 289143 108158
rect 266537 107946 266603 107949
rect 263948 107944 266603 107946
rect 263948 107888 266542 107944
rect 266598 107888 266603 107944
rect 263948 107886 266603 107888
rect 266537 107883 266603 107886
rect 303797 107810 303863 107813
rect 277350 107750 290076 107810
rect 301852 107808 303863 107810
rect 301852 107752 303802 107808
rect 303858 107752 303863 107808
rect 301852 107750 303863 107752
rect 271321 107674 271387 107677
rect 277350 107674 277410 107750
rect 303797 107747 303863 107750
rect 271321 107672 277410 107674
rect 271321 107616 271326 107672
rect 271382 107616 277410 107672
rect 271321 107614 277410 107616
rect 271321 107611 271387 107614
rect 249701 107538 249767 107541
rect 285070 107538 285076 107540
rect 249701 107536 252172 107538
rect 249701 107480 249706 107536
rect 249762 107480 252172 107536
rect 249701 107478 252172 107480
rect 263948 107478 285076 107538
rect 249701 107475 249767 107478
rect 285070 107476 285076 107478
rect 285140 107476 285146 107540
rect 287973 107402 288039 107405
rect 287973 107400 290076 107402
rect 287973 107344 287978 107400
rect 288034 107344 290076 107400
rect 287973 107342 290076 107344
rect 287973 107339 288039 107342
rect 266353 107130 266419 107133
rect 263948 107128 266419 107130
rect 263948 107072 266358 107128
rect 266414 107072 266419 107128
rect 263948 107070 266419 107072
rect 266353 107067 266419 107070
rect 288341 106994 288407 106997
rect 303797 106994 303863 106997
rect 288341 106992 290076 106994
rect 288341 106936 288346 106992
rect 288402 106936 290076 106992
rect 288341 106934 290076 106936
rect 301852 106992 303863 106994
rect 301852 106936 303802 106992
rect 303858 106936 303863 106992
rect 301852 106934 303863 106936
rect 288341 106931 288407 106934
rect 303797 106931 303863 106934
rect 249517 106858 249583 106861
rect 249517 106856 252172 106858
rect 249517 106800 249522 106856
rect 249578 106800 252172 106856
rect 249517 106798 252172 106800
rect 249517 106795 249583 106798
rect 266445 106586 266511 106589
rect 263948 106584 266511 106586
rect 263948 106528 266450 106584
rect 266506 106528 266511 106584
rect 263948 106526 266511 106528
rect 266445 106523 266511 106526
rect 277350 106390 290076 106450
rect 276841 106314 276907 106317
rect 277350 106314 277410 106390
rect 276841 106312 277410 106314
rect 276841 106256 276846 106312
rect 276902 106256 277410 106312
rect 276841 106254 277410 106256
rect 276841 106251 276907 106254
rect 248781 106178 248847 106181
rect 266302 106178 266308 106180
rect 248781 106176 252172 106178
rect 248781 106120 248786 106176
rect 248842 106120 252172 106176
rect 248781 106118 252172 106120
rect 263948 106118 266308 106178
rect 248781 106115 248847 106118
rect 266302 106116 266308 106118
rect 266372 106116 266378 106180
rect 280286 106116 280292 106180
rect 280356 106178 280362 106180
rect 281441 106178 281507 106181
rect 303654 106178 303660 106180
rect 280356 106176 281507 106178
rect 280356 106120 281446 106176
rect 281502 106120 281507 106176
rect 280356 106118 281507 106120
rect 301852 106118 303660 106178
rect 280356 106116 280362 106118
rect 281441 106115 281507 106118
rect 303654 106116 303660 106118
rect 303724 106116 303730 106180
rect 288341 106042 288407 106045
rect 288341 106040 290076 106042
rect 288341 105984 288346 106040
rect 288402 105984 290076 106040
rect 288341 105982 290076 105984
rect 288341 105979 288407 105982
rect 249701 105634 249767 105637
rect 266353 105634 266419 105637
rect 249701 105632 252172 105634
rect 249701 105576 249706 105632
rect 249762 105576 252172 105632
rect 249701 105574 252172 105576
rect 263948 105632 266419 105634
rect 263948 105576 266358 105632
rect 266414 105576 266419 105632
rect 263948 105574 266419 105576
rect 249701 105571 249767 105574
rect 266353 105571 266419 105574
rect 287973 105634 288039 105637
rect 287973 105632 290076 105634
rect 287973 105576 287978 105632
rect 288034 105576 290076 105632
rect 287973 105574 290076 105576
rect 287973 105571 288039 105574
rect 267038 105436 267044 105500
rect 267108 105498 267114 105500
rect 284017 105498 284083 105501
rect 303705 105498 303771 105501
rect 267108 105496 284083 105498
rect 267108 105440 284022 105496
rect 284078 105440 284083 105496
rect 267108 105438 284083 105440
rect 301852 105496 303771 105498
rect 301852 105440 303710 105496
rect 303766 105440 303771 105496
rect 301852 105438 303771 105440
rect 267108 105436 267114 105438
rect 284017 105435 284083 105438
rect 303705 105435 303771 105438
rect 264053 105362 264119 105365
rect 264053 105360 264162 105362
rect 264053 105304 264058 105360
rect 264114 105304 264162 105360
rect 264053 105299 264162 105304
rect 264102 105226 264162 105299
rect 263948 105166 264162 105226
rect 268377 105226 268443 105229
rect 268377 105224 290076 105226
rect 268377 105168 268382 105224
rect 268438 105168 290076 105224
rect 268377 105166 290076 105168
rect 268377 105163 268443 105166
rect 249609 104954 249675 104957
rect 249609 104952 252172 104954
rect 249609 104896 249614 104952
rect 249670 104896 252172 104952
rect 249609 104894 252172 104896
rect 249609 104891 249675 104894
rect 272558 104756 272564 104820
rect 272628 104818 272634 104820
rect 273161 104818 273227 104821
rect 272628 104816 273227 104818
rect 272628 104760 273166 104816
rect 273222 104760 273227 104816
rect 272628 104758 273227 104760
rect 272628 104756 272634 104758
rect 273161 104755 273227 104758
rect 268326 104682 268332 104684
rect 263948 104622 268332 104682
rect 268326 104620 268332 104622
rect 268396 104620 268402 104684
rect 290046 104546 290106 104788
rect 304349 104682 304415 104685
rect 301852 104680 304415 104682
rect 301852 104624 304354 104680
rect 304410 104624 304415 104680
rect 301852 104622 304415 104624
rect 304349 104619 304415 104622
rect 277350 104486 290106 104546
rect 203517 104274 203583 104277
rect 218697 104274 218763 104277
rect 203517 104272 218763 104274
rect 203517 104216 203522 104272
rect 203578 104216 218702 104272
rect 218758 104216 218763 104272
rect 203517 104214 218763 104216
rect 203517 104211 203583 104214
rect 218697 104211 218763 104214
rect 249701 104274 249767 104277
rect 271086 104274 271092 104276
rect 249701 104272 252172 104274
rect 249701 104216 249706 104272
rect 249762 104216 252172 104272
rect 249701 104214 252172 104216
rect 263948 104214 271092 104274
rect 249701 104211 249767 104214
rect 271086 104212 271092 104214
rect 271156 104212 271162 104276
rect 209129 104138 209195 104141
rect 249609 104138 249675 104141
rect 209129 104136 249675 104138
rect 209129 104080 209134 104136
rect 209190 104080 249614 104136
rect 249670 104080 249675 104136
rect 209129 104078 249675 104080
rect 209129 104075 209195 104078
rect 249609 104075 249675 104078
rect 274173 104002 274239 104005
rect 277350 104002 277410 104486
rect 274173 104000 277410 104002
rect 274173 103944 274178 104000
rect 274234 103944 277410 104000
rect 274173 103942 277410 103944
rect 288525 104002 288591 104005
rect 290046 104002 290106 104380
rect 303797 104002 303863 104005
rect 288525 104000 290106 104002
rect 288525 103944 288530 104000
rect 288586 103944 290106 104000
rect 288525 103942 290106 103944
rect 301852 104000 303863 104002
rect 301852 103944 303802 104000
rect 303858 103944 303863 104000
rect 301852 103942 303863 103944
rect 274173 103939 274239 103942
rect 288525 103939 288591 103942
rect 303797 103939 303863 103942
rect 270125 103866 270191 103869
rect 270125 103864 290076 103866
rect 270125 103808 270130 103864
rect 270186 103808 290076 103864
rect 270125 103806 290076 103808
rect 270125 103803 270191 103806
rect 266353 103730 266419 103733
rect 263948 103728 266419 103730
rect 263948 103672 266358 103728
rect 266414 103672 266419 103728
rect 263948 103670 266419 103672
rect 266353 103667 266419 103670
rect 248505 103594 248571 103597
rect 282269 103594 282335 103597
rect 288525 103594 288591 103597
rect 248505 103592 252172 103594
rect 248505 103536 248510 103592
rect 248566 103536 252172 103592
rect 248505 103534 252172 103536
rect 282269 103592 288591 103594
rect 282269 103536 282274 103592
rect 282330 103536 288530 103592
rect 288586 103536 288591 103592
rect 282269 103534 288591 103536
rect 248505 103531 248571 103534
rect 282269 103531 282335 103534
rect 288525 103531 288591 103534
rect 288341 103458 288407 103461
rect 288341 103456 290076 103458
rect 288341 103400 288346 103456
rect 288402 103400 290076 103456
rect 288341 103398 290076 103400
rect 288341 103395 288407 103398
rect 266353 103322 266419 103325
rect 263948 103320 266419 103322
rect 263948 103264 266358 103320
rect 266414 103264 266419 103320
rect 263948 103262 266419 103264
rect 266353 103259 266419 103262
rect 303613 103186 303679 103189
rect 301852 103184 303679 103186
rect 301852 103128 303618 103184
rect 303674 103128 303679 103184
rect 301852 103126 303679 103128
rect 303613 103123 303679 103126
rect 249701 102914 249767 102917
rect 249701 102912 252172 102914
rect 249701 102856 249706 102912
rect 249762 102856 252172 102912
rect 249701 102854 252172 102856
rect 249701 102851 249767 102854
rect 266445 102778 266511 102781
rect 290598 102780 290658 103020
rect 263948 102776 266511 102778
rect 263948 102720 266450 102776
rect 266506 102720 266511 102776
rect 263948 102718 266511 102720
rect 266445 102715 266511 102718
rect 290590 102716 290596 102780
rect 290660 102716 290666 102780
rect 288249 102642 288315 102645
rect 288249 102640 290076 102642
rect 288249 102584 288254 102640
rect 288310 102584 290076 102640
rect 288249 102582 290076 102584
rect 288249 102579 288315 102582
rect 268285 102506 268351 102509
rect 269062 102506 269068 102508
rect 268285 102504 269068 102506
rect 268285 102448 268290 102504
rect 268346 102448 269068 102504
rect 268285 102446 269068 102448
rect 268285 102443 268351 102446
rect 269062 102444 269068 102446
rect 269132 102444 269138 102508
rect 282913 102506 282979 102509
rect 287973 102506 288039 102509
rect 282913 102504 288039 102506
rect 282913 102448 282918 102504
rect 282974 102448 287978 102504
rect 288034 102448 288039 102504
rect 282913 102446 288039 102448
rect 282913 102443 282979 102446
rect 287973 102443 288039 102446
rect 67265 102370 67331 102373
rect 68142 102370 68816 102376
rect 265617 102370 265683 102373
rect 67265 102368 68816 102370
rect 67265 102312 67270 102368
rect 67326 102316 68816 102368
rect 263948 102368 265683 102370
rect 67326 102312 68202 102316
rect 67265 102310 68202 102312
rect 263948 102312 265622 102368
rect 265678 102312 265683 102368
rect 263948 102310 265683 102312
rect 67265 102307 67331 102310
rect 265617 102307 265683 102310
rect 269062 102308 269068 102372
rect 269132 102370 269138 102372
rect 270217 102370 270283 102373
rect 269132 102368 270283 102370
rect 269132 102312 270222 102368
rect 270278 102312 270283 102368
rect 269132 102310 270283 102312
rect 301852 102310 306390 102370
rect 269132 102308 269138 102310
rect 270217 102307 270283 102310
rect 249241 102234 249307 102237
rect 249241 102232 252172 102234
rect 249241 102176 249246 102232
rect 249302 102176 252172 102232
rect 249241 102174 252172 102176
rect 249241 102171 249307 102174
rect 267958 102172 267964 102236
rect 268028 102234 268034 102236
rect 269021 102234 269087 102237
rect 268028 102232 269087 102234
rect 268028 102176 269026 102232
rect 269082 102176 269087 102232
rect 268028 102174 269087 102176
rect 268028 102172 268034 102174
rect 269021 102171 269087 102174
rect 269849 102234 269915 102237
rect 306330 102234 306390 102310
rect 316166 102234 316172 102236
rect 269849 102232 290076 102234
rect 269849 102176 269854 102232
rect 269910 102176 290076 102232
rect 269849 102174 290076 102176
rect 306330 102174 316172 102234
rect 269849 102171 269915 102174
rect 316166 102172 316172 102174
rect 316236 102172 316242 102236
rect 266445 102098 266511 102101
rect 280838 102098 280844 102100
rect 266445 102096 280844 102098
rect 266445 102040 266450 102096
rect 266506 102040 280844 102096
rect 266445 102038 280844 102040
rect 266445 102035 266511 102038
rect 280838 102036 280844 102038
rect 280908 102036 280914 102100
rect 266353 101826 266419 101829
rect 263948 101824 266419 101826
rect 263948 101768 266358 101824
rect 266414 101768 266419 101824
rect 263948 101766 266419 101768
rect 266353 101763 266419 101766
rect 287605 101826 287671 101829
rect 287605 101824 290076 101826
rect 287605 101768 287610 101824
rect 287666 101768 290076 101824
rect 287605 101766 290076 101768
rect 287605 101763 287671 101766
rect 303705 101690 303771 101693
rect 301852 101688 303771 101690
rect 301852 101632 303710 101688
rect 303766 101632 303771 101688
rect 301852 101630 303771 101632
rect 303705 101627 303771 101630
rect 248781 101554 248847 101557
rect 267089 101554 267155 101557
rect 248781 101552 252172 101554
rect 248781 101496 248786 101552
rect 248842 101496 252172 101552
rect 248781 101494 252172 101496
rect 265206 101552 267155 101554
rect 265206 101496 267094 101552
rect 267150 101496 267155 101552
rect 265206 101494 267155 101496
rect 248781 101491 248847 101494
rect 169017 101418 169083 101421
rect 248505 101418 248571 101421
rect 265206 101418 265266 101494
rect 267089 101491 267155 101494
rect 169017 101416 248571 101418
rect 169017 101360 169022 101416
rect 169078 101360 248510 101416
rect 248566 101360 248571 101416
rect 169017 101358 248571 101360
rect 263948 101358 265266 101418
rect 266629 101418 266695 101421
rect 286174 101418 286180 101420
rect 266629 101416 286180 101418
rect 266629 101360 266634 101416
rect 266690 101360 286180 101416
rect 266629 101358 286180 101360
rect 169017 101355 169083 101358
rect 248505 101355 248571 101358
rect 266629 101355 266695 101358
rect 286174 101356 286180 101358
rect 286244 101356 286250 101420
rect 288341 101282 288407 101285
rect 288341 101280 290076 101282
rect 288341 101224 288346 101280
rect 288402 101224 290076 101280
rect 288341 101222 290076 101224
rect 288341 101219 288407 101222
rect 249149 101010 249215 101013
rect 271229 101010 271295 101013
rect 272558 101010 272564 101012
rect 249149 101008 252172 101010
rect 249149 100952 249154 101008
rect 249210 100952 252172 101008
rect 249149 100950 252172 100952
rect 271229 101008 272564 101010
rect 271229 100952 271234 101008
rect 271290 100952 272564 101008
rect 271229 100950 272564 100952
rect 249149 100947 249215 100950
rect 271229 100947 271295 100950
rect 272558 100948 272564 100950
rect 272628 100948 272634 101012
rect 284334 100948 284340 101012
rect 284404 101010 284410 101012
rect 285581 101010 285647 101013
rect 284404 101008 285647 101010
rect 284404 100952 285586 101008
rect 285642 100952 285647 101008
rect 284404 100950 285647 100952
rect 284404 100948 284410 100950
rect 285581 100947 285647 100950
rect 266445 100874 266511 100877
rect 263948 100872 266511 100874
rect 263948 100816 266450 100872
rect 266506 100816 266511 100872
rect 263948 100814 266511 100816
rect 266445 100811 266511 100814
rect 270534 100812 270540 100876
rect 270604 100874 270610 100876
rect 271413 100874 271479 100877
rect 270604 100872 271479 100874
rect 270604 100816 271418 100872
rect 271474 100816 271479 100872
rect 270604 100814 271479 100816
rect 270604 100812 270610 100814
rect 271413 100811 271479 100814
rect 272057 100874 272123 100877
rect 272057 100872 290076 100874
rect 272057 100816 272062 100872
rect 272118 100816 290076 100872
rect 272057 100814 290076 100816
rect 272057 100811 272123 100814
rect 67633 100738 67699 100741
rect 68142 100738 68816 100744
rect 67633 100736 68816 100738
rect 67633 100680 67638 100736
rect 67694 100684 68816 100736
rect 67694 100680 68202 100684
rect 67633 100678 68202 100680
rect 67633 100675 67699 100678
rect 301270 100605 301330 100844
rect 301270 100600 301379 100605
rect 301270 100544 301318 100600
rect 301374 100544 301379 100600
rect 301270 100542 301379 100544
rect 301313 100539 301379 100542
rect 266353 100466 266419 100469
rect 263948 100464 266419 100466
rect 263948 100408 266358 100464
rect 266414 100408 266419 100464
rect 263948 100406 266419 100408
rect 266353 100403 266419 100406
rect 288249 100466 288315 100469
rect 288249 100464 290076 100466
rect 288249 100408 288254 100464
rect 288310 100408 290076 100464
rect 288249 100406 290076 100408
rect 288249 100403 288315 100406
rect 249701 100330 249767 100333
rect 249701 100328 252172 100330
rect 249701 100272 249706 100328
rect 249762 100272 252172 100328
rect 249701 100270 252172 100272
rect 249701 100267 249767 100270
rect 266537 100058 266603 100061
rect 273846 100058 273852 100060
rect 266537 100056 273852 100058
rect 266537 100000 266542 100056
rect 266598 100000 273852 100056
rect 266537 99998 273852 100000
rect 266537 99995 266603 99998
rect 273846 99996 273852 99998
rect 273916 99996 273922 100060
rect 266445 99922 266511 99925
rect 263948 99920 266511 99922
rect 263948 99864 266450 99920
rect 266506 99864 266511 99920
rect 263948 99862 266511 99864
rect 266445 99859 266511 99862
rect 286174 99724 286180 99788
rect 286244 99786 286250 99788
rect 290046 99786 290106 100028
rect 286244 99726 290106 99786
rect 286244 99724 286250 99726
rect 301454 99653 301514 100164
rect 249517 99650 249583 99653
rect 288341 99650 288407 99653
rect 249517 99648 252172 99650
rect 249517 99592 249522 99648
rect 249578 99592 252172 99648
rect 249517 99590 252172 99592
rect 288341 99648 290076 99650
rect 288341 99592 288346 99648
rect 288402 99592 290076 99648
rect 288341 99590 290076 99592
rect 301454 99648 301563 99653
rect 301454 99592 301502 99648
rect 301558 99592 301563 99648
rect 301454 99590 301563 99592
rect 249517 99587 249583 99590
rect 288341 99587 288407 99590
rect 301497 99587 301563 99590
rect 266629 99514 266695 99517
rect 263948 99512 266695 99514
rect 263948 99456 266634 99512
rect 266690 99456 266695 99512
rect 263948 99454 266695 99456
rect 266629 99451 266695 99454
rect 583109 99514 583175 99517
rect 583520 99514 584960 99604
rect 583109 99512 584960 99514
rect 583109 99456 583114 99512
rect 583170 99456 584960 99512
rect 583109 99454 584960 99456
rect 583109 99451 583175 99454
rect 303613 99378 303679 99381
rect 301852 99376 303679 99378
rect 301852 99320 303618 99376
rect 303674 99320 303679 99376
rect 583520 99364 584960 99454
rect 301852 99318 303679 99320
rect 303613 99315 303679 99318
rect 264094 99044 264100 99108
rect 264164 99106 264170 99108
rect 264881 99106 264947 99109
rect 264164 99104 264947 99106
rect 264164 99048 264886 99104
rect 264942 99048 264947 99104
rect 264164 99046 264947 99048
rect 264164 99044 264170 99046
rect 264881 99043 264947 99046
rect 249609 98970 249675 98973
rect 265566 98970 265572 98972
rect 249609 98968 252172 98970
rect 249609 98912 249614 98968
rect 249670 98912 252172 98968
rect 249609 98910 252172 98912
rect 263948 98910 265572 98970
rect 249609 98907 249675 98910
rect 265566 98908 265572 98910
rect 265636 98908 265642 98972
rect 273846 98772 273852 98836
rect 273916 98834 273922 98836
rect 277025 98834 277091 98837
rect 273916 98832 277091 98834
rect 273916 98776 277030 98832
rect 277086 98776 277091 98832
rect 273916 98774 277091 98776
rect 273916 98772 273922 98774
rect 277025 98771 277091 98774
rect 288525 98834 288591 98837
rect 290046 98834 290106 99212
rect 288525 98832 290106 98834
rect 288525 98776 288530 98832
rect 288586 98776 290106 98832
rect 288525 98774 290106 98776
rect 288525 98771 288591 98774
rect 234061 98698 234127 98701
rect 250713 98698 250779 98701
rect 234061 98696 250779 98698
rect 234061 98640 234066 98696
rect 234122 98640 250718 98696
rect 250774 98640 250779 98696
rect 234061 98638 250779 98640
rect 234061 98635 234127 98638
rect 250713 98635 250779 98638
rect 266353 98698 266419 98701
rect 283782 98698 283788 98700
rect 266353 98696 283788 98698
rect 266353 98640 266358 98696
rect 266414 98640 283788 98696
rect 266353 98638 283788 98640
rect 266353 98635 266419 98638
rect 283782 98636 283788 98638
rect 283852 98636 283858 98700
rect 283925 98698 283991 98701
rect 283925 98696 290076 98698
rect 283925 98640 283930 98696
rect 283986 98640 290076 98696
rect 283925 98638 290076 98640
rect 283925 98635 283991 98638
rect 266537 98562 266603 98565
rect 302233 98562 302299 98565
rect 263948 98560 266603 98562
rect 263948 98504 266542 98560
rect 266598 98504 266603 98560
rect 263948 98502 266603 98504
rect 301852 98560 302299 98562
rect 301852 98504 302238 98560
rect 302294 98504 302299 98560
rect 301852 98502 302299 98504
rect 266537 98499 266603 98502
rect 302233 98499 302299 98502
rect 249701 98290 249767 98293
rect 282453 98290 282519 98293
rect 288525 98290 288591 98293
rect 249701 98288 252172 98290
rect 249701 98232 249706 98288
rect 249762 98232 252172 98288
rect 249701 98230 252172 98232
rect 282453 98288 288591 98290
rect 282453 98232 282458 98288
rect 282514 98232 288530 98288
rect 288586 98232 288591 98288
rect 282453 98230 288591 98232
rect 249701 98227 249767 98230
rect 282453 98227 282519 98230
rect 288525 98227 288591 98230
rect 266445 98018 266511 98021
rect 263948 98016 266511 98018
rect 263948 97960 266450 98016
rect 266506 97960 266511 98016
rect 263948 97958 266511 97960
rect 266445 97955 266511 97958
rect 283966 97956 283972 98020
rect 284036 98018 284042 98020
rect 284109 98018 284175 98021
rect 284036 98016 284175 98018
rect 284036 97960 284114 98016
rect 284170 97960 284175 98016
rect 284036 97958 284175 97960
rect 284036 97956 284042 97958
rect 284109 97955 284175 97958
rect 287789 98018 287855 98021
rect 290046 98018 290106 98260
rect 287789 98016 290106 98018
rect 287789 97960 287794 98016
rect 287850 97960 290106 98016
rect 287789 97958 290106 97960
rect 287789 97955 287855 97958
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 249701 97610 249767 97613
rect 266353 97610 266419 97613
rect 249701 97608 252172 97610
rect 249701 97552 249706 97608
rect 249762 97552 252172 97608
rect 249701 97550 252172 97552
rect 263948 97608 266419 97610
rect 263948 97552 266358 97608
rect 266414 97552 266419 97608
rect 263948 97550 266419 97552
rect 249701 97547 249767 97550
rect 266353 97547 266419 97550
rect 286593 97610 286659 97613
rect 290046 97610 290106 97852
rect 286593 97608 290106 97610
rect 286593 97552 286598 97608
rect 286654 97552 290106 97608
rect 286593 97550 290106 97552
rect 286593 97547 286659 97550
rect 287881 97474 287947 97477
rect 287881 97472 290076 97474
rect 287881 97416 287886 97472
rect 287942 97416 290076 97472
rect 287881 97414 290076 97416
rect 287881 97411 287947 97414
rect 301454 97341 301514 97852
rect 266905 97338 266971 97341
rect 276606 97338 276612 97340
rect 266905 97336 276612 97338
rect 266905 97280 266910 97336
rect 266966 97280 276612 97336
rect 266905 97278 276612 97280
rect 266905 97275 266971 97278
rect 276606 97276 276612 97278
rect 276676 97276 276682 97340
rect 301405 97336 301514 97341
rect 301405 97280 301410 97336
rect 301466 97280 301514 97336
rect 301405 97278 301514 97280
rect 301405 97275 301471 97278
rect 166206 97140 166212 97204
rect 166276 97202 166282 97204
rect 184381 97202 184447 97205
rect 166276 97200 184447 97202
rect 166276 97144 184386 97200
rect 184442 97144 184447 97200
rect 166276 97142 184447 97144
rect 166276 97140 166282 97142
rect 184381 97139 184447 97142
rect 196566 97140 196572 97204
rect 196636 97202 196642 97204
rect 252502 97202 252508 97204
rect 196636 97142 252508 97202
rect 196636 97140 196642 97142
rect 252502 97140 252508 97142
rect 252572 97140 252578 97204
rect 264329 97202 264395 97205
rect 276238 97202 276244 97204
rect 264329 97200 276244 97202
rect 264329 97144 264334 97200
rect 264390 97144 276244 97200
rect 264329 97142 276244 97144
rect 264329 97139 264395 97142
rect 276238 97140 276244 97142
rect 276308 97140 276314 97204
rect 267641 97066 267707 97069
rect 263948 97064 267707 97066
rect 263948 97008 267646 97064
rect 267702 97008 267707 97064
rect 263948 97006 267707 97008
rect 267641 97003 267707 97006
rect 288341 97066 288407 97069
rect 288341 97064 290076 97066
rect 288341 97008 288346 97064
rect 288402 97008 290076 97064
rect 288341 97006 290076 97008
rect 288341 97003 288407 97006
rect 249241 96930 249307 96933
rect 249241 96928 252172 96930
rect 249241 96872 249246 96928
rect 249302 96872 252172 96928
rect 249241 96870 252172 96872
rect 249241 96867 249307 96870
rect 301270 96661 301330 97036
rect 264145 96658 264211 96661
rect 266905 96658 266971 96661
rect 263948 96656 266971 96658
rect 263948 96600 264150 96656
rect 264206 96600 266910 96656
rect 266966 96600 266971 96656
rect 263948 96598 266971 96600
rect 264145 96595 264211 96598
rect 266905 96595 266971 96598
rect 276790 96596 276796 96660
rect 276860 96658 276866 96660
rect 276860 96598 290076 96658
rect 301270 96656 301379 96661
rect 301270 96600 301318 96656
rect 301374 96600 301379 96656
rect 301270 96598 301379 96600
rect 276860 96596 276866 96598
rect 301313 96595 301379 96598
rect 270718 96460 270724 96524
rect 270788 96522 270794 96524
rect 271781 96522 271847 96525
rect 270788 96520 271847 96522
rect 270788 96464 271786 96520
rect 271842 96464 271847 96520
rect 270788 96462 271847 96464
rect 270788 96460 270794 96462
rect 271781 96459 271847 96462
rect 249333 96386 249399 96389
rect 303889 96386 303955 96389
rect 249333 96384 252172 96386
rect 249333 96328 249338 96384
rect 249394 96328 252172 96384
rect 249333 96326 252172 96328
rect 301852 96384 303955 96386
rect 301852 96328 303894 96384
rect 303950 96328 303955 96384
rect 301852 96326 303955 96328
rect 249333 96323 249399 96326
rect 303889 96323 303955 96326
rect 266445 96250 266511 96253
rect 263948 96248 266511 96250
rect 263948 96192 266450 96248
rect 266506 96192 266511 96248
rect 263948 96190 266511 96192
rect 266445 96187 266511 96190
rect 257889 95980 257955 95981
rect 261017 95980 261083 95981
rect 257838 95978 257844 95980
rect 257798 95918 257844 95978
rect 257908 95976 257955 95980
rect 260966 95978 260972 95980
rect 257950 95920 257955 95976
rect 257838 95916 257844 95918
rect 257908 95916 257955 95920
rect 260926 95918 260972 95978
rect 261036 95976 261083 95980
rect 261078 95920 261083 95976
rect 260966 95916 260972 95918
rect 261036 95916 261083 95920
rect 257889 95915 257955 95916
rect 261017 95915 261083 95916
rect 262857 95978 262923 95981
rect 270534 95978 270540 95980
rect 262857 95976 270540 95978
rect 262857 95920 262862 95976
rect 262918 95920 270540 95976
rect 262857 95918 270540 95920
rect 262857 95915 262923 95918
rect 270534 95916 270540 95918
rect 270604 95916 270610 95980
rect 199469 95842 199535 95845
rect 249517 95842 249583 95845
rect 199469 95840 249583 95842
rect 199469 95784 199474 95840
rect 199530 95784 249522 95840
rect 249578 95784 249583 95840
rect 199469 95782 249583 95784
rect 199469 95779 199535 95782
rect 249517 95779 249583 95782
rect 257797 95842 257863 95845
rect 259310 95842 259316 95844
rect 257797 95840 259316 95842
rect 257797 95784 257802 95840
rect 257858 95784 259316 95840
rect 257797 95782 259316 95784
rect 257797 95779 257863 95782
rect 259310 95780 259316 95782
rect 259380 95780 259386 95844
rect 263041 95842 263107 95845
rect 278998 95842 279004 95844
rect 263041 95840 279004 95842
rect 263041 95784 263046 95840
rect 263102 95784 279004 95840
rect 263041 95782 279004 95784
rect 263041 95779 263107 95782
rect 278998 95780 279004 95782
rect 279068 95780 279074 95844
rect 290598 95706 290658 96220
rect 291101 95706 291167 95709
rect 290598 95704 291167 95706
rect 290598 95648 291106 95704
rect 291162 95648 291167 95704
rect 290598 95646 291167 95648
rect 291101 95643 291167 95646
rect 67265 95162 67331 95165
rect 165521 95162 165587 95165
rect 67265 95160 165587 95162
rect 67265 95104 67270 95160
rect 67326 95104 165526 95160
rect 165582 95104 165587 95160
rect 67265 95102 165587 95104
rect 67265 95099 67331 95102
rect 165521 95099 165587 95102
rect 227478 95100 227484 95164
rect 227548 95162 227554 95164
rect 301313 95162 301379 95165
rect 227548 95160 301379 95162
rect 227548 95104 301318 95160
rect 301374 95104 301379 95160
rect 227548 95102 301379 95104
rect 227548 95100 227554 95102
rect 301313 95099 301379 95102
rect 113136 94964 113142 95028
rect 113206 95026 113212 95028
rect 114502 95026 114508 95028
rect 113206 94966 114508 95026
rect 113206 94964 113212 94966
rect 114502 94964 114508 94966
rect 114572 94964 114578 95028
rect 151302 94964 151308 95028
rect 151372 95026 151378 95028
rect 151760 95026 151766 95028
rect 151372 94966 151766 95026
rect 151372 94964 151378 94966
rect 151760 94964 151766 94966
rect 151830 94964 151836 95028
rect 246297 95026 246363 95029
rect 301405 95026 301471 95029
rect 246297 95024 301471 95026
rect 246297 94968 246302 95024
rect 246358 94968 301410 95024
rect 301466 94968 301471 95024
rect 246297 94966 301471 94968
rect 246297 94963 246363 94966
rect 301405 94963 301471 94966
rect 289813 94892 289879 94893
rect 289813 94890 289860 94892
rect 289768 94888 289860 94890
rect 289768 94832 289818 94888
rect 289768 94830 289860 94832
rect 289813 94828 289860 94830
rect 289924 94828 289930 94892
rect 289813 94827 289879 94828
rect 124029 94756 124095 94757
rect 124016 94692 124022 94756
rect 124086 94754 124095 94756
rect 124086 94752 124178 94754
rect 124090 94696 124178 94752
rect 124086 94694 124178 94696
rect 124086 94692 124095 94694
rect 124029 94691 124095 94692
rect 262949 94482 263015 94485
rect 284293 94482 284359 94485
rect 262949 94480 284359 94482
rect 262949 94424 262954 94480
rect 263010 94424 284298 94480
rect 284354 94424 284359 94480
rect 262949 94422 284359 94424
rect 262949 94419 263015 94422
rect 284293 94419 284359 94422
rect 131982 94012 131988 94076
rect 132052 94074 132058 94076
rect 175917 94074 175983 94077
rect 132052 94072 175983 94074
rect 132052 94016 175922 94072
rect 175978 94016 175983 94072
rect 132052 94014 175983 94016
rect 132052 94012 132058 94014
rect 175917 94011 175983 94014
rect 96654 93876 96660 93940
rect 96724 93938 96730 93940
rect 229737 93938 229803 93941
rect 96724 93936 229803 93938
rect 96724 93880 229742 93936
rect 229798 93880 229803 93936
rect 96724 93878 229803 93880
rect 96724 93876 96730 93878
rect 229737 93875 229803 93878
rect 99230 93740 99236 93804
rect 99300 93802 99306 93804
rect 250621 93802 250687 93805
rect 99300 93800 250687 93802
rect 99300 93744 250626 93800
rect 250682 93744 250687 93800
rect 99300 93742 250687 93744
rect 99300 93740 99306 93742
rect 250621 93739 250687 93742
rect 99598 93604 99604 93668
rect 99668 93666 99674 93668
rect 172053 93666 172119 93669
rect 99668 93664 172119 93666
rect 99668 93608 172058 93664
rect 172114 93608 172119 93664
rect 99668 93606 172119 93608
rect 99668 93604 99674 93606
rect 172053 93603 172119 93606
rect 205398 93604 205404 93668
rect 205468 93666 205474 93668
rect 302233 93666 302299 93669
rect 205468 93664 302299 93666
rect 205468 93608 302238 93664
rect 302294 93608 302299 93664
rect 205468 93606 302299 93608
rect 205468 93604 205474 93606
rect 302233 93603 302299 93606
rect 119705 93532 119771 93533
rect 121729 93532 121795 93533
rect 119654 93530 119660 93532
rect 119614 93470 119660 93530
rect 119724 93528 119771 93532
rect 121678 93530 121684 93532
rect 119766 93472 119771 93528
rect 119654 93468 119660 93470
rect 119724 93468 119771 93472
rect 121638 93470 121684 93530
rect 121748 93528 121795 93532
rect 267733 93530 267799 93533
rect 121790 93472 121795 93528
rect 121678 93468 121684 93470
rect 121748 93468 121795 93472
rect 119705 93467 119771 93468
rect 121729 93467 121795 93468
rect 238710 93528 267799 93530
rect 238710 93472 267738 93528
rect 267794 93472 267799 93528
rect 238710 93470 267799 93472
rect 110137 93260 110203 93261
rect 110086 93258 110092 93260
rect 110046 93198 110092 93258
rect 110156 93256 110203 93260
rect 110198 93200 110203 93256
rect 110086 93196 110092 93198
rect 110156 93196 110203 93200
rect 110137 93195 110203 93196
rect 158713 93122 158779 93125
rect 168649 93122 168715 93125
rect 158713 93120 168715 93122
rect 158713 93064 158718 93120
rect 158774 93064 168654 93120
rect 168710 93064 168715 93120
rect 158713 93062 168715 93064
rect 158713 93059 158779 93062
rect 168649 93059 168715 93062
rect 229829 93122 229895 93125
rect 238518 93122 238524 93124
rect 229829 93120 238524 93122
rect 229829 93064 229834 93120
rect 229890 93064 238524 93120
rect 229829 93062 238524 93064
rect 229829 93059 229895 93062
rect 238518 93060 238524 93062
rect 238588 93122 238594 93124
rect 238710 93122 238770 93470
rect 267733 93467 267799 93470
rect 238588 93062 238770 93122
rect 238588 93060 238594 93062
rect 86718 92380 86724 92444
rect 86788 92442 86794 92444
rect 86861 92442 86927 92445
rect 86788 92440 86927 92442
rect 86788 92384 86866 92440
rect 86922 92384 86927 92440
rect 86788 92382 86927 92384
rect 86788 92380 86794 92382
rect 86861 92379 86927 92382
rect 88926 92380 88932 92444
rect 88996 92442 89002 92444
rect 89069 92442 89135 92445
rect 88996 92440 89135 92442
rect 88996 92384 89074 92440
rect 89130 92384 89135 92440
rect 88996 92382 89135 92384
rect 88996 92380 89002 92382
rect 89069 92379 89135 92382
rect 109166 92380 109172 92444
rect 109236 92442 109242 92444
rect 109953 92442 110019 92445
rect 109236 92440 110019 92442
rect 109236 92384 109958 92440
rect 110014 92384 110019 92440
rect 109236 92382 110019 92384
rect 109236 92380 109242 92382
rect 109953 92379 110019 92382
rect 111190 92380 111196 92444
rect 111260 92442 111266 92444
rect 111609 92442 111675 92445
rect 111260 92440 111675 92442
rect 111260 92384 111614 92440
rect 111670 92384 111675 92440
rect 111260 92382 111675 92384
rect 111260 92380 111266 92382
rect 111609 92379 111675 92382
rect 114461 92444 114527 92445
rect 136081 92444 136147 92445
rect 151353 92444 151419 92445
rect 114461 92440 114508 92444
rect 114572 92442 114578 92444
rect 136030 92442 136036 92444
rect 114461 92384 114466 92440
rect 114461 92380 114508 92384
rect 114572 92382 114618 92442
rect 135990 92382 136036 92442
rect 136100 92440 136147 92444
rect 151302 92442 151308 92444
rect 136142 92384 136147 92440
rect 114572 92380 114578 92382
rect 136030 92380 136036 92382
rect 136100 92380 136147 92384
rect 151262 92382 151308 92442
rect 151372 92440 151419 92444
rect 151414 92384 151419 92440
rect 151302 92380 151308 92382
rect 151372 92380 151419 92384
rect 114461 92379 114527 92380
rect 136081 92379 136147 92380
rect 151353 92379 151419 92380
rect 126881 92306 126947 92309
rect 206277 92306 206343 92309
rect 126881 92304 206343 92306
rect 126881 92248 126886 92304
rect 126942 92248 206282 92304
rect 206338 92248 206343 92304
rect 126881 92246 206343 92248
rect 126881 92243 126947 92246
rect 206277 92243 206343 92246
rect 120206 92108 120212 92172
rect 120276 92170 120282 92172
rect 164969 92170 165035 92173
rect 120276 92168 165035 92170
rect 120276 92112 164974 92168
rect 165030 92112 165035 92168
rect 120276 92110 165035 92112
rect 120276 92108 120282 92110
rect 164969 92107 165035 92110
rect 130745 92036 130811 92037
rect 130694 92034 130700 92036
rect 130654 91974 130700 92034
rect 130764 92032 130811 92036
rect 130806 91976 130811 92032
rect 130694 91972 130700 91974
rect 130764 91972 130811 91976
rect 130745 91971 130811 91972
rect 105670 91836 105676 91900
rect 105740 91898 105746 91900
rect 126605 91898 126671 91901
rect 105740 91896 126671 91898
rect 105740 91840 126610 91896
rect 126666 91840 126671 91896
rect 105740 91838 126671 91840
rect 105740 91836 105746 91838
rect 126605 91835 126671 91838
rect 258809 91898 258875 91901
rect 282453 91898 282519 91901
rect 258809 91896 282519 91898
rect 258809 91840 258814 91896
rect 258870 91840 282458 91896
rect 282514 91840 282519 91896
rect 258809 91838 282519 91840
rect 258809 91835 258875 91838
rect 282453 91835 282519 91838
rect 84326 91700 84332 91764
rect 84396 91762 84402 91764
rect 105537 91762 105603 91765
rect 84396 91760 105603 91762
rect 84396 91704 105542 91760
rect 105598 91704 105603 91760
rect 84396 91702 105603 91704
rect 84396 91700 84402 91702
rect 105537 91699 105603 91702
rect 106406 91700 106412 91764
rect 106476 91762 106482 91764
rect 107469 91762 107535 91765
rect 114921 91764 114987 91765
rect 114870 91762 114876 91764
rect 106476 91760 107535 91762
rect 106476 91704 107474 91760
rect 107530 91704 107535 91760
rect 106476 91702 107535 91704
rect 114830 91702 114876 91762
rect 114940 91760 114987 91764
rect 114982 91704 114987 91760
rect 106476 91700 106482 91702
rect 107469 91699 107535 91702
rect 114870 91700 114876 91702
rect 114940 91700 114987 91704
rect 116710 91700 116716 91764
rect 116780 91762 116786 91764
rect 198089 91762 198155 91765
rect 299473 91762 299539 91765
rect 116780 91702 122850 91762
rect 116780 91700 116786 91702
rect 114921 91699 114987 91700
rect 106774 91564 106780 91628
rect 106844 91626 106850 91628
rect 117221 91626 117287 91629
rect 106844 91624 117287 91626
rect 106844 91568 117226 91624
rect 117282 91568 117287 91624
rect 106844 91566 117287 91568
rect 106844 91564 106850 91566
rect 117221 91563 117287 91566
rect 98494 91428 98500 91492
rect 98564 91490 98570 91492
rect 98729 91490 98795 91493
rect 98564 91488 98795 91490
rect 98564 91432 98734 91488
rect 98790 91432 98795 91488
rect 98564 91430 98795 91432
rect 98564 91428 98570 91430
rect 98729 91427 98795 91430
rect 101857 91490 101923 91493
rect 101990 91490 101996 91492
rect 101857 91488 101996 91490
rect 101857 91432 101862 91488
rect 101918 91432 101996 91488
rect 101857 91430 101996 91432
rect 101857 91427 101923 91430
rect 101990 91428 101996 91430
rect 102060 91428 102066 91492
rect 122790 91490 122850 91702
rect 198089 91760 299539 91762
rect 198089 91704 198094 91760
rect 198150 91704 299478 91760
rect 299534 91704 299539 91760
rect 198089 91702 299539 91704
rect 198089 91699 198155 91702
rect 299473 91699 299539 91702
rect 125726 91564 125732 91628
rect 125796 91626 125802 91628
rect 126881 91626 126947 91629
rect 125796 91624 126947 91626
rect 125796 91568 126886 91624
rect 126942 91568 126947 91624
rect 125796 91566 126947 91568
rect 125796 91564 125802 91566
rect 126881 91563 126947 91566
rect 245009 91490 245075 91493
rect 122790 91488 245075 91490
rect 122790 91432 245014 91488
rect 245070 91432 245075 91488
rect 122790 91430 245075 91432
rect 245009 91427 245075 91430
rect 93894 91292 93900 91356
rect 93964 91354 93970 91356
rect 95049 91354 95115 91357
rect 93964 91352 95115 91354
rect 93964 91296 95054 91352
rect 95110 91296 95115 91352
rect 93964 91294 95115 91296
rect 93964 91292 93970 91294
rect 95049 91291 95115 91294
rect 101806 91292 101812 91356
rect 101876 91354 101882 91356
rect 102041 91354 102107 91357
rect 101876 91352 102107 91354
rect 101876 91296 102046 91352
rect 102102 91296 102107 91352
rect 101876 91294 102107 91296
rect 101876 91292 101882 91294
rect 102041 91291 102107 91294
rect 107694 91292 107700 91356
rect 107764 91354 107770 91356
rect 108849 91354 108915 91357
rect 107764 91352 108915 91354
rect 107764 91296 108854 91352
rect 108910 91296 108915 91352
rect 107764 91294 108915 91296
rect 107764 91292 107770 91294
rect 108849 91291 108915 91294
rect 115422 91292 115428 91356
rect 115492 91354 115498 91356
rect 115749 91354 115815 91357
rect 115492 91352 115815 91354
rect 115492 91296 115754 91352
rect 115810 91296 115815 91352
rect 115492 91294 115815 91296
rect 115492 91292 115498 91294
rect 115749 91291 115815 91294
rect 117998 91292 118004 91356
rect 118068 91354 118074 91356
rect 118509 91354 118575 91357
rect 122833 91356 122899 91357
rect 125409 91356 125475 91357
rect 118068 91352 118575 91354
rect 118068 91296 118514 91352
rect 118570 91296 118575 91352
rect 118068 91294 118575 91296
rect 118068 91292 118074 91294
rect 118509 91291 118575 91294
rect 122782 91292 122788 91356
rect 122852 91354 122899 91356
rect 125358 91354 125364 91356
rect 122852 91352 122944 91354
rect 122894 91296 122944 91352
rect 122852 91294 122944 91296
rect 125318 91294 125364 91354
rect 125428 91352 125475 91356
rect 125470 91296 125475 91352
rect 122852 91292 122899 91294
rect 125358 91292 125364 91294
rect 125428 91292 125475 91296
rect 126462 91292 126468 91356
rect 126532 91354 126538 91356
rect 126697 91354 126763 91357
rect 126532 91352 126763 91354
rect 126532 91296 126702 91352
rect 126758 91296 126763 91352
rect 126532 91294 126763 91296
rect 126532 91292 126538 91294
rect 122833 91291 122899 91292
rect 125409 91291 125475 91292
rect 126697 91291 126763 91294
rect 151629 91356 151695 91357
rect 151629 91352 151676 91356
rect 151740 91354 151746 91356
rect 151629 91296 151634 91352
rect 151629 91292 151676 91296
rect 151740 91294 151786 91354
rect 151740 91292 151746 91294
rect 151629 91291 151695 91292
rect 74758 91156 74764 91220
rect 74828 91218 74834 91220
rect 75821 91218 75887 91221
rect 74828 91216 75887 91218
rect 74828 91160 75826 91216
rect 75882 91160 75887 91216
rect 74828 91158 75887 91160
rect 74828 91156 74834 91158
rect 75821 91155 75887 91158
rect 85798 91156 85804 91220
rect 85868 91218 85874 91220
rect 86769 91218 86835 91221
rect 85868 91216 86835 91218
rect 85868 91160 86774 91216
rect 86830 91160 86835 91216
rect 85868 91158 86835 91160
rect 85868 91156 85874 91158
rect 86769 91155 86835 91158
rect 88006 91156 88012 91220
rect 88076 91218 88082 91220
rect 88149 91218 88215 91221
rect 88076 91216 88215 91218
rect 88076 91160 88154 91216
rect 88210 91160 88215 91216
rect 88076 91158 88215 91160
rect 88076 91156 88082 91158
rect 88149 91155 88215 91158
rect 90214 91156 90220 91220
rect 90284 91218 90290 91220
rect 91001 91218 91067 91221
rect 90284 91216 91067 91218
rect 90284 91160 91006 91216
rect 91062 91160 91067 91216
rect 90284 91158 91067 91160
rect 90284 91156 90290 91158
rect 91001 91155 91067 91158
rect 91318 91156 91324 91220
rect 91388 91218 91394 91220
rect 91921 91218 91987 91221
rect 91388 91216 91987 91218
rect 91388 91160 91926 91216
rect 91982 91160 91987 91216
rect 91388 91158 91987 91160
rect 91388 91156 91394 91158
rect 91921 91155 91987 91158
rect 92606 91156 92612 91220
rect 92676 91218 92682 91220
rect 93209 91218 93275 91221
rect 92676 91216 93275 91218
rect 92676 91160 93214 91216
rect 93270 91160 93275 91216
rect 92676 91158 93275 91160
rect 92676 91156 92682 91158
rect 93209 91155 93275 91158
rect 94998 91156 95004 91220
rect 95068 91218 95074 91220
rect 95141 91218 95207 91221
rect 95068 91216 95207 91218
rect 95068 91160 95146 91216
rect 95202 91160 95207 91216
rect 95068 91158 95207 91160
rect 95068 91156 95074 91158
rect 95141 91155 95207 91158
rect 96286 91156 96292 91220
rect 96356 91218 96362 91220
rect 96521 91218 96587 91221
rect 96356 91216 96587 91218
rect 96356 91160 96526 91216
rect 96582 91160 96587 91216
rect 96356 91158 96587 91160
rect 96356 91156 96362 91158
rect 96521 91155 96587 91158
rect 97206 91156 97212 91220
rect 97276 91218 97282 91220
rect 97901 91218 97967 91221
rect 97276 91216 97967 91218
rect 97276 91160 97906 91216
rect 97962 91160 97967 91216
rect 97276 91158 97967 91160
rect 97276 91156 97282 91158
rect 97901 91155 97967 91158
rect 98126 91156 98132 91220
rect 98196 91218 98202 91220
rect 99189 91218 99255 91221
rect 98196 91216 99255 91218
rect 98196 91160 99194 91216
rect 99250 91160 99255 91216
rect 98196 91158 99255 91160
rect 98196 91156 98202 91158
rect 99189 91155 99255 91158
rect 100518 91156 100524 91220
rect 100588 91218 100594 91220
rect 100661 91218 100727 91221
rect 100588 91216 100727 91218
rect 100588 91160 100666 91216
rect 100722 91160 100727 91216
rect 100588 91158 100727 91160
rect 100588 91156 100594 91158
rect 100661 91155 100727 91158
rect 100886 91156 100892 91220
rect 100956 91218 100962 91220
rect 101949 91218 102015 91221
rect 102593 91220 102659 91221
rect 102542 91218 102548 91220
rect 100956 91216 102015 91218
rect 100956 91160 101954 91216
rect 102010 91160 102015 91216
rect 100956 91158 102015 91160
rect 102502 91158 102548 91218
rect 102612 91216 102659 91220
rect 102654 91160 102659 91216
rect 100956 91156 100962 91158
rect 101949 91155 102015 91158
rect 102542 91156 102548 91158
rect 102612 91156 102659 91160
rect 102726 91156 102732 91220
rect 102796 91218 102802 91220
rect 103421 91218 103487 91221
rect 104249 91220 104315 91221
rect 104198 91218 104204 91220
rect 102796 91216 103487 91218
rect 102796 91160 103426 91216
rect 103482 91160 103487 91216
rect 102796 91158 103487 91160
rect 104158 91158 104204 91218
rect 104268 91216 104315 91220
rect 104310 91160 104315 91216
rect 102796 91156 102802 91158
rect 102593 91155 102659 91156
rect 103421 91155 103487 91158
rect 104198 91156 104204 91158
rect 104268 91156 104315 91160
rect 104566 91156 104572 91220
rect 104636 91218 104642 91220
rect 104801 91218 104867 91221
rect 104636 91216 104867 91218
rect 104636 91160 104806 91216
rect 104862 91160 104867 91216
rect 104636 91158 104867 91160
rect 104636 91156 104642 91158
rect 104249 91155 104315 91156
rect 104801 91155 104867 91158
rect 105486 91156 105492 91220
rect 105556 91156 105562 91220
rect 108062 91156 108068 91220
rect 108132 91218 108138 91220
rect 108941 91218 109007 91221
rect 108132 91216 109007 91218
rect 108132 91160 108946 91216
rect 109002 91160 109007 91216
rect 108132 91158 109007 91160
rect 108132 91156 108138 91158
rect 105494 91082 105554 91156
rect 108941 91155 109007 91158
rect 109534 91156 109540 91220
rect 109604 91218 109610 91220
rect 110321 91218 110387 91221
rect 109604 91216 110387 91218
rect 109604 91160 110326 91216
rect 110382 91160 110387 91216
rect 109604 91158 110387 91160
rect 109604 91156 109610 91158
rect 110321 91155 110387 91158
rect 110638 91156 110644 91220
rect 110708 91218 110714 91220
rect 111149 91218 111215 91221
rect 110708 91216 111215 91218
rect 110708 91160 111154 91216
rect 111210 91160 111215 91216
rect 110708 91158 111215 91160
rect 110708 91156 110714 91158
rect 111149 91155 111215 91158
rect 111926 91156 111932 91220
rect 111996 91218 112002 91220
rect 112069 91218 112135 91221
rect 111996 91216 112135 91218
rect 111996 91160 112074 91216
rect 112130 91160 112135 91216
rect 111996 91158 112135 91160
rect 111996 91156 112002 91158
rect 112069 91155 112135 91158
rect 112294 91156 112300 91220
rect 112364 91218 112370 91220
rect 112989 91218 113055 91221
rect 112364 91216 113055 91218
rect 112364 91160 112994 91216
rect 113050 91160 113055 91216
rect 112364 91158 113055 91160
rect 112364 91156 112370 91158
rect 112989 91155 113055 91158
rect 113214 91156 113220 91220
rect 113284 91218 113290 91220
rect 113449 91218 113515 91221
rect 114277 91220 114343 91221
rect 115841 91220 115907 91221
rect 114277 91218 114324 91220
rect 113284 91216 113515 91218
rect 113284 91160 113454 91216
rect 113510 91160 113515 91216
rect 113284 91158 113515 91160
rect 114232 91216 114324 91218
rect 114232 91160 114282 91216
rect 114232 91158 114324 91160
rect 113284 91156 113290 91158
rect 113449 91155 113515 91158
rect 114277 91156 114324 91158
rect 114388 91156 114394 91220
rect 115790 91218 115796 91220
rect 115750 91158 115796 91218
rect 115860 91216 115907 91220
rect 115902 91160 115907 91216
rect 115790 91156 115796 91158
rect 115860 91156 115907 91160
rect 117078 91156 117084 91220
rect 117148 91218 117154 91220
rect 117221 91218 117287 91221
rect 117148 91216 117287 91218
rect 117148 91160 117226 91216
rect 117282 91160 117287 91216
rect 117148 91158 117287 91160
rect 117148 91156 117154 91158
rect 114277 91155 114343 91156
rect 115841 91155 115907 91156
rect 117221 91155 117287 91158
rect 118182 91156 118188 91220
rect 118252 91218 118258 91220
rect 118601 91218 118667 91221
rect 118252 91216 118667 91218
rect 118252 91160 118606 91216
rect 118662 91160 118667 91216
rect 118252 91158 118667 91160
rect 118252 91156 118258 91158
rect 118601 91155 118667 91158
rect 119286 91156 119292 91220
rect 119356 91218 119362 91220
rect 119981 91218 120047 91221
rect 119356 91216 120047 91218
rect 119356 91160 119986 91216
rect 120042 91160 120047 91216
rect 119356 91158 120047 91160
rect 119356 91156 119362 91158
rect 119981 91155 120047 91158
rect 120574 91156 120580 91220
rect 120644 91218 120650 91220
rect 121361 91218 121427 91221
rect 120644 91216 121427 91218
rect 120644 91160 121366 91216
rect 121422 91160 121427 91216
rect 120644 91158 121427 91160
rect 120644 91156 120650 91158
rect 121361 91155 121427 91158
rect 122046 91156 122052 91220
rect 122116 91218 122122 91220
rect 122741 91218 122807 91221
rect 122116 91216 122807 91218
rect 122116 91160 122746 91216
rect 122802 91160 122807 91216
rect 122116 91158 122807 91160
rect 122116 91156 122122 91158
rect 122741 91155 122807 91158
rect 123150 91156 123156 91220
rect 123220 91218 123226 91220
rect 124121 91218 124187 91221
rect 123220 91216 124187 91218
rect 123220 91160 124126 91216
rect 124182 91160 124187 91216
rect 123220 91158 124187 91160
rect 123220 91156 123226 91158
rect 124121 91155 124187 91158
rect 124438 91156 124444 91220
rect 124508 91218 124514 91220
rect 125501 91218 125567 91221
rect 124508 91216 125567 91218
rect 124508 91160 125506 91216
rect 125562 91160 125567 91216
rect 124508 91158 125567 91160
rect 124508 91156 124514 91158
rect 125501 91155 125567 91158
rect 126646 91156 126652 91220
rect 126716 91218 126722 91220
rect 126789 91218 126855 91221
rect 126716 91216 126855 91218
rect 126716 91160 126794 91216
rect 126850 91160 126855 91216
rect 126716 91158 126855 91160
rect 126716 91156 126722 91158
rect 126789 91155 126855 91158
rect 127566 91156 127572 91220
rect 127636 91218 127642 91220
rect 127985 91218 128051 91221
rect 127636 91216 128051 91218
rect 127636 91160 127990 91216
rect 128046 91160 128051 91216
rect 127636 91158 128051 91160
rect 127636 91156 127642 91158
rect 127985 91155 128051 91158
rect 129406 91156 129412 91220
rect 129476 91218 129482 91220
rect 129641 91218 129707 91221
rect 129476 91216 129707 91218
rect 129476 91160 129646 91216
rect 129702 91160 129707 91216
rect 129476 91158 129707 91160
rect 129476 91156 129482 91158
rect 129641 91155 129707 91158
rect 133086 91156 133092 91220
rect 133156 91218 133162 91220
rect 133781 91218 133847 91221
rect 134425 91220 134491 91221
rect 134374 91218 134380 91220
rect 133156 91216 133847 91218
rect 133156 91160 133786 91216
rect 133842 91160 133847 91216
rect 133156 91158 133847 91160
rect 134334 91158 134380 91218
rect 134444 91216 134491 91220
rect 134486 91160 134491 91216
rect 133156 91156 133162 91158
rect 133781 91155 133847 91158
rect 134374 91156 134380 91158
rect 134444 91156 134491 91160
rect 151486 91156 151492 91220
rect 151556 91218 151562 91220
rect 151721 91218 151787 91221
rect 151556 91216 151787 91218
rect 151556 91160 151726 91216
rect 151782 91160 151787 91216
rect 151556 91158 151787 91160
rect 151556 91156 151562 91158
rect 134425 91155 134491 91156
rect 151721 91155 151787 91158
rect 151854 91156 151860 91220
rect 151924 91218 151930 91220
rect 153101 91218 153167 91221
rect 151924 91216 153167 91218
rect 151924 91160 153106 91216
rect 153162 91160 153167 91216
rect 151924 91158 153167 91160
rect 151924 91156 151930 91158
rect 153101 91155 153167 91158
rect 238201 91082 238267 91085
rect 105494 91080 238267 91082
rect 105494 91024 238206 91080
rect 238262 91024 238267 91080
rect 105494 91022 238267 91024
rect 238201 91019 238267 91022
rect 254577 90538 254643 90541
rect 271505 90538 271571 90541
rect 254577 90536 271571 90538
rect 254577 90480 254582 90536
rect 254638 90480 271510 90536
rect 271566 90480 271571 90536
rect 254577 90478 271571 90480
rect 254577 90475 254643 90478
rect 271505 90475 271571 90478
rect 130745 90402 130811 90405
rect 151077 90402 151143 90405
rect 130745 90400 151143 90402
rect 130745 90344 130750 90400
rect 130806 90344 151082 90400
rect 151138 90344 151143 90400
rect 130745 90342 151143 90344
rect 130745 90339 130811 90342
rect 151077 90339 151143 90342
rect 163497 90402 163563 90405
rect 180333 90402 180399 90405
rect 163497 90400 180399 90402
rect 163497 90344 163502 90400
rect 163558 90344 180338 90400
rect 180394 90344 180399 90400
rect 163497 90342 180399 90344
rect 163497 90339 163563 90342
rect 180333 90339 180399 90342
rect 226977 90402 227043 90405
rect 304257 90402 304323 90405
rect 226977 90400 304323 90402
rect 226977 90344 226982 90400
rect 227038 90344 304262 90400
rect 304318 90344 304323 90400
rect 226977 90342 304323 90344
rect 226977 90339 227043 90342
rect 304257 90339 304323 90342
rect 114921 89722 114987 89725
rect 184289 89722 184355 89725
rect 114921 89720 184355 89722
rect 114921 89664 114926 89720
rect 114982 89664 184294 89720
rect 184350 89664 184355 89720
rect 114921 89662 184355 89664
rect 114921 89659 114987 89662
rect 184289 89659 184355 89662
rect 110137 89586 110203 89589
rect 170489 89586 170555 89589
rect 110137 89584 170555 89586
rect 110137 89528 110142 89584
rect 110198 89528 170494 89584
rect 170550 89528 170555 89584
rect 110137 89526 170555 89528
rect 110137 89523 110203 89526
rect 170489 89523 170555 89526
rect 249057 89178 249123 89181
rect 274030 89178 274036 89180
rect 249057 89176 274036 89178
rect 249057 89120 249062 89176
rect 249118 89120 274036 89176
rect 249057 89118 274036 89120
rect 249057 89115 249123 89118
rect 274030 89116 274036 89118
rect 274100 89116 274106 89180
rect 162209 89042 162275 89045
rect 231209 89042 231275 89045
rect 162209 89040 231275 89042
rect 162209 88984 162214 89040
rect 162270 88984 231214 89040
rect 231270 88984 231275 89040
rect 162209 88982 231275 88984
rect 162209 88979 162275 88982
rect 231209 88979 231275 88982
rect 236637 89042 236703 89045
rect 298737 89042 298803 89045
rect 236637 89040 298803 89042
rect 236637 88984 236642 89040
rect 236698 88984 298742 89040
rect 298798 88984 298803 89040
rect 236637 88982 298803 88984
rect 236637 88979 236703 88982
rect 298737 88979 298803 88982
rect 91921 88226 91987 88229
rect 166349 88226 166415 88229
rect 91921 88224 166415 88226
rect 91921 88168 91926 88224
rect 91982 88168 166354 88224
rect 166410 88168 166415 88224
rect 91921 88166 166415 88168
rect 91921 88163 91987 88166
rect 166349 88163 166415 88166
rect 259310 88164 259316 88228
rect 259380 88226 259386 88228
rect 303654 88226 303660 88228
rect 259380 88166 303660 88226
rect 259380 88164 259386 88166
rect 303654 88164 303660 88166
rect 303724 88164 303730 88228
rect 111149 88090 111215 88093
rect 171777 88090 171843 88093
rect 111149 88088 171843 88090
rect 111149 88032 111154 88088
rect 111210 88032 171782 88088
rect 171838 88032 171843 88088
rect 111149 88030 171843 88032
rect 111149 88027 111215 88030
rect 171777 88027 171843 88030
rect 134425 87954 134491 87957
rect 167913 87954 167979 87957
rect 134425 87952 167979 87954
rect 134425 87896 134430 87952
rect 134486 87896 167918 87952
rect 167974 87896 167979 87952
rect 134425 87894 167979 87896
rect 134425 87891 134491 87894
rect 167913 87891 167979 87894
rect 236637 87682 236703 87685
rect 267774 87682 267780 87684
rect 236637 87680 267780 87682
rect 236637 87624 236642 87680
rect 236698 87624 267780 87680
rect 236637 87622 267780 87624
rect 236637 87619 236703 87622
rect 267774 87620 267780 87622
rect 267844 87620 267850 87684
rect 232589 87546 232655 87549
rect 280889 87546 280955 87549
rect 232589 87544 280955 87546
rect 232589 87488 232594 87544
rect 232650 87488 280894 87544
rect 280950 87488 280955 87544
rect 232589 87486 280955 87488
rect 232589 87483 232655 87486
rect 280889 87483 280955 87486
rect 101857 86866 101923 86869
rect 169109 86866 169175 86869
rect 101857 86864 169175 86866
rect 101857 86808 101862 86864
rect 101918 86808 169114 86864
rect 169170 86808 169175 86864
rect 101857 86806 169175 86808
rect 101857 86803 101923 86806
rect 169109 86803 169175 86806
rect 112069 86730 112135 86733
rect 164877 86730 164943 86733
rect 112069 86728 164943 86730
rect 112069 86672 112074 86728
rect 112130 86672 164882 86728
rect 164938 86672 164943 86728
rect 112069 86670 164943 86672
rect 112069 86667 112135 86670
rect 164877 86667 164943 86670
rect 126605 86594 126671 86597
rect 173249 86594 173315 86597
rect 126605 86592 173315 86594
rect 126605 86536 126610 86592
rect 126666 86536 173254 86592
rect 173310 86536 173315 86592
rect 126605 86534 173315 86536
rect 126605 86531 126671 86534
rect 173249 86531 173315 86534
rect 238109 86186 238175 86189
rect 267958 86186 267964 86188
rect 238109 86184 267964 86186
rect 238109 86128 238114 86184
rect 238170 86128 267964 86184
rect 238109 86126 267964 86128
rect 238109 86123 238175 86126
rect 267958 86124 267964 86126
rect 268028 86124 268034 86188
rect 268653 86186 268719 86189
rect 287881 86186 287947 86189
rect 268653 86184 287947 86186
rect 268653 86128 268658 86184
rect 268714 86128 287886 86184
rect 287942 86128 287947 86184
rect 268653 86126 287947 86128
rect 268653 86123 268719 86126
rect 287881 86123 287947 86126
rect 583293 86186 583359 86189
rect 583520 86186 584960 86276
rect 583293 86184 584960 86186
rect 583293 86128 583298 86184
rect 583354 86128 584960 86184
rect 583293 86126 584960 86128
rect 583293 86123 583359 86126
rect 583520 86036 584960 86126
rect 93209 85506 93275 85509
rect 191281 85506 191347 85509
rect 93209 85504 191347 85506
rect 93209 85448 93214 85504
rect 93270 85448 191286 85504
rect 191342 85448 191347 85504
rect 93209 85446 191347 85448
rect 93209 85443 93275 85446
rect 191281 85443 191347 85446
rect 106181 85370 106247 85373
rect 174721 85370 174787 85373
rect 106181 85368 174787 85370
rect 106181 85312 106186 85368
rect 106242 85312 174726 85368
rect 174782 85312 174787 85368
rect 106181 85310 174787 85312
rect 106181 85307 106247 85310
rect 174721 85307 174787 85310
rect 104249 85234 104315 85237
rect 167821 85234 167887 85237
rect 104249 85232 167887 85234
rect 104249 85176 104254 85232
rect 104310 85176 167826 85232
rect 167882 85176 167887 85232
rect 104249 85174 167887 85176
rect 104249 85171 104315 85174
rect 167821 85171 167887 85174
rect 196801 84826 196867 84829
rect 279693 84826 279759 84829
rect 196801 84824 279759 84826
rect -960 84690 480 84780
rect 196801 84768 196806 84824
rect 196862 84768 279698 84824
rect 279754 84768 279759 84824
rect 196801 84766 279759 84768
rect 196801 84763 196867 84766
rect 279693 84763 279759 84766
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 115749 84146 115815 84149
rect 203609 84146 203675 84149
rect 115749 84144 203675 84146
rect 115749 84088 115754 84144
rect 115810 84088 203614 84144
rect 203670 84088 203675 84144
rect 115749 84086 203675 84088
rect 115749 84083 115815 84086
rect 203609 84083 203675 84086
rect 122741 84010 122807 84013
rect 166206 84010 166212 84012
rect 122741 84008 166212 84010
rect 122741 83952 122746 84008
rect 122802 83952 166212 84008
rect 122741 83950 166212 83952
rect 122741 83947 122807 83950
rect 166206 83948 166212 83950
rect 166276 83948 166282 84012
rect 22001 83466 22067 83469
rect 283966 83466 283972 83468
rect 22001 83464 283972 83466
rect 22001 83408 22006 83464
rect 22062 83408 283972 83464
rect 22001 83406 283972 83408
rect 22001 83403 22067 83406
rect 283966 83404 283972 83406
rect 284036 83404 284042 83468
rect 111057 82786 111123 82789
rect 181529 82786 181595 82789
rect 111057 82784 181595 82786
rect 111057 82728 111062 82784
rect 111118 82728 181534 82784
rect 181590 82728 181595 82784
rect 111057 82726 181595 82728
rect 111057 82723 111123 82726
rect 181529 82723 181595 82726
rect 243629 82378 243695 82381
rect 270718 82378 270724 82380
rect 243629 82376 270724 82378
rect 243629 82320 243634 82376
rect 243690 82320 270724 82376
rect 243629 82318 270724 82320
rect 243629 82315 243695 82318
rect 270718 82316 270724 82318
rect 270788 82316 270794 82380
rect 122097 82242 122163 82245
rect 287697 82242 287763 82245
rect 122097 82240 287763 82242
rect 122097 82184 122102 82240
rect 122158 82184 287702 82240
rect 287758 82184 287763 82240
rect 122097 82182 287763 82184
rect 122097 82179 122163 82182
rect 287697 82179 287763 82182
rect 34421 82106 34487 82109
rect 284937 82106 285003 82109
rect 34421 82104 285003 82106
rect 34421 82048 34426 82104
rect 34482 82048 284942 82104
rect 284998 82048 285003 82104
rect 34421 82046 285003 82048
rect 34421 82043 34487 82046
rect 284937 82043 285003 82046
rect 67449 81426 67515 81429
rect 169017 81426 169083 81429
rect 67449 81424 169083 81426
rect 67449 81368 67454 81424
rect 67510 81368 169022 81424
rect 169078 81368 169083 81424
rect 67449 81366 169083 81368
rect 67449 81363 67515 81366
rect 169017 81363 169083 81366
rect 105537 81290 105603 81293
rect 177481 81290 177547 81293
rect 105537 81288 177547 81290
rect 105537 81232 105542 81288
rect 105598 81232 177486 81288
rect 177542 81232 177547 81288
rect 105537 81230 177547 81232
rect 105537 81227 105603 81230
rect 177481 81227 177547 81230
rect 245009 80882 245075 80885
rect 290590 80882 290596 80884
rect 245009 80880 290596 80882
rect 245009 80824 245014 80880
rect 245070 80824 290596 80880
rect 245009 80822 290596 80824
rect 245009 80819 245075 80822
rect 290590 80820 290596 80822
rect 290660 80820 290666 80884
rect 99281 80746 99347 80749
rect 286409 80746 286475 80749
rect 99281 80744 286475 80746
rect 99281 80688 99286 80744
rect 99342 80688 286414 80744
rect 286470 80688 286475 80744
rect 99281 80686 286475 80688
rect 99281 80683 99347 80686
rect 286409 80683 286475 80686
rect 99189 80066 99255 80069
rect 188521 80066 188587 80069
rect 99189 80064 188587 80066
rect 99189 80008 99194 80064
rect 99250 80008 188526 80064
rect 188582 80008 188587 80064
rect 99189 80006 188587 80008
rect 99189 80003 99255 80006
rect 188521 80003 188587 80006
rect 35801 79522 35867 79525
rect 271270 79522 271276 79524
rect 35801 79520 271276 79522
rect 35801 79464 35806 79520
rect 35862 79464 271276 79520
rect 35801 79462 271276 79464
rect 35801 79459 35867 79462
rect 271270 79460 271276 79462
rect 271340 79460 271346 79524
rect 50889 79386 50955 79389
rect 289169 79386 289235 79389
rect 50889 79384 289235 79386
rect 50889 79328 50894 79384
rect 50950 79328 289174 79384
rect 289230 79328 289235 79384
rect 50889 79326 289235 79328
rect 50889 79323 50955 79326
rect 289169 79323 289235 79326
rect 22737 78026 22803 78029
rect 287789 78026 287855 78029
rect 22737 78024 287855 78026
rect 22737 77968 22742 78024
rect 22798 77968 287794 78024
rect 287850 77968 287855 78024
rect 22737 77966 287855 77968
rect 22737 77963 22803 77966
rect 287789 77963 287855 77966
rect 16481 77890 16547 77893
rect 286593 77890 286659 77893
rect 16481 77888 286659 77890
rect 16481 77832 16486 77888
rect 16542 77832 286598 77888
rect 286654 77832 286659 77888
rect 16481 77830 286659 77832
rect 16481 77827 16547 77830
rect 286593 77827 286659 77830
rect 151077 76802 151143 76805
rect 289813 76802 289879 76805
rect 151077 76800 289879 76802
rect 151077 76744 151082 76800
rect 151138 76744 289818 76800
rect 289874 76744 289879 76800
rect 151077 76742 289879 76744
rect 151077 76739 151143 76742
rect 289813 76739 289879 76742
rect 70209 76666 70275 76669
rect 282310 76666 282316 76668
rect 70209 76664 282316 76666
rect 70209 76608 70214 76664
rect 70270 76608 282316 76664
rect 70209 76606 282316 76608
rect 70209 76603 70275 76606
rect 282310 76604 282316 76606
rect 282380 76604 282386 76668
rect 4061 76530 4127 76533
rect 276790 76530 276796 76532
rect 4061 76528 276796 76530
rect 4061 76472 4066 76528
rect 4122 76472 276796 76528
rect 4061 76470 276796 76472
rect 4061 76467 4127 76470
rect 276790 76468 276796 76470
rect 276860 76468 276866 76532
rect 59169 75306 59235 75309
rect 249793 75306 249859 75309
rect 59169 75304 249859 75306
rect 59169 75248 59174 75304
rect 59230 75248 249798 75304
rect 249854 75248 249859 75304
rect 59169 75246 249859 75248
rect 59169 75243 59235 75246
rect 249793 75243 249859 75246
rect 88241 75170 88307 75173
rect 289261 75170 289327 75173
rect 88241 75168 289327 75170
rect 88241 75112 88246 75168
rect 88302 75112 289266 75168
rect 289322 75112 289327 75168
rect 88241 75110 289327 75112
rect 88241 75107 88307 75110
rect 289261 75107 289327 75110
rect 107009 74490 107075 74493
rect 171961 74490 172027 74493
rect 107009 74488 172027 74490
rect 107009 74432 107014 74488
rect 107070 74432 171966 74488
rect 172022 74432 172027 74488
rect 107009 74430 172027 74432
rect 107009 74427 107075 74430
rect 171961 74427 172027 74430
rect 100661 74354 100727 74357
rect 164969 74354 165035 74357
rect 100661 74352 165035 74354
rect 100661 74296 100666 74352
rect 100722 74296 164974 74352
rect 165030 74296 165035 74352
rect 100661 74294 165035 74296
rect 100661 74291 100727 74294
rect 164969 74291 165035 74294
rect 224217 74082 224283 74085
rect 269614 74082 269620 74084
rect 224217 74080 269620 74082
rect 224217 74024 224222 74080
rect 224278 74024 269620 74080
rect 224217 74022 269620 74024
rect 224217 74019 224283 74022
rect 269614 74020 269620 74022
rect 269684 74020 269690 74084
rect 214557 73946 214623 73949
rect 267038 73946 267044 73948
rect 214557 73944 267044 73946
rect 214557 73888 214562 73944
rect 214618 73888 267044 73944
rect 214557 73886 267044 73888
rect 214557 73883 214623 73886
rect 267038 73884 267044 73886
rect 267108 73884 267114 73948
rect 202229 73810 202295 73813
rect 299565 73810 299631 73813
rect 202229 73808 299631 73810
rect 202229 73752 202234 73808
rect 202290 73752 299570 73808
rect 299626 73752 299631 73808
rect 202229 73750 299631 73752
rect 202229 73747 202295 73750
rect 299565 73747 299631 73750
rect 582557 72994 582623 72997
rect 583520 72994 584960 73084
rect 582557 72992 584960 72994
rect 582557 72936 582562 72992
rect 582618 72936 584960 72992
rect 582557 72934 584960 72936
rect 582557 72931 582623 72934
rect 583520 72844 584960 72934
rect 95141 72586 95207 72589
rect 265709 72586 265775 72589
rect 95141 72584 265775 72586
rect 95141 72528 95146 72584
rect 95202 72528 265714 72584
rect 265770 72528 265775 72584
rect 95141 72526 265775 72528
rect 95141 72523 95207 72526
rect 265709 72523 265775 72526
rect 53741 72450 53807 72453
rect 289813 72450 289879 72453
rect 53741 72448 289879 72450
rect 53741 72392 53746 72448
rect 53802 72392 289818 72448
rect 289874 72392 289879 72448
rect 53741 72390 289879 72392
rect 53741 72387 53807 72390
rect 289813 72387 289879 72390
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 56501 71226 56567 71229
rect 248413 71226 248479 71229
rect 56501 71224 248479 71226
rect 56501 71168 56506 71224
rect 56562 71168 248418 71224
rect 248474 71168 248479 71224
rect 56501 71166 248479 71168
rect 56501 71163 56567 71166
rect 248413 71163 248479 71166
rect 79961 71090 80027 71093
rect 285121 71090 285187 71093
rect 79961 71088 285187 71090
rect 79961 71032 79966 71088
rect 80022 71032 285126 71088
rect 285182 71032 285187 71088
rect 79961 71030 285187 71032
rect 79961 71027 80027 71030
rect 285121 71027 285187 71030
rect 62021 69730 62087 69733
rect 255313 69730 255379 69733
rect 62021 69728 255379 69730
rect 62021 69672 62026 69728
rect 62082 69672 255318 69728
rect 255374 69672 255379 69728
rect 62021 69670 255379 69672
rect 62021 69667 62087 69670
rect 255313 69667 255379 69670
rect 13721 69594 13787 69597
rect 280286 69594 280292 69596
rect 13721 69592 280292 69594
rect 13721 69536 13726 69592
rect 13782 69536 280292 69592
rect 13721 69534 280292 69536
rect 13721 69531 13787 69534
rect 280286 69532 280292 69534
rect 280356 69532 280362 69596
rect 64413 68370 64479 68373
rect 262213 68370 262279 68373
rect 64413 68368 262279 68370
rect 64413 68312 64418 68368
rect 64474 68312 262218 68368
rect 262274 68312 262279 68368
rect 64413 68310 262279 68312
rect 64413 68307 64479 68310
rect 262213 68307 262279 68310
rect 19241 68234 19307 68237
rect 275369 68234 275435 68237
rect 19241 68232 275435 68234
rect 19241 68176 19246 68232
rect 19302 68176 275374 68232
rect 275430 68176 275435 68232
rect 19241 68174 275435 68176
rect 19241 68171 19307 68174
rect 275369 68171 275435 68174
rect 147029 67010 147095 67013
rect 262949 67010 263015 67013
rect 147029 67008 263015 67010
rect 147029 66952 147034 67008
rect 147090 66952 262954 67008
rect 263010 66952 263015 67008
rect 147029 66950 263015 66952
rect 147029 66947 147095 66950
rect 262949 66947 263015 66950
rect 41321 66874 41387 66877
rect 284293 66874 284359 66877
rect 41321 66872 284359 66874
rect 41321 66816 41326 66872
rect 41382 66816 284298 66872
rect 284354 66816 284359 66872
rect 41321 66814 284359 66816
rect 41321 66811 41387 66814
rect 284293 66811 284359 66814
rect 67541 66194 67607 66197
rect 249149 66194 249215 66197
rect 67541 66192 249215 66194
rect 67541 66136 67546 66192
rect 67602 66136 249154 66192
rect 249210 66136 249215 66192
rect 67541 66134 249215 66136
rect 67541 66131 67607 66134
rect 249149 66131 249215 66134
rect 60641 65514 60707 65517
rect 311893 65514 311959 65517
rect 60641 65512 311959 65514
rect 60641 65456 60646 65512
rect 60702 65456 311898 65512
rect 311954 65456 311959 65512
rect 60641 65454 311959 65456
rect 60641 65451 60707 65454
rect 311893 65451 311959 65454
rect 116577 64290 116643 64293
rect 257337 64290 257403 64293
rect 116577 64288 257403 64290
rect 116577 64232 116582 64288
rect 116638 64232 257342 64288
rect 257398 64232 257403 64288
rect 116577 64230 257403 64232
rect 116577 64227 116643 64230
rect 257337 64227 257403 64230
rect 53741 64154 53807 64157
rect 289118 64154 289124 64156
rect 53741 64152 289124 64154
rect 53741 64096 53746 64152
rect 53802 64096 289124 64152
rect 53741 64094 289124 64096
rect 53741 64091 53807 64094
rect 289118 64092 289124 64094
rect 289188 64092 289194 64156
rect 255405 63610 255471 63613
rect 259494 63610 259500 63612
rect 255405 63608 259500 63610
rect 255405 63552 255410 63608
rect 255466 63552 259500 63608
rect 255405 63550 259500 63552
rect 255405 63547 255471 63550
rect 259494 63548 259500 63550
rect 259564 63548 259570 63612
rect 67633 63474 67699 63477
rect 249241 63474 249307 63477
rect 67633 63472 249307 63474
rect 67633 63416 67638 63472
rect 67694 63416 249246 63472
rect 249302 63416 249307 63472
rect 67633 63414 249307 63416
rect 67633 63411 67699 63414
rect 249241 63411 249307 63414
rect 48129 62794 48195 62797
rect 285029 62794 285095 62797
rect 48129 62792 285095 62794
rect 48129 62736 48134 62792
rect 48190 62736 285034 62792
rect 285090 62736 285095 62792
rect 48129 62734 285095 62736
rect 48129 62731 48195 62734
rect 285029 62731 285095 62734
rect 235993 61570 236059 61573
rect 255405 61570 255471 61573
rect 235993 61568 255471 61570
rect 235993 61512 235998 61568
rect 236054 61512 255410 61568
rect 255466 61512 255471 61568
rect 235993 61510 255471 61512
rect 235993 61507 236059 61510
rect 255405 61507 255471 61510
rect 78581 61434 78647 61437
rect 277894 61434 277900 61436
rect 78581 61432 277900 61434
rect 78581 61376 78586 61432
rect 78642 61376 277900 61432
rect 78581 61374 277900 61376
rect 78581 61371 78647 61374
rect 277894 61372 277900 61374
rect 277964 61372 277970 61436
rect 66161 60074 66227 60077
rect 281073 60074 281139 60077
rect 66161 60072 281139 60074
rect 66161 60016 66166 60072
rect 66222 60016 281078 60072
rect 281134 60016 281139 60072
rect 66161 60014 281139 60016
rect 66161 60011 66227 60014
rect 281073 60011 281139 60014
rect 26141 59938 26207 59941
rect 283925 59938 283991 59941
rect 26141 59936 283991 59938
rect 26141 59880 26146 59936
rect 26202 59880 283930 59936
rect 283986 59880 283991 59936
rect 26141 59878 283991 59880
rect 26141 59875 26207 59878
rect 283925 59875 283991 59878
rect 583017 59666 583083 59669
rect 583520 59666 584960 59756
rect 583017 59664 584960 59666
rect 583017 59608 583022 59664
rect 583078 59608 584960 59664
rect 583017 59606 584960 59608
rect 583017 59603 583083 59606
rect 583520 59516 584960 59606
rect 100661 58714 100727 58717
rect 282126 58714 282132 58716
rect 100661 58712 282132 58714
rect -960 58578 480 58668
rect 100661 58656 100666 58712
rect 100722 58656 282132 58712
rect 100661 58654 282132 58656
rect 100661 58651 100727 58654
rect 282126 58652 282132 58654
rect 282196 58652 282202 58716
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 73061 58578 73127 58581
rect 276841 58578 276907 58581
rect 73061 58576 276907 58578
rect 73061 58520 73066 58576
rect 73122 58520 276846 58576
rect 276902 58520 276907 58576
rect 73061 58518 276907 58520
rect 73061 58515 73127 58518
rect 276841 58515 276907 58518
rect 103421 57218 103487 57221
rect 266854 57218 266860 57220
rect 103421 57216 266860 57218
rect 103421 57160 103426 57216
rect 103482 57160 266860 57216
rect 103421 57158 266860 57160
rect 103421 57155 103487 57158
rect 266854 57156 266860 57158
rect 266924 57156 266930 57220
rect 33041 55994 33107 55997
rect 151077 55994 151143 55997
rect 33041 55992 151143 55994
rect 33041 55936 33046 55992
rect 33102 55936 151082 55992
rect 151138 55936 151143 55992
rect 33041 55934 151143 55936
rect 33041 55931 33107 55934
rect 151077 55931 151143 55934
rect 111701 55858 111767 55861
rect 279601 55858 279667 55861
rect 111701 55856 279667 55858
rect 111701 55800 111706 55856
rect 111762 55800 279606 55856
rect 279662 55800 279667 55856
rect 111701 55798 279667 55800
rect 111701 55795 111767 55798
rect 279601 55795 279667 55798
rect 59261 54498 59327 54501
rect 106917 54498 106983 54501
rect 59261 54496 106983 54498
rect 59261 54440 59266 54496
rect 59322 54440 106922 54496
rect 106978 54440 106983 54496
rect 59261 54438 106983 54440
rect 59261 54435 59327 54438
rect 106917 54435 106983 54438
rect 108297 54498 108363 54501
rect 287094 54498 287100 54500
rect 108297 54496 287100 54498
rect 108297 54440 108302 54496
rect 108358 54440 287100 54496
rect 108297 54438 287100 54440
rect 108297 54435 108363 54438
rect 287094 54436 287100 54438
rect 287164 54436 287170 54500
rect 15101 53138 15167 53141
rect 269062 53138 269068 53140
rect 15101 53136 269068 53138
rect 15101 53080 15106 53136
rect 15162 53080 269068 53136
rect 15101 53078 269068 53080
rect 15101 53075 15167 53078
rect 269062 53076 269068 53078
rect 269132 53076 269138 53140
rect 64781 51778 64847 51781
rect 265750 51778 265756 51780
rect 64781 51776 265756 51778
rect 64781 51720 64786 51776
rect 64842 51720 265756 51776
rect 64781 51718 265756 51720
rect 64781 51715 64847 51718
rect 265750 51716 265756 51718
rect 265820 51716 265826 51780
rect 62021 50282 62087 50285
rect 264094 50282 264100 50284
rect 62021 50280 264100 50282
rect 62021 50224 62026 50280
rect 62082 50224 264100 50280
rect 62021 50222 264100 50224
rect 62021 50219 62087 50222
rect 264094 50220 264100 50222
rect 264164 50220 264170 50284
rect 17861 48922 17927 48925
rect 286174 48922 286180 48924
rect 17861 48920 286180 48922
rect 17861 48864 17866 48920
rect 17922 48864 286180 48920
rect 17861 48862 286180 48864
rect 17861 48859 17927 48862
rect 286174 48860 286180 48862
rect 286244 48860 286250 48924
rect 61878 47500 61884 47564
rect 61948 47562 61954 47564
rect 324405 47562 324471 47565
rect 61948 47560 324471 47562
rect 61948 47504 324410 47560
rect 324466 47504 324471 47560
rect 61948 47502 324471 47504
rect 61948 47500 61954 47502
rect 324405 47499 324471 47502
rect 582833 46338 582899 46341
rect 583520 46338 584960 46428
rect 582833 46336 584960 46338
rect 582833 46280 582838 46336
rect 582894 46280 584960 46336
rect 582833 46278 584960 46280
rect 582833 46275 582899 46278
rect 38561 46202 38627 46205
rect 282177 46202 282243 46205
rect 38561 46200 282243 46202
rect 38561 46144 38566 46200
rect 38622 46144 282182 46200
rect 282238 46144 282243 46200
rect 583520 46188 584960 46278
rect 38561 46142 282243 46144
rect 38561 46139 38627 46142
rect 282177 46139 282243 46142
rect -960 45522 480 45612
rect 2773 45522 2839 45525
rect -960 45520 2839 45522
rect -960 45464 2778 45520
rect 2834 45464 2839 45520
rect -960 45462 2839 45464
rect -960 45372 480 45462
rect 2773 45459 2839 45462
rect 42701 44842 42767 44845
rect 284334 44842 284340 44844
rect 42701 44840 284340 44842
rect 42701 44784 42706 44840
rect 42762 44784 284340 44840
rect 42701 44782 284340 44784
rect 42701 44779 42767 44782
rect 284334 44780 284340 44782
rect 284404 44780 284410 44844
rect 193857 43482 193923 43485
rect 256693 43482 256759 43485
rect 193857 43480 256759 43482
rect 193857 43424 193862 43480
rect 193918 43424 256698 43480
rect 256754 43424 256759 43480
rect 193857 43422 256759 43424
rect 193857 43419 193923 43422
rect 256693 43419 256759 43422
rect 151077 40626 151143 40629
rect 243629 40626 243695 40629
rect 151077 40624 243695 40626
rect 151077 40568 151082 40624
rect 151138 40568 243634 40624
rect 243690 40568 243695 40624
rect 151077 40566 243695 40568
rect 151077 40563 151143 40566
rect 243629 40563 243695 40566
rect 33777 39266 33843 39269
rect 258809 39266 258875 39269
rect 33777 39264 258875 39266
rect 33777 39208 33782 39264
rect 33838 39208 258814 39264
rect 258870 39208 258875 39264
rect 33777 39206 258875 39208
rect 33777 39203 33843 39206
rect 258809 39203 258875 39206
rect 29637 37906 29703 37909
rect 287646 37906 287652 37908
rect 29637 37904 287652 37906
rect 29637 37848 29642 37904
rect 29698 37848 287652 37904
rect 29637 37846 287652 37848
rect 29637 37843 29703 37846
rect 287646 37844 287652 37846
rect 287716 37844 287722 37908
rect 57789 35186 57855 35189
rect 263910 35186 263916 35188
rect 57789 35184 263916 35186
rect 57789 35128 57794 35184
rect 57850 35128 263916 35184
rect 57789 35126 263916 35128
rect 57789 35123 57855 35126
rect 263910 35124 263916 35126
rect 263980 35124 263986 35188
rect 52361 33826 52427 33829
rect 307753 33826 307819 33829
rect 52361 33824 307819 33826
rect 52361 33768 52366 33824
rect 52422 33768 307758 33824
rect 307814 33768 307819 33824
rect 52361 33766 307819 33768
rect 52361 33763 52427 33766
rect 307753 33763 307819 33766
rect 582741 33146 582807 33149
rect 583520 33146 584960 33236
rect 582741 33144 584960 33146
rect 582741 33088 582746 33144
rect 582802 33088 584960 33144
rect 582741 33086 584960 33088
rect 582741 33083 582807 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 57881 32466 57947 32469
rect 236637 32466 236703 32469
rect 57881 32464 236703 32466
rect 57881 32408 57886 32464
rect 57942 32408 236642 32464
rect 236698 32408 236703 32464
rect 57881 32406 236703 32408
rect 57881 32403 57947 32406
rect 236637 32403 236703 32406
rect 28901 30970 28967 30973
rect 273897 30970 273963 30973
rect 28901 30968 273963 30970
rect 28901 30912 28906 30968
rect 28962 30912 273902 30968
rect 273958 30912 273963 30968
rect 28901 30910 273963 30912
rect 28901 30907 28967 30910
rect 273897 30907 273963 30910
rect 55121 29610 55187 29613
rect 310513 29610 310579 29613
rect 55121 29608 310579 29610
rect 55121 29552 55126 29608
rect 55182 29552 310518 29608
rect 310574 29552 310579 29608
rect 55121 29550 310579 29552
rect 55121 29547 55187 29550
rect 310513 29547 310579 29550
rect 104157 28250 104223 28253
rect 238109 28250 238175 28253
rect 104157 28248 238175 28250
rect 104157 28192 104162 28248
rect 104218 28192 238114 28248
rect 238170 28192 238175 28248
rect 104157 28190 238175 28192
rect 104157 28187 104223 28190
rect 238109 28187 238175 28190
rect 66110 26828 66116 26892
rect 66180 26890 66186 26892
rect 296713 26890 296779 26893
rect 66180 26888 296779 26890
rect 66180 26832 296718 26888
rect 296774 26832 296779 26888
rect 66180 26830 296779 26832
rect 66180 26828 66186 26830
rect 296713 26827 296779 26830
rect 43897 25530 43963 25533
rect 278773 25530 278839 25533
rect 43897 25528 278839 25530
rect 43897 25472 43902 25528
rect 43958 25472 278778 25528
rect 278834 25472 278839 25528
rect 43897 25470 278839 25472
rect 43897 25467 43963 25470
rect 278773 25467 278839 25470
rect 228449 24170 228515 24173
rect 285673 24170 285739 24173
rect 228449 24168 285739 24170
rect 228449 24112 228454 24168
rect 228510 24112 285678 24168
rect 285734 24112 285739 24168
rect 228449 24110 285739 24112
rect 228449 24107 228515 24110
rect 285673 24107 285739 24110
rect 46841 22674 46907 22677
rect 258717 22674 258783 22677
rect 46841 22672 258783 22674
rect 46841 22616 46846 22672
rect 46902 22616 258722 22672
rect 258778 22616 258783 22672
rect 46841 22614 258783 22616
rect 46841 22611 46907 22614
rect 258717 22611 258783 22614
rect 24761 21314 24827 21317
rect 273846 21314 273852 21316
rect 24761 21312 273852 21314
rect 24761 21256 24766 21312
rect 24822 21256 273852 21312
rect 24761 21254 273852 21256
rect 24761 21251 24827 21254
rect 273846 21252 273852 21254
rect 273916 21252 273922 21316
rect 67766 19892 67772 19956
rect 67836 19954 67842 19956
rect 276105 19954 276171 19957
rect 67836 19952 276171 19954
rect 67836 19896 276110 19952
rect 276166 19896 276171 19952
rect 67836 19894 276171 19896
rect 67836 19892 67842 19894
rect 276105 19891 276171 19894
rect 582465 19818 582531 19821
rect 583520 19818 584960 19908
rect 582465 19816 584960 19818
rect 582465 19760 582470 19816
rect 582526 19760 584960 19816
rect 582465 19758 584960 19760
rect 582465 19755 582531 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 6821 18594 6887 18597
rect 260966 18594 260972 18596
rect 6821 18592 260972 18594
rect 6821 18536 6826 18592
rect 6882 18536 260972 18592
rect 6821 18534 260972 18536
rect 6821 18531 6887 18534
rect 260966 18532 260972 18534
rect 261036 18532 261042 18596
rect 86769 17234 86835 17237
rect 284886 17234 284892 17236
rect 86769 17232 284892 17234
rect 86769 17176 86774 17232
rect 86830 17176 284892 17232
rect 86769 17174 284892 17176
rect 86769 17171 86835 17174
rect 284886 17172 284892 17174
rect 284956 17172 284962 17236
rect 105537 15874 105603 15877
rect 285622 15874 285628 15876
rect 105537 15872 285628 15874
rect 105537 15816 105542 15872
rect 105598 15816 285628 15872
rect 105537 15814 285628 15816
rect 105537 15811 105603 15814
rect 285622 15812 285628 15814
rect 285692 15812 285698 15876
rect 186814 14452 186820 14516
rect 186884 14514 186890 14516
rect 261753 14514 261819 14517
rect 186884 14512 261819 14514
rect 186884 14456 261758 14512
rect 261814 14456 261819 14512
rect 186884 14454 261819 14456
rect 186884 14452 186890 14454
rect 261753 14451 261819 14454
rect 195237 13154 195303 13157
rect 268377 13154 268443 13157
rect 195237 13152 268443 13154
rect 195237 13096 195242 13152
rect 195298 13096 268382 13152
rect 268438 13096 268443 13152
rect 195237 13094 268443 13096
rect 195237 13091 195303 13094
rect 268377 13091 268443 13094
rect 180057 13018 180123 13021
rect 292573 13018 292639 13021
rect 180057 13016 292639 13018
rect 180057 12960 180062 13016
rect 180118 12960 292578 13016
rect 292634 12960 292639 13016
rect 180057 12958 292639 12960
rect 180057 12955 180123 12958
rect 292573 12955 292639 12958
rect 220077 11658 220143 11661
rect 288985 11658 289051 11661
rect 220077 11656 289051 11658
rect 220077 11600 220082 11656
rect 220138 11600 288990 11656
rect 289046 11600 289051 11656
rect 220077 11598 289051 11600
rect 220077 11595 220143 11598
rect 288985 11595 289051 11598
rect 298093 11658 298159 11661
rect 317454 11658 317460 11660
rect 298093 11656 317460 11658
rect 298093 11600 298098 11656
rect 298154 11600 317460 11656
rect 298093 11598 317460 11600
rect 298093 11595 298159 11598
rect 317454 11596 317460 11598
rect 317524 11596 317530 11660
rect 132953 10298 133019 10301
rect 165654 10298 165660 10300
rect 132953 10296 165660 10298
rect 132953 10240 132958 10296
rect 133014 10240 165660 10296
rect 132953 10238 165660 10240
rect 132953 10235 133019 10238
rect 165654 10236 165660 10238
rect 165724 10236 165730 10300
rect 191046 10236 191052 10300
rect 191116 10298 191122 10300
rect 280797 10298 280863 10301
rect 191116 10296 280863 10298
rect 191116 10240 280802 10296
rect 280858 10240 280863 10296
rect 191116 10238 280863 10240
rect 191116 10236 191122 10238
rect 280797 10235 280863 10238
rect 170254 8876 170260 8940
rect 170324 8938 170330 8940
rect 310237 8938 310303 8941
rect 170324 8936 310303 8938
rect 170324 8880 310242 8936
rect 310298 8880 310303 8936
rect 170324 8878 310303 8880
rect 170324 8876 170330 8878
rect 310237 8875 310303 8878
rect 240225 7034 240291 7037
rect 313825 7034 313891 7037
rect 240225 7032 313891 7034
rect 240225 6976 240230 7032
rect 240286 6976 313830 7032
rect 313886 6976 313891 7032
rect 240225 6974 313891 6976
rect 240225 6971 240291 6974
rect 313825 6971 313891 6974
rect 582649 6626 582715 6629
rect 583520 6626 584960 6716
rect 582649 6624 584960 6626
rect -960 6490 480 6580
rect 582649 6568 582654 6624
rect 582710 6568 584960 6624
rect 582649 6566 584960 6568
rect 582649 6563 582715 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 177297 6218 177363 6221
rect 242893 6218 242959 6221
rect 177297 6216 242959 6218
rect 177297 6160 177302 6216
rect 177358 6160 242898 6216
rect 242954 6160 242959 6216
rect 177297 6158 242959 6160
rect 177297 6155 177363 6158
rect 242893 6155 242959 6158
rect 247677 6218 247743 6221
rect 254669 6218 254735 6221
rect 247677 6216 254735 6218
rect 247677 6160 247682 6216
rect 247738 6160 254674 6216
rect 254730 6160 254735 6216
rect 247677 6158 254735 6160
rect 247677 6155 247743 6158
rect 254669 6155 254735 6158
rect 136449 4858 136515 4861
rect 168414 4858 168420 4860
rect 136449 4856 168420 4858
rect 136449 4800 136454 4856
rect 136510 4800 168420 4856
rect 136449 4798 168420 4800
rect 136449 4795 136515 4798
rect 168414 4796 168420 4798
rect 168484 4796 168490 4860
rect 218697 4858 218763 4861
rect 266537 4858 266603 4861
rect 218697 4856 266603 4858
rect 218697 4800 218702 4856
rect 218758 4800 266542 4856
rect 266598 4800 266603 4856
rect 218697 4798 266603 4800
rect 218697 4795 218763 4798
rect 266537 4795 266603 4798
rect 322054 4796 322060 4860
rect 322124 4858 322130 4860
rect 329189 4858 329255 4861
rect 322124 4856 329255 4858
rect 322124 4800 329194 4856
rect 329250 4800 329255 4856
rect 322124 4798 329255 4800
rect 322124 4796 322130 4798
rect 329189 4795 329255 4798
rect 173157 4042 173223 4045
rect 240225 4042 240291 4045
rect 173157 4040 240291 4042
rect 173157 3984 173162 4040
rect 173218 3984 240230 4040
rect 240286 3984 240291 4040
rect 173157 3982 240291 3984
rect 173157 3979 173223 3982
rect 240225 3979 240291 3982
rect 277158 3980 277164 4044
rect 277228 4042 277234 4044
rect 278313 4042 278379 4045
rect 277228 4040 278379 4042
rect 277228 3984 278318 4040
rect 278374 3984 278379 4040
rect 277228 3982 278379 3984
rect 277228 3980 277234 3982
rect 278313 3979 278379 3982
rect 309726 3980 309732 4044
rect 309796 4042 309802 4044
rect 317321 4042 317387 4045
rect 309796 4040 317387 4042
rect 309796 3984 317326 4040
rect 317382 3984 317387 4040
rect 309796 3982 317387 3984
rect 309796 3980 309802 3982
rect 317321 3979 317387 3982
rect 82077 3634 82143 3637
rect 126237 3634 126303 3637
rect 82077 3632 126303 3634
rect 82077 3576 82082 3632
rect 82138 3576 126242 3632
rect 126298 3576 126303 3632
rect 82077 3574 126303 3576
rect 82077 3571 82143 3574
rect 126237 3571 126303 3574
rect 351637 3634 351703 3637
rect 358813 3634 358879 3637
rect 351637 3632 358879 3634
rect 351637 3576 351642 3632
rect 351698 3576 358818 3632
rect 358874 3576 358879 3632
rect 351637 3574 358879 3576
rect 351637 3571 351703 3574
rect 358813 3571 358879 3574
rect 121085 3498 121151 3501
rect 191097 3498 191163 3501
rect 121085 3496 191163 3498
rect 121085 3440 121090 3496
rect 121146 3440 191102 3496
rect 191158 3440 191163 3496
rect 121085 3438 191163 3440
rect 121085 3435 121151 3438
rect 191097 3435 191163 3438
rect 252502 3436 252508 3500
rect 252572 3498 252578 3500
rect 253473 3498 253539 3501
rect 252572 3496 253539 3498
rect 252572 3440 253478 3496
rect 253534 3440 253539 3496
rect 252572 3438 253539 3440
rect 252572 3436 252578 3438
rect 253473 3435 253539 3438
rect 288934 3436 288940 3500
rect 289004 3498 289010 3500
rect 294873 3498 294939 3501
rect 289004 3496 294939 3498
rect 289004 3440 294878 3496
rect 294934 3440 294939 3496
rect 289004 3438 294939 3440
rect 289004 3436 289010 3438
rect 294873 3435 294939 3438
rect 307937 3498 308003 3501
rect 313222 3498 313228 3500
rect 307937 3496 313228 3498
rect 307937 3440 307942 3496
rect 307998 3440 313228 3496
rect 307937 3438 313228 3440
rect 307937 3435 308003 3438
rect 313222 3436 313228 3438
rect 313292 3436 313298 3500
rect 320214 3436 320220 3500
rect 320284 3498 320290 3500
rect 320909 3498 320975 3501
rect 320284 3496 320975 3498
rect 320284 3440 320914 3496
rect 320970 3440 320975 3496
rect 320284 3438 320975 3440
rect 320284 3436 320290 3438
rect 320909 3435 320975 3438
rect 322105 3498 322171 3501
rect 322974 3498 322980 3500
rect 322105 3496 322980 3498
rect 322105 3440 322110 3496
rect 322166 3440 322980 3496
rect 322105 3438 322980 3440
rect 322105 3435 322171 3438
rect 322974 3436 322980 3438
rect 323044 3436 323050 3500
rect 348049 3498 348115 3501
rect 357433 3498 357499 3501
rect 348049 3496 357499 3498
rect 348049 3440 348054 3496
rect 348110 3440 357438 3496
rect 357494 3440 357499 3496
rect 348049 3438 357499 3440
rect 348049 3435 348115 3438
rect 357433 3435 357499 3438
rect 19425 3362 19491 3365
rect 108297 3362 108363 3365
rect 19425 3360 108363 3362
rect 19425 3304 19430 3360
rect 19486 3304 108302 3360
rect 108358 3304 108363 3360
rect 19425 3302 108363 3304
rect 19425 3299 19491 3302
rect 108297 3299 108363 3302
rect 125869 3362 125935 3365
rect 232497 3362 232563 3365
rect 125869 3360 232563 3362
rect 125869 3304 125874 3360
rect 125930 3304 232502 3360
rect 232558 3304 232563 3360
rect 125869 3302 232563 3304
rect 125869 3299 125935 3302
rect 232497 3299 232563 3302
rect 243537 3362 243603 3365
rect 258257 3362 258323 3365
rect 243537 3360 258323 3362
rect 243537 3304 243542 3360
rect 243598 3304 258262 3360
rect 258318 3304 258323 3360
rect 243537 3302 258323 3304
rect 243537 3299 243603 3302
rect 258257 3299 258323 3302
rect 271321 3362 271387 3365
rect 274817 3362 274883 3365
rect 271321 3360 274883 3362
rect 271321 3304 271326 3360
rect 271382 3304 274822 3360
rect 274878 3304 274883 3360
rect 271321 3302 274883 3304
rect 271321 3299 271387 3302
rect 274817 3299 274883 3302
rect 275134 3300 275140 3364
rect 275204 3362 275210 3364
rect 280705 3362 280771 3365
rect 275204 3360 280771 3362
rect 275204 3304 280710 3360
rect 280766 3304 280771 3360
rect 275204 3302 280771 3304
rect 275204 3300 275210 3302
rect 280705 3299 280771 3302
rect 344553 3362 344619 3365
rect 356053 3362 356119 3365
rect 344553 3360 356119 3362
rect 344553 3304 344558 3360
rect 344614 3304 356058 3360
rect 356114 3304 356119 3360
rect 344553 3302 356119 3304
rect 344553 3299 344619 3302
rect 356053 3299 356119 3302
rect 48221 2002 48287 2005
rect 318517 2002 318583 2005
rect 48221 2000 318583 2002
rect 48221 1944 48226 2000
rect 48282 1944 318522 2000
rect 318578 1944 318583 2000
rect 48221 1942 318583 1944
rect 48221 1939 48287 1942
rect 318517 1939 318583 1942
<< via3 >>
rect 69612 702476 69676 702540
rect 76052 699756 76116 699820
rect 88196 588508 88260 588572
rect 159220 586468 159284 586532
rect 88196 585652 88260 585716
rect 67772 583748 67836 583812
rect 69428 581844 69492 581908
rect 119476 580212 119540 580276
rect 111012 553420 111076 553484
rect 66668 550836 66732 550900
rect 99972 550700 100036 550764
rect 109356 546484 109420 546548
rect 76052 538052 76116 538116
rect 69612 535528 69676 535532
rect 69612 535472 69662 535528
rect 69662 535472 69676 535528
rect 69612 535468 69676 535472
rect 71820 535468 71884 535532
rect 122604 469780 122668 469844
rect 106412 467060 106476 467124
rect 96844 462844 96908 462908
rect 120212 462844 120276 462908
rect 89668 461484 89732 461548
rect 111748 461484 111812 461548
rect 92612 460124 92676 460188
rect 102732 460124 102796 460188
rect 104940 459580 105004 459644
rect 107700 458764 107764 458828
rect 67772 457404 67836 457468
rect 98132 457404 98196 457468
rect 91140 456180 91204 456244
rect 100708 456044 100772 456108
rect 115980 456044 116044 456108
rect 148180 455500 148244 455564
rect 121684 451828 121748 451892
rect 172468 449984 172532 449988
rect 172468 449928 172518 449984
rect 172518 449928 172532 449984
rect 172468 449924 172532 449928
rect 95188 449108 95252 449172
rect 160692 448564 160756 448628
rect 123340 447612 123404 447676
rect 96476 446388 96540 446452
rect 90220 445844 90284 445908
rect 95004 445708 95068 445772
rect 96660 445768 96724 445772
rect 96660 445712 96674 445768
rect 96674 445712 96724 445768
rect 96660 445708 96724 445712
rect 99052 445708 99116 445772
rect 110644 445708 110708 445772
rect 114324 445708 114388 445772
rect 118556 445708 118620 445772
rect 109172 444620 109236 444684
rect 119844 444620 119908 444684
rect 68876 444212 68940 444276
rect 123340 444212 123404 444276
rect 120028 442716 120092 442780
rect 143580 442308 143644 442372
rect 165660 441628 165724 441692
rect 122788 435236 122852 435300
rect 120396 434692 120460 434756
rect 120212 431428 120276 431492
rect 122604 425580 122668 425644
rect 66668 410484 66732 410548
rect 69244 408172 69308 408236
rect 121684 403684 121748 403748
rect 140820 401644 140884 401708
rect 61884 393272 61948 393276
rect 61884 393216 61934 393272
rect 61934 393216 61948 393272
rect 61884 393212 61948 393216
rect 113036 391988 113100 392052
rect 92612 390900 92676 390964
rect 102732 390900 102796 390964
rect 100708 390552 100772 390556
rect 100708 390496 100722 390552
rect 100722 390496 100772 390552
rect 100708 390492 100772 390496
rect 69612 390356 69676 390420
rect 71820 390416 71884 390420
rect 71820 390360 71870 390416
rect 71870 390360 71884 390416
rect 71820 390356 71884 390360
rect 89668 390356 89732 390420
rect 91140 390356 91204 390420
rect 96844 390356 96908 390420
rect 98132 390356 98196 390420
rect 104940 390356 105004 390420
rect 106412 390356 106476 390420
rect 107700 390356 107764 390420
rect 109356 390356 109420 390420
rect 115980 390416 116044 390420
rect 115980 390360 115994 390416
rect 115994 390360 116044 390416
rect 115980 390356 116044 390360
rect 120212 390416 120276 390420
rect 120212 390360 120262 390416
rect 120262 390360 120276 390416
rect 120212 390356 120276 390360
rect 111012 389404 111076 389468
rect 96476 389132 96540 389196
rect 95188 388996 95252 389060
rect 111748 389056 111812 389060
rect 111748 389000 111798 389056
rect 111798 389000 111812 389056
rect 111748 388996 111812 389000
rect 137140 388724 137204 388788
rect 99972 388316 100036 388380
rect 122604 387092 122668 387156
rect 114324 386276 114388 386340
rect 109172 383012 109236 383076
rect 95188 382876 95252 382940
rect 68692 378660 68756 378724
rect 68876 377300 68940 377364
rect 90220 371316 90284 371380
rect 95004 369820 95068 369884
rect 96660 369004 96724 369068
rect 99052 368324 99116 368388
rect 110644 367644 110708 367708
rect 138060 366284 138124 366348
rect 207980 365740 208044 365804
rect 118556 365604 118620 365668
rect 184060 364516 184124 364580
rect 233740 361660 233804 361724
rect 156460 360844 156524 360908
rect 120028 360300 120092 360364
rect 248460 360300 248524 360364
rect 322980 360164 323044 360228
rect 317460 358804 317524 358868
rect 151860 355540 151924 355604
rect 136036 355404 136100 355468
rect 113036 353636 113100 353700
rect 69796 352548 69860 352612
rect 231900 351868 231964 351932
rect 70164 351052 70228 351116
rect 229692 350780 229756 350844
rect 139716 349828 139780 349892
rect 67772 349692 67836 349756
rect 188292 349148 188356 349212
rect 277164 346428 277228 346492
rect 203012 345612 203076 345676
rect 133092 345204 133156 345268
rect 203012 345068 203076 345132
rect 240732 342212 240796 342276
rect 155172 341124 155236 341188
rect 244228 340852 244292 340916
rect 212580 339628 212644 339692
rect 230980 339492 231044 339556
rect 66668 335956 66732 336020
rect 84700 330516 84764 330580
rect 196572 330244 196636 330308
rect 154068 330108 154132 330172
rect 69612 329972 69676 330036
rect 70164 329972 70228 330036
rect 133092 329836 133156 329900
rect 133092 328476 133156 328540
rect 67588 328340 67652 328404
rect 68692 328340 68756 328404
rect 84700 327660 84764 327724
rect 154252 327660 154316 327724
rect 150388 327524 150452 327588
rect 155724 327524 155788 327588
rect 68692 327388 68756 327452
rect 66116 327116 66180 327180
rect 67220 326980 67284 327044
rect 77156 327116 77220 327180
rect 83964 327176 84028 327180
rect 83964 327120 83978 327176
rect 83978 327120 84028 327176
rect 83964 327116 84028 327120
rect 143396 326980 143460 327044
rect 154252 325212 154316 325276
rect 155724 324940 155788 325004
rect 154252 323580 154316 323644
rect 161980 323172 162044 323236
rect 155172 320724 155236 320788
rect 170260 320316 170324 320380
rect 156460 318684 156524 318748
rect 320220 316644 320284 316708
rect 222332 315284 222396 315348
rect 61884 313380 61948 313444
rect 270724 310660 270788 310724
rect 269068 309300 269132 309364
rect 67220 307940 67284 308004
rect 258396 307804 258460 307868
rect 315988 306640 316052 306644
rect 315988 306584 316002 306640
rect 316002 306584 316052 306640
rect 315988 306580 316052 306584
rect 322060 306444 322124 306508
rect 315988 306368 316052 306372
rect 315988 306312 316002 306368
rect 316002 306312 316052 306368
rect 315988 306308 316052 306312
rect 160692 303724 160756 303788
rect 218652 303724 218716 303788
rect 161980 302772 162044 302836
rect 227852 302772 227916 302836
rect 186820 301004 186884 301068
rect 287100 298420 287164 298484
rect 65932 297332 65996 297396
rect 237420 297332 237484 297396
rect 273300 296788 273364 296852
rect 316172 296788 316236 296852
rect 315988 296516 316052 296580
rect 180012 295972 180076 296036
rect 69428 295428 69492 295492
rect 161980 293524 162044 293588
rect 242940 293116 243004 293180
rect 284340 292708 284404 292772
rect 178540 292572 178604 292636
rect 66668 292164 66732 292228
rect 223620 291892 223684 291956
rect 270540 289988 270604 290052
rect 306420 287676 306484 287740
rect 191052 287268 191116 287332
rect 315988 287192 316052 287196
rect 315988 287136 316002 287192
rect 316002 287136 316052 287192
rect 315988 287132 316052 287136
rect 315988 287056 316052 287060
rect 315988 287000 316002 287056
rect 316002 287000 316052 287056
rect 315988 286996 316052 287000
rect 223804 285772 223868 285836
rect 223620 285636 223684 285700
rect 197308 284684 197372 284748
rect 245700 284548 245764 284612
rect 217548 284276 217612 284340
rect 224908 284276 224972 284340
rect 238524 284276 238588 284340
rect 216444 284004 216508 284068
rect 205404 283928 205468 283932
rect 205404 283872 205418 283928
rect 205418 283872 205468 283928
rect 205404 283868 205468 283872
rect 212396 283868 212460 283932
rect 214420 283928 214484 283932
rect 214420 283872 214470 283928
rect 214470 283872 214484 283928
rect 214420 283868 214484 283872
rect 215524 283868 215588 283932
rect 227484 283868 227548 283932
rect 237236 283868 237300 283932
rect 244228 284140 244292 284204
rect 244228 284004 244292 284068
rect 245700 282100 245764 282164
rect 244412 281012 244476 281076
rect 197308 280876 197372 280940
rect 67772 279380 67836 279444
rect 316172 277476 316236 277540
rect 315988 277400 316052 277404
rect 315988 277344 316002 277400
rect 316002 277344 316052 277400
rect 315988 277340 316052 277344
rect 248460 275300 248524 275364
rect 67772 268772 67836 268836
rect 316172 267820 316236 267884
rect 67956 267684 68020 267748
rect 316172 267684 316236 267748
rect 197124 267140 197188 267204
rect 244228 267004 244292 267068
rect 66668 266868 66732 266932
rect 199884 265236 199948 265300
rect 154620 260748 154684 260812
rect 61884 255988 61948 256052
rect 69428 253948 69492 254012
rect 67404 251908 67468 251972
rect 199516 248372 199580 248436
rect 200068 248372 200132 248436
rect 315988 248432 316052 248436
rect 315988 248376 316002 248432
rect 316002 248376 316052 248432
rect 315988 248372 316052 248376
rect 316172 248236 316236 248300
rect 200068 247556 200132 247620
rect 243492 246196 243556 246260
rect 69428 245924 69492 245988
rect 298140 244836 298204 244900
rect 154252 244564 154316 244628
rect 69244 244292 69308 244356
rect 67772 243476 67836 243540
rect 155172 243476 155236 243540
rect 245884 242932 245948 242996
rect 136036 242040 136100 242044
rect 136036 241984 136050 242040
rect 136050 241984 136100 242040
rect 136036 241980 136100 241984
rect 138060 241980 138124 242044
rect 151860 241844 151924 241908
rect 69244 241708 69308 241772
rect 172468 241768 172532 241772
rect 172468 241712 172518 241768
rect 172518 241712 172532 241768
rect 172468 241708 172532 241712
rect 148180 241496 148244 241500
rect 148180 241440 148194 241496
rect 148194 241440 148244 241496
rect 148180 241436 148244 241440
rect 195836 241436 195900 241500
rect 67404 241300 67468 241364
rect 195836 240620 195900 240684
rect 199884 240212 199948 240276
rect 245700 240212 245764 240276
rect 224908 240076 224972 240140
rect 227852 240076 227916 240140
rect 231900 240136 231964 240140
rect 231900 240080 231950 240136
rect 231950 240080 231964 240136
rect 231900 240076 231964 240080
rect 237420 240076 237484 240140
rect 315988 238776 316052 238780
rect 315988 238720 316002 238776
rect 316002 238720 316052 238776
rect 315988 238716 316052 238720
rect 203012 238580 203076 238644
rect 212580 238580 212644 238644
rect 222332 238580 222396 238644
rect 229692 238580 229756 238644
rect 233740 238580 233804 238644
rect 241284 238580 241348 238644
rect 315988 238640 316052 238644
rect 315988 238584 316002 238640
rect 316002 238584 316052 238640
rect 315988 238580 316052 238584
rect 218652 238444 218716 238508
rect 230980 238172 231044 238236
rect 223620 238036 223684 238100
rect 212580 237356 212644 237420
rect 137140 237220 137204 237284
rect 180012 237220 180076 237284
rect 207980 237220 208044 237284
rect 223620 237220 223684 237284
rect 137140 236948 137204 237012
rect 186268 236540 186332 236604
rect 67956 235860 68020 235924
rect 186268 235588 186332 235652
rect 139716 233956 139780 234020
rect 215524 233820 215588 233884
rect 143580 232868 143644 232932
rect 197124 231568 197188 231572
rect 197124 231512 197138 231568
rect 197138 231512 197188 231568
rect 197124 231508 197188 231512
rect 154620 231372 154684 231436
rect 245884 230420 245948 230484
rect 154068 230284 154132 230348
rect 278820 229876 278884 229940
rect 195836 229740 195900 229804
rect 316172 229060 316236 229124
rect 155172 228924 155236 228988
rect 316172 228924 316236 228988
rect 84700 227428 84764 227492
rect 245700 227428 245764 227492
rect 140820 224708 140884 224772
rect 276244 223484 276308 223548
rect 199516 222940 199580 223004
rect 217548 222260 217612 222324
rect 69796 222124 69860 222188
rect 273484 220220 273548 220284
rect 315988 219464 316052 219468
rect 315988 219408 316002 219464
rect 316002 219408 316052 219464
rect 315988 219404 316052 219408
rect 315988 219132 316052 219196
rect 77156 218588 77220 218652
rect 302188 216684 302252 216748
rect 178540 216412 178604 216476
rect 276612 215868 276676 215932
rect 65932 214508 65996 214572
rect 269252 213828 269316 213892
rect 277532 210564 277596 210628
rect 284524 210428 284588 210492
rect 310468 210292 310532 210356
rect 315988 209808 316052 209812
rect 315988 209752 316002 209808
rect 316002 209752 316052 209808
rect 315988 209748 316052 209752
rect 315988 209476 316052 209540
rect 66668 208932 66732 208996
rect 214420 207028 214484 207092
rect 154620 206212 154684 206276
rect 161980 206212 162044 206276
rect 69612 204172 69676 204236
rect 212580 204172 212644 204236
rect 213132 204172 213196 204236
rect 309180 202268 309244 202332
rect 315988 200152 316052 200156
rect 315988 200096 316002 200152
rect 316002 200096 316052 200152
rect 315988 200092 316052 200096
rect 315988 199820 316052 199884
rect 281764 199412 281828 199476
rect 150388 197916 150452 197980
rect 159220 197916 159284 197980
rect 168420 197916 168484 197980
rect 285812 196692 285876 196756
rect 242940 195876 243004 195940
rect 285628 195332 285692 195396
rect 241284 194108 241348 194172
rect 265756 193972 265820 194036
rect 309732 193836 309796 193900
rect 266308 193216 266372 193220
rect 266308 193160 266358 193216
rect 266358 193160 266372 193216
rect 266308 193156 266372 193160
rect 188292 192612 188356 192676
rect 83964 192476 84028 192540
rect 281580 192476 281644 192540
rect 280292 190572 280356 190636
rect 304948 190436 305012 190500
rect 315988 190496 316052 190500
rect 315988 190440 316002 190496
rect 316002 190440 316052 190496
rect 315988 190436 316052 190440
rect 315988 190360 316052 190364
rect 315988 190304 316002 190360
rect 316002 190304 316052 190360
rect 315988 190300 316052 190304
rect 133092 189892 133156 189956
rect 143396 189756 143460 189820
rect 275140 189620 275204 189684
rect 312308 189620 312372 189684
rect 272564 188396 272628 188460
rect 316172 188396 316236 188460
rect 313228 188260 313292 188324
rect 267780 185812 267844 185876
rect 237236 185676 237300 185740
rect 288940 185540 289004 185604
rect 216444 181324 216508 181388
rect 302372 181324 302436 181388
rect 315988 180916 316052 180980
rect 267964 180780 268028 180844
rect 315988 180704 316052 180708
rect 315988 180648 316002 180704
rect 316002 180648 316052 180704
rect 315988 180644 316052 180648
rect 305132 180100 305196 180164
rect 280292 179964 280356 180028
rect 301820 179964 301884 180028
rect 308628 178604 308692 178668
rect 110644 178196 110708 178260
rect 263916 178196 263980 178260
rect 290596 178060 290660 178124
rect 97028 177924 97092 177988
rect 100708 177516 100772 177580
rect 104572 177516 104636 177580
rect 105676 177516 105740 177580
rect 106964 177516 107028 177580
rect 113220 177516 113284 177580
rect 116900 177576 116964 177580
rect 116900 177520 116950 177576
rect 116950 177520 116964 177576
rect 116900 177516 116964 177520
rect 119476 177516 119540 177580
rect 120764 177516 120828 177580
rect 125732 177516 125796 177580
rect 129412 177516 129476 177580
rect 148180 177516 148244 177580
rect 258212 177516 258276 177580
rect 301268 177380 301332 177444
rect 112116 177108 112180 177172
rect 118372 177108 118436 177172
rect 108068 176972 108132 177036
rect 98316 176836 98380 176900
rect 101996 176760 102060 176764
rect 101996 176704 102046 176760
rect 102046 176704 102060 176760
rect 101996 176700 102060 176704
rect 115796 176760 115860 176764
rect 115796 176704 115846 176760
rect 115846 176704 115860 176760
rect 115796 176700 115860 176704
rect 124444 176760 124508 176764
rect 124444 176704 124494 176760
rect 124494 176704 124508 176760
rect 124444 176700 124508 176704
rect 127020 176700 127084 176764
rect 132356 176760 132420 176764
rect 132356 176704 132406 176760
rect 132406 176704 132420 176760
rect 132356 176700 132420 176704
rect 134380 176760 134444 176764
rect 134380 176704 134430 176760
rect 134430 176704 134444 176760
rect 134380 176700 134444 176704
rect 136036 176760 136100 176764
rect 136036 176704 136086 176760
rect 136086 176704 136100 176760
rect 136036 176700 136100 176704
rect 158852 176700 158916 176764
rect 265020 176700 265084 176764
rect 276612 176700 276676 176764
rect 306604 176564 306668 176628
rect 99420 176428 99484 176492
rect 103284 176428 103348 176492
rect 298140 175944 298204 175948
rect 298140 175888 298190 175944
rect 298190 175888 298204 175944
rect 298140 175884 298204 175888
rect 130700 175808 130764 175812
rect 130700 175752 130750 175808
rect 130750 175752 130764 175808
rect 130700 175748 130764 175752
rect 114324 175612 114388 175676
rect 164740 175612 164804 175676
rect 121868 175476 121932 175540
rect 109540 175340 109604 175404
rect 123070 174992 123134 174996
rect 123070 174936 123114 174992
rect 123114 174936 123134 174992
rect 123070 174932 123134 174936
rect 128102 174796 128166 174860
rect 133276 174660 133340 174724
rect 301268 173708 301332 173772
rect 266860 172484 266924 172548
rect 267964 172484 268028 172548
rect 315988 171260 316052 171324
rect 315988 171048 316052 171052
rect 315988 170992 316002 171048
rect 316002 170992 316052 171048
rect 315988 170988 316052 170992
rect 269252 169084 269316 169148
rect 305132 167860 305196 167924
rect 270356 166500 270420 166564
rect 268332 166228 268396 166292
rect 265020 165548 265084 165612
rect 272564 165548 272628 165612
rect 265572 164868 265636 164932
rect 164740 164324 164804 164388
rect 306604 164324 306668 164388
rect 273484 164248 273548 164252
rect 273484 164192 273498 164248
rect 273498 164192 273548 164248
rect 273484 164188 273548 164192
rect 269068 163780 269132 163844
rect 269620 163372 269684 163436
rect 270724 162692 270788 162756
rect 283788 162692 283852 162756
rect 276244 162420 276308 162484
rect 315988 161604 316052 161668
rect 274036 161468 274100 161532
rect 315988 161196 316052 161260
rect 267780 160108 267844 160172
rect 266308 159020 266372 159084
rect 270356 157388 270420 157452
rect 278820 157448 278884 157452
rect 278820 157392 278834 157448
rect 278834 157392 278884 157448
rect 278820 157388 278884 157392
rect 288388 157388 288452 157452
rect 268516 156844 268580 156908
rect 267044 156572 267108 156636
rect 266860 156164 266924 156228
rect 273484 155952 273548 155956
rect 273484 155896 273498 155952
rect 273498 155896 273548 155952
rect 273484 155892 273548 155896
rect 273300 154804 273364 154868
rect 265020 154456 265084 154460
rect 265020 154400 265070 154456
rect 265070 154400 265084 154456
rect 265020 154396 265084 154400
rect 265756 154260 265820 154324
rect 280108 153716 280172 153780
rect 280660 153308 280724 153372
rect 276796 152084 276860 152148
rect 315988 151872 316052 151876
rect 315988 151816 316002 151872
rect 316002 151816 316052 151872
rect 315988 151812 316052 151816
rect 315988 151540 316052 151604
rect 268332 151268 268396 151332
rect 266860 151132 266924 151196
rect 264100 150996 264164 151060
rect 269804 150996 269868 151060
rect 285812 150996 285876 151060
rect 264100 150452 264164 150516
rect 284524 150452 284588 150516
rect 268700 149908 268764 149972
rect 272564 149772 272628 149836
rect 283788 149636 283852 149700
rect 285076 149228 285140 149292
rect 267044 147732 267108 147796
rect 301820 147052 301884 147116
rect 281764 146372 281828 146436
rect 268516 145828 268580 145892
rect 271092 145828 271156 145892
rect 268332 145692 268396 145756
rect 284340 145556 284404 145620
rect 264100 145284 264164 145348
rect 278820 144740 278884 144804
rect 280292 144740 280356 144804
rect 184060 142700 184124 142764
rect 280844 143108 280908 143172
rect 267228 142700 267292 142764
rect 306420 142700 306484 142764
rect 265020 142428 265084 142492
rect 286180 142156 286244 142220
rect 315988 142216 316052 142220
rect 315988 142160 316002 142216
rect 316002 142160 316052 142216
rect 315988 142156 316052 142160
rect 315988 142080 316052 142084
rect 315988 142024 316002 142080
rect 316002 142024 316052 142080
rect 315988 142020 316052 142024
rect 213132 141340 213196 141404
rect 273852 141340 273916 141404
rect 277532 140932 277596 140996
rect 283788 140932 283852 140996
rect 273484 140796 273548 140860
rect 269804 140660 269868 140724
rect 288204 140388 288268 140452
rect 302372 140388 302436 140452
rect 270356 139980 270420 140044
rect 282500 139708 282564 139772
rect 285628 139436 285692 139500
rect 269804 138620 269868 138684
rect 288388 138348 288452 138412
rect 270356 138212 270420 138276
rect 290596 137940 290660 138004
rect 270540 137804 270604 137868
rect 281580 136852 281644 136916
rect 287100 136988 287164 137052
rect 282316 136852 282380 136916
rect 302188 136580 302252 136644
rect 278636 135628 278700 135692
rect 284892 135356 284956 135420
rect 278820 135220 278884 135284
rect 287836 134812 287900 134876
rect 278636 134540 278700 134604
rect 271644 134404 271708 134468
rect 288204 134404 288268 134468
rect 277900 134132 277964 134196
rect 290228 133724 290292 133788
rect 212396 133044 212460 133108
rect 265756 132772 265820 132836
rect 315988 132636 316052 132700
rect 315988 132424 316052 132428
rect 315988 132368 316002 132424
rect 316002 132368 316052 132424
rect 315988 132364 316052 132368
rect 282500 131684 282564 131748
rect 289124 131412 289188 131476
rect 286548 130324 286612 130388
rect 289860 128828 289924 128892
rect 287652 128420 287716 128484
rect 282316 128284 282380 128348
rect 269620 128148 269684 128212
rect 270356 127060 270420 127124
rect 308628 126788 308692 126852
rect 267228 124476 267292 124540
rect 266860 123524 266924 123588
rect 274036 123388 274100 123452
rect 315988 122980 316052 123044
rect 315988 122768 316052 122772
rect 315988 122712 316002 122768
rect 316002 122712 316052 122768
rect 315988 122708 316052 122712
rect 282316 122164 282380 122228
rect 266860 122028 266924 122092
rect 273300 121620 273364 121684
rect 269804 121212 269868 121276
rect 304948 120668 305012 120732
rect 279004 120260 279068 120324
rect 282316 119444 282380 119508
rect 276796 118084 276860 118148
rect 266308 117948 266372 118012
rect 276244 117948 276308 118012
rect 273300 117872 273364 117876
rect 273300 117816 273314 117872
rect 273314 117816 273364 117872
rect 273300 117812 273364 117816
rect 274036 117812 274100 117876
rect 310468 116180 310532 116244
rect 271644 115772 271708 115836
rect 286548 115772 286612 115836
rect 271276 114820 271340 114884
rect 269068 114684 269132 114748
rect 264100 113732 264164 113796
rect 287836 113188 287900 113252
rect 290044 113052 290108 113116
rect 268700 111964 268764 112028
rect 285628 111964 285692 112028
rect 287100 111964 287164 112028
rect 280660 111692 280724 111756
rect 267780 110468 267844 110532
rect 269620 109652 269684 109716
rect 309180 109380 309244 109444
rect 270356 109108 270420 109172
rect 312308 109108 312372 109172
rect 272564 108836 272628 108900
rect 285076 107476 285140 107540
rect 266308 106116 266372 106180
rect 280292 106116 280356 106180
rect 303660 106116 303724 106180
rect 267044 105436 267108 105500
rect 272564 104756 272628 104820
rect 268332 104620 268396 104684
rect 271092 104212 271156 104276
rect 290596 102716 290660 102780
rect 269068 102444 269132 102508
rect 269068 102308 269132 102372
rect 267964 102172 268028 102236
rect 316172 102172 316236 102236
rect 280844 102036 280908 102100
rect 286180 101356 286244 101420
rect 272564 100948 272628 101012
rect 284340 100948 284404 101012
rect 270540 100812 270604 100876
rect 273852 99996 273916 100060
rect 286180 99724 286244 99788
rect 264100 99044 264164 99108
rect 265572 98908 265636 98972
rect 273852 98772 273916 98836
rect 283788 98636 283852 98700
rect 283972 97956 284036 98020
rect 276612 97276 276676 97340
rect 166212 97140 166276 97204
rect 196572 97140 196636 97204
rect 252508 97140 252572 97204
rect 276244 97140 276308 97204
rect 276796 96596 276860 96660
rect 270724 96460 270788 96524
rect 257844 95976 257908 95980
rect 257844 95920 257894 95976
rect 257894 95920 257908 95976
rect 257844 95916 257908 95920
rect 260972 95976 261036 95980
rect 260972 95920 261022 95976
rect 261022 95920 261036 95976
rect 260972 95916 261036 95920
rect 270540 95916 270604 95980
rect 259316 95780 259380 95844
rect 279004 95780 279068 95844
rect 227484 95100 227548 95164
rect 113142 94964 113206 95028
rect 114508 94964 114572 95028
rect 151308 94964 151372 95028
rect 151766 94964 151830 95028
rect 289860 94888 289924 94892
rect 289860 94832 289874 94888
rect 289874 94832 289924 94888
rect 289860 94828 289924 94832
rect 124022 94752 124086 94756
rect 124022 94696 124034 94752
rect 124034 94696 124086 94752
rect 124022 94692 124086 94696
rect 131988 94012 132052 94076
rect 96660 93876 96724 93940
rect 99236 93740 99300 93804
rect 99604 93604 99668 93668
rect 205404 93604 205468 93668
rect 119660 93528 119724 93532
rect 119660 93472 119710 93528
rect 119710 93472 119724 93528
rect 119660 93468 119724 93472
rect 121684 93528 121748 93532
rect 121684 93472 121734 93528
rect 121734 93472 121748 93528
rect 121684 93468 121748 93472
rect 110092 93256 110156 93260
rect 110092 93200 110142 93256
rect 110142 93200 110156 93256
rect 110092 93196 110156 93200
rect 238524 93060 238588 93124
rect 86724 92380 86788 92444
rect 88932 92380 88996 92444
rect 109172 92380 109236 92444
rect 111196 92380 111260 92444
rect 114508 92440 114572 92444
rect 114508 92384 114522 92440
rect 114522 92384 114572 92440
rect 114508 92380 114572 92384
rect 136036 92440 136100 92444
rect 136036 92384 136086 92440
rect 136086 92384 136100 92440
rect 136036 92380 136100 92384
rect 151308 92440 151372 92444
rect 151308 92384 151358 92440
rect 151358 92384 151372 92440
rect 151308 92380 151372 92384
rect 120212 92108 120276 92172
rect 130700 92032 130764 92036
rect 130700 91976 130750 92032
rect 130750 91976 130764 92032
rect 130700 91972 130764 91976
rect 105676 91836 105740 91900
rect 84332 91700 84396 91764
rect 106412 91700 106476 91764
rect 114876 91760 114940 91764
rect 114876 91704 114926 91760
rect 114926 91704 114940 91760
rect 114876 91700 114940 91704
rect 116716 91700 116780 91764
rect 106780 91564 106844 91628
rect 98500 91428 98564 91492
rect 101996 91428 102060 91492
rect 125732 91564 125796 91628
rect 93900 91292 93964 91356
rect 101812 91292 101876 91356
rect 107700 91292 107764 91356
rect 115428 91292 115492 91356
rect 118004 91292 118068 91356
rect 122788 91352 122852 91356
rect 122788 91296 122838 91352
rect 122838 91296 122852 91352
rect 122788 91292 122852 91296
rect 125364 91352 125428 91356
rect 125364 91296 125414 91352
rect 125414 91296 125428 91352
rect 125364 91292 125428 91296
rect 126468 91292 126532 91356
rect 151676 91352 151740 91356
rect 151676 91296 151690 91352
rect 151690 91296 151740 91352
rect 151676 91292 151740 91296
rect 74764 91156 74828 91220
rect 85804 91156 85868 91220
rect 88012 91156 88076 91220
rect 90220 91156 90284 91220
rect 91324 91156 91388 91220
rect 92612 91156 92676 91220
rect 95004 91156 95068 91220
rect 96292 91156 96356 91220
rect 97212 91156 97276 91220
rect 98132 91156 98196 91220
rect 100524 91156 100588 91220
rect 100892 91156 100956 91220
rect 102548 91216 102612 91220
rect 102548 91160 102598 91216
rect 102598 91160 102612 91216
rect 102548 91156 102612 91160
rect 102732 91156 102796 91220
rect 104204 91216 104268 91220
rect 104204 91160 104254 91216
rect 104254 91160 104268 91216
rect 104204 91156 104268 91160
rect 104572 91156 104636 91220
rect 105492 91156 105556 91220
rect 108068 91156 108132 91220
rect 109540 91156 109604 91220
rect 110644 91156 110708 91220
rect 111932 91156 111996 91220
rect 112300 91156 112364 91220
rect 113220 91156 113284 91220
rect 114324 91216 114388 91220
rect 114324 91160 114338 91216
rect 114338 91160 114388 91216
rect 114324 91156 114388 91160
rect 115796 91216 115860 91220
rect 115796 91160 115846 91216
rect 115846 91160 115860 91216
rect 115796 91156 115860 91160
rect 117084 91156 117148 91220
rect 118188 91156 118252 91220
rect 119292 91156 119356 91220
rect 120580 91156 120644 91220
rect 122052 91156 122116 91220
rect 123156 91156 123220 91220
rect 124444 91156 124508 91220
rect 126652 91156 126716 91220
rect 127572 91156 127636 91220
rect 129412 91156 129476 91220
rect 133092 91156 133156 91220
rect 134380 91216 134444 91220
rect 134380 91160 134430 91216
rect 134430 91160 134444 91216
rect 134380 91156 134444 91160
rect 151492 91156 151556 91220
rect 151860 91156 151924 91220
rect 274036 89116 274100 89180
rect 259316 88164 259380 88228
rect 303660 88164 303724 88228
rect 267780 87620 267844 87684
rect 267964 86124 268028 86188
rect 166212 83948 166276 84012
rect 283972 83404 284036 83468
rect 270724 82316 270788 82380
rect 290596 80820 290660 80884
rect 271276 79460 271340 79524
rect 282316 76604 282380 76668
rect 276796 76468 276860 76532
rect 269620 74020 269684 74084
rect 267044 73884 267108 73948
rect 280292 69532 280356 69596
rect 289124 64092 289188 64156
rect 259500 63548 259564 63612
rect 277900 61372 277964 61436
rect 282132 58652 282196 58716
rect 266860 57156 266924 57220
rect 287100 54436 287164 54500
rect 269068 53076 269132 53140
rect 265756 51716 265820 51780
rect 264100 50220 264164 50284
rect 286180 48860 286244 48924
rect 61884 47500 61948 47564
rect 284340 44780 284404 44844
rect 287652 37844 287716 37908
rect 263916 35124 263980 35188
rect 66116 26828 66180 26892
rect 273852 21252 273916 21316
rect 67772 19892 67836 19956
rect 260972 18532 261036 18596
rect 284892 17172 284956 17236
rect 285628 15812 285692 15876
rect 186820 14452 186884 14516
rect 317460 11596 317524 11660
rect 165660 10236 165724 10300
rect 191052 10236 191116 10300
rect 170260 8876 170324 8940
rect 168420 4796 168484 4860
rect 322060 4796 322124 4860
rect 277164 3980 277228 4044
rect 309732 3980 309796 4044
rect 252508 3436 252572 3500
rect 288940 3436 289004 3500
rect 313228 3436 313292 3500
rect 320220 3436 320284 3500
rect 322980 3436 323044 3500
rect 275140 3300 275204 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 69611 702540 69677 702541
rect 69611 702476 69612 702540
rect 69676 702476 69677 702540
rect 69611 702475 69677 702476
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 591166 67574 608058
rect 69614 586530 69674 702475
rect 73794 687454 74414 704282
rect 76051 699820 76117 699821
rect 76051 699756 76052 699820
rect 76116 699756 76117 699820
rect 76051 699755 76117 699756
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 591166 74414 614898
rect 69430 586470 69674 586530
rect 67771 583812 67837 583813
rect 67771 583748 67772 583812
rect 67836 583748 67837 583812
rect 67771 583747 67837 583748
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 66667 550900 66733 550901
rect 66667 550836 66668 550900
rect 66732 550836 66733 550900
rect 66667 550835 66733 550836
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 61883 393276 61949 393277
rect 61883 393212 61884 393276
rect 61948 393212 61949 393276
rect 61883 393211 61949 393212
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 61886 313445 61946 393211
rect 63234 388894 63854 424338
rect 66670 410549 66730 550835
rect 66954 536614 67574 537166
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 446407 67574 464058
rect 67774 457469 67834 583747
rect 69430 581909 69490 586470
rect 69427 581908 69493 581909
rect 69427 581844 69428 581908
rect 69492 581844 69493 581908
rect 69427 581843 69493 581844
rect 72679 579454 72999 579486
rect 72679 579218 72721 579454
rect 72957 579218 72999 579454
rect 72679 579134 72999 579218
rect 72679 578898 72721 579134
rect 72957 578898 72999 579134
rect 72679 578866 72999 578898
rect 75644 561454 75964 561486
rect 75644 561218 75686 561454
rect 75922 561218 75964 561454
rect 75644 561134 75964 561218
rect 75644 560898 75686 561134
rect 75922 560898 75964 561134
rect 75644 560866 75964 560898
rect 72679 543454 72999 543486
rect 72679 543218 72721 543454
rect 72957 543218 72999 543454
rect 72679 543134 72999 543218
rect 72679 542898 72721 543134
rect 72957 542898 72999 543134
rect 72679 542866 72999 542898
rect 76054 538117 76114 699755
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 591166 78134 618618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 591166 81854 622338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 591166 85574 626058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 88195 588572 88261 588573
rect 88195 588508 88196 588572
rect 88260 588508 88261 588572
rect 88195 588507 88261 588508
rect 88198 585717 88258 588507
rect 88195 585716 88261 585717
rect 88195 585652 88196 585716
rect 88260 585652 88261 585716
rect 88195 585651 88261 585652
rect 78609 579454 78929 579486
rect 78609 579218 78651 579454
rect 78887 579218 78929 579454
rect 78609 579134 78929 579218
rect 78609 578898 78651 579134
rect 78887 578898 78929 579134
rect 78609 578866 78929 578898
rect 84540 579454 84860 579486
rect 84540 579218 84582 579454
rect 84818 579218 84860 579454
rect 84540 579134 84860 579218
rect 84540 578898 84582 579134
rect 84818 578898 84860 579134
rect 84540 578866 84860 578898
rect 81575 561454 81895 561486
rect 81575 561218 81617 561454
rect 81853 561218 81895 561454
rect 81575 561134 81895 561218
rect 81575 560898 81617 561134
rect 81853 560898 81895 561134
rect 81575 560866 81895 560898
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 78609 543454 78929 543486
rect 78609 543218 78651 543454
rect 78887 543218 78929 543454
rect 78609 543134 78929 543218
rect 78609 542898 78651 543134
rect 78887 542898 78929 543134
rect 78609 542866 78929 542898
rect 84540 543454 84860 543486
rect 84540 543218 84582 543454
rect 84818 543218 84860 543454
rect 84540 543134 84860 543218
rect 84540 542898 84582 543134
rect 84818 542898 84860 543134
rect 84540 542866 84860 542898
rect 76051 538116 76117 538117
rect 76051 538052 76052 538116
rect 76116 538052 76117 538116
rect 76051 538051 76117 538052
rect 69611 535532 69677 535533
rect 69611 535468 69612 535532
rect 69676 535468 69677 535532
rect 69611 535467 69677 535468
rect 71819 535532 71885 535533
rect 71819 535468 71820 535532
rect 71884 535468 71885 535532
rect 71819 535467 71885 535468
rect 67771 457468 67837 457469
rect 67771 457404 67772 457468
rect 67836 457404 67837 457468
rect 67771 457403 67837 457404
rect 68875 444276 68941 444277
rect 68875 444212 68876 444276
rect 68940 444212 68941 444276
rect 68875 444211 68941 444212
rect 66667 410548 66733 410549
rect 66667 410484 66668 410548
rect 66732 410484 66733 410548
rect 66667 410483 66733 410484
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 66954 356614 67574 388356
rect 68691 378724 68757 378725
rect 68691 378660 68692 378724
rect 68756 378660 68757 378724
rect 68691 378659 68757 378660
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66667 336020 66733 336021
rect 66667 335956 66668 336020
rect 66732 335956 66733 336020
rect 66667 335955 66733 335956
rect 66115 327180 66181 327181
rect 66115 327116 66116 327180
rect 66180 327116 66181 327180
rect 66115 327115 66181 327116
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 61883 313444 61949 313445
rect 61883 313380 61884 313444
rect 61948 313380 61949 313444
rect 61883 313379 61949 313380
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 63234 280894 63854 316338
rect 65931 297396 65997 297397
rect 65931 297332 65932 297396
rect 65996 297332 65997 297396
rect 65931 297331 65997 297332
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 61883 256052 61949 256053
rect 61883 255988 61884 256052
rect 61948 255988 61949 256052
rect 61883 255987 61949 255988
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 61886 47565 61946 255987
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 65934 214573 65994 297331
rect 65931 214572 65997 214573
rect 65931 214508 65932 214572
rect 65996 214508 65997 214572
rect 65931 214507 65997 214508
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 61883 47564 61949 47565
rect 61883 47500 61884 47564
rect 61948 47500 61949 47564
rect 61883 47499 61949 47500
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 66118 26893 66178 327115
rect 66670 292229 66730 335955
rect 66954 329592 67574 356058
rect 67771 349756 67837 349757
rect 67771 349692 67772 349756
rect 67836 349692 67837 349756
rect 67771 349691 67837 349692
rect 67587 328404 67653 328405
rect 67587 328340 67588 328404
rect 67652 328340 67653 328404
rect 67587 328339 67653 328340
rect 67219 327044 67285 327045
rect 67219 326980 67220 327044
rect 67284 326980 67285 327044
rect 67219 326979 67285 326980
rect 67222 308005 67282 326979
rect 67219 308004 67285 308005
rect 67219 307940 67220 308004
rect 67284 307940 67285 308004
rect 67219 307939 67285 307940
rect 66667 292228 66733 292229
rect 66667 292164 66668 292228
rect 66732 292164 66733 292228
rect 66667 292163 66733 292164
rect 67590 277410 67650 328339
rect 67774 279445 67834 349691
rect 68694 328405 68754 378659
rect 68878 377365 68938 444211
rect 69614 414030 69674 535467
rect 69062 413970 69674 414030
rect 69062 405650 69122 413970
rect 69246 408310 69674 408370
rect 69246 408237 69306 408310
rect 69243 408236 69309 408237
rect 69243 408172 69244 408236
rect 69308 408172 69309 408236
rect 69243 408171 69309 408172
rect 69614 407826 69674 408310
rect 69614 407766 70226 407826
rect 69062 405590 69674 405650
rect 69614 404290 69674 405590
rect 70166 404370 70226 407766
rect 69062 404230 69674 404290
rect 69982 404310 70226 404370
rect 69062 396130 69122 404230
rect 69982 400890 70042 404310
rect 69798 400830 70042 400890
rect 69062 396070 69674 396130
rect 69614 390421 69674 396070
rect 69611 390420 69677 390421
rect 69611 390356 69612 390420
rect 69676 390356 69677 390420
rect 69611 390355 69677 390356
rect 68875 377364 68941 377365
rect 68875 377300 68876 377364
rect 68940 377300 68941 377364
rect 68875 377299 68941 377300
rect 69798 352613 69858 400830
rect 71822 390421 71882 535467
rect 73794 507454 74414 537166
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 446407 74414 470898
rect 77514 511174 78134 537166
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 446407 78134 474618
rect 81234 514894 81854 537166
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 446407 81854 478338
rect 84954 518614 85574 537166
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446407 85574 482058
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 89667 461548 89733 461549
rect 89667 461484 89668 461548
rect 89732 461484 89733 461548
rect 89667 461483 89733 461484
rect 72978 435454 73298 435486
rect 72978 435218 73020 435454
rect 73256 435218 73298 435454
rect 72978 435134 73298 435218
rect 72978 434898 73020 435134
rect 73256 434898 73298 435134
rect 72978 434866 73298 434898
rect 88338 417454 88658 417486
rect 88338 417218 88380 417454
rect 88616 417218 88658 417454
rect 88338 417134 88658 417218
rect 88338 416898 88380 417134
rect 88616 416898 88658 417134
rect 88338 416866 88658 416898
rect 72978 399454 73298 399486
rect 72978 399218 73020 399454
rect 73256 399218 73298 399454
rect 72978 399134 73298 399218
rect 72978 398898 73020 399134
rect 73256 398898 73298 399134
rect 72978 398866 73298 398898
rect 89670 390421 89730 461483
rect 91139 456244 91205 456245
rect 91139 456180 91140 456244
rect 91204 456180 91205 456244
rect 91139 456179 91205 456180
rect 90219 445908 90285 445909
rect 90219 445844 90220 445908
rect 90284 445844 90285 445908
rect 90219 445843 90285 445844
rect 71819 390420 71885 390421
rect 71819 390356 71820 390420
rect 71884 390356 71885 390420
rect 71819 390355 71885 390356
rect 89667 390420 89733 390421
rect 89667 390356 89668 390420
rect 89732 390356 89733 390420
rect 89667 390355 89733 390356
rect 73794 363454 74414 388356
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 69795 352612 69861 352613
rect 69795 352548 69796 352612
rect 69860 352548 69861 352612
rect 69795 352547 69861 352548
rect 70163 351116 70229 351117
rect 70163 351052 70164 351116
rect 70228 351052 70229 351116
rect 70163 351051 70229 351052
rect 70166 330037 70226 351051
rect 69611 330036 69677 330037
rect 69611 329972 69612 330036
rect 69676 329972 69677 330036
rect 69611 329971 69677 329972
rect 70163 330036 70229 330037
rect 70163 329972 70164 330036
rect 70228 329972 70229 330036
rect 70163 329971 70229 329972
rect 68691 328404 68757 328405
rect 68691 328340 68692 328404
rect 68756 328340 68757 328404
rect 68691 328339 68757 328340
rect 68694 327453 68754 328339
rect 68691 327452 68757 327453
rect 68691 327388 68692 327452
rect 68756 327388 68757 327452
rect 68691 327387 68757 327388
rect 69614 296730 69674 329971
rect 73794 329592 74414 362898
rect 77514 367174 78134 388356
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 329592 78134 330618
rect 81234 370894 81854 388356
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 329592 81854 334338
rect 84954 374614 85574 388356
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 90222 371381 90282 445843
rect 91142 390421 91202 456179
rect 91794 453454 92414 488898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 92611 460188 92677 460189
rect 92611 460124 92612 460188
rect 92676 460124 92677 460188
rect 92611 460123 92677 460124
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 446407 92414 452898
rect 92614 390965 92674 460123
rect 95514 457174 96134 492618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 99971 550764 100037 550765
rect 99971 550700 99972 550764
rect 100036 550700 100037 550764
rect 99971 550699 100037 550700
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 96843 462908 96909 462909
rect 96843 462844 96844 462908
rect 96908 462844 96909 462908
rect 96843 462843 96909 462844
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95187 449172 95253 449173
rect 95187 449108 95188 449172
rect 95252 449108 95253 449172
rect 95187 449107 95253 449108
rect 95003 445772 95069 445773
rect 95003 445708 95004 445772
rect 95068 445708 95069 445772
rect 95003 445707 95069 445708
rect 92611 390964 92677 390965
rect 92611 390900 92612 390964
rect 92676 390900 92677 390964
rect 92611 390899 92677 390900
rect 91139 390420 91205 390421
rect 91139 390356 91140 390420
rect 91204 390356 91205 390420
rect 91139 390355 91205 390356
rect 91794 381454 92414 388356
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 90219 371380 90285 371381
rect 90219 371316 90220 371380
rect 90284 371316 90285 371380
rect 90219 371315 90285 371316
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84699 330580 84765 330581
rect 84699 330516 84700 330580
rect 84764 330516 84765 330580
rect 84699 330515 84765 330516
rect 84702 327725 84762 330515
rect 84954 329592 85574 338058
rect 91794 345454 92414 380898
rect 95006 369885 95066 445707
rect 95190 389061 95250 449107
rect 95514 446407 96134 456618
rect 96475 446452 96541 446453
rect 96475 446388 96476 446452
rect 96540 446388 96541 446452
rect 96475 446387 96541 446388
rect 96478 389197 96538 446387
rect 96659 445772 96725 445773
rect 96659 445708 96660 445772
rect 96724 445708 96725 445772
rect 96659 445707 96725 445708
rect 96475 389196 96541 389197
rect 96475 389132 96476 389196
rect 96540 389132 96541 389196
rect 96475 389131 96541 389132
rect 95187 389060 95253 389061
rect 95187 388996 95188 389060
rect 95252 388996 95253 389060
rect 95187 388995 95253 388996
rect 95190 382941 95250 388995
rect 95514 385174 96134 388356
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95187 382940 95253 382941
rect 95187 382876 95188 382940
rect 95252 382876 95253 382940
rect 95187 382875 95253 382876
rect 95003 369884 95069 369885
rect 95003 369820 95004 369884
rect 95068 369820 95069 369884
rect 95003 369819 95069 369820
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 329592 92414 344898
rect 95514 349174 96134 384618
rect 96662 369069 96722 445707
rect 96846 390421 96906 462843
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 98131 457468 98197 457469
rect 98131 457404 98132 457468
rect 98196 457404 98197 457468
rect 98131 457403 98197 457404
rect 98134 390421 98194 457403
rect 99234 446407 99854 460338
rect 99051 445772 99117 445773
rect 99051 445708 99052 445772
rect 99116 445708 99117 445772
rect 99051 445707 99117 445708
rect 96843 390420 96909 390421
rect 96843 390356 96844 390420
rect 96908 390356 96909 390420
rect 96843 390355 96909 390356
rect 98131 390420 98197 390421
rect 98131 390356 98132 390420
rect 98196 390356 98197 390420
rect 98131 390355 98197 390356
rect 96659 369068 96725 369069
rect 96659 369004 96660 369068
rect 96724 369004 96725 369068
rect 96659 369003 96725 369004
rect 99054 368389 99114 445707
rect 99974 388381 100034 550699
rect 102954 536614 103574 572058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109355 546548 109421 546549
rect 109355 546484 109356 546548
rect 109420 546484 109421 546548
rect 109355 546483 109421 546484
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 106411 467124 106477 467125
rect 106411 467060 106412 467124
rect 106476 467060 106477 467124
rect 106411 467059 106477 467060
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102731 460188 102797 460189
rect 102731 460124 102732 460188
rect 102796 460124 102797 460188
rect 102731 460123 102797 460124
rect 100707 456108 100773 456109
rect 100707 456044 100708 456108
rect 100772 456044 100773 456108
rect 100707 456043 100773 456044
rect 100710 390557 100770 456043
rect 102734 390965 102794 460123
rect 102954 446407 103574 464058
rect 104939 459644 105005 459645
rect 104939 459580 104940 459644
rect 105004 459580 105005 459644
rect 104939 459579 105005 459580
rect 103698 435454 104018 435486
rect 103698 435218 103740 435454
rect 103976 435218 104018 435454
rect 103698 435134 104018 435218
rect 103698 434898 103740 435134
rect 103976 434898 104018 435134
rect 103698 434866 104018 434898
rect 103698 399454 104018 399486
rect 103698 399218 103740 399454
rect 103976 399218 104018 399454
rect 103698 399134 104018 399218
rect 103698 398898 103740 399134
rect 103976 398898 104018 399134
rect 103698 398866 104018 398898
rect 102731 390964 102797 390965
rect 102731 390900 102732 390964
rect 102796 390900 102797 390964
rect 102731 390899 102797 390900
rect 100707 390556 100773 390557
rect 100707 390492 100708 390556
rect 100772 390492 100773 390556
rect 100707 390491 100773 390492
rect 104942 390421 105002 459579
rect 106414 390421 106474 467059
rect 107699 458828 107765 458829
rect 107699 458764 107700 458828
rect 107764 458764 107765 458828
rect 107699 458763 107765 458764
rect 107702 390421 107762 458763
rect 109171 444684 109237 444685
rect 109171 444620 109172 444684
rect 109236 444620 109237 444684
rect 109171 444619 109237 444620
rect 104939 390420 105005 390421
rect 104939 390356 104940 390420
rect 105004 390356 105005 390420
rect 104939 390355 105005 390356
rect 106411 390420 106477 390421
rect 106411 390356 106412 390420
rect 106476 390356 106477 390420
rect 106411 390355 106477 390356
rect 107699 390420 107765 390421
rect 107699 390356 107700 390420
rect 107764 390356 107765 390420
rect 107699 390355 107765 390356
rect 99971 388380 100037 388381
rect 99051 368388 99117 368389
rect 99051 368324 99052 368388
rect 99116 368324 99117 368388
rect 99051 368323 99117 368324
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 329592 96134 348618
rect 99234 352894 99854 388356
rect 99971 388316 99972 388380
rect 100036 388316 100037 388380
rect 99971 388315 100037 388316
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 329592 99854 352338
rect 102954 356614 103574 388356
rect 109174 383077 109234 444619
rect 109358 390421 109418 546483
rect 109794 543454 110414 578898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 111011 553484 111077 553485
rect 111011 553420 111012 553484
rect 111076 553420 111077 553484
rect 111011 553419 111077 553420
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 446407 110414 470898
rect 110643 445772 110709 445773
rect 110643 445708 110644 445772
rect 110708 445708 110709 445772
rect 110643 445707 110709 445708
rect 109355 390420 109421 390421
rect 109355 390356 109356 390420
rect 109420 390356 109421 390420
rect 109355 390355 109421 390356
rect 109171 383076 109237 383077
rect 109171 383012 109172 383076
rect 109236 383012 109237 383076
rect 109171 383011 109237 383012
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 329592 103574 356058
rect 109794 363454 110414 388356
rect 110646 367709 110706 445707
rect 111014 389469 111074 553419
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 111747 461548 111813 461549
rect 111747 461484 111748 461548
rect 111812 461484 111813 461548
rect 111747 461483 111813 461484
rect 111011 389468 111077 389469
rect 111011 389404 111012 389468
rect 111076 389404 111077 389468
rect 111011 389403 111077 389404
rect 111750 389061 111810 461483
rect 113514 446407 114134 474618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 119475 580276 119541 580277
rect 119475 580212 119476 580276
rect 119540 580212 119541 580276
rect 119475 580211 119541 580212
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 115979 456108 116045 456109
rect 115979 456044 115980 456108
rect 116044 456044 116045 456108
rect 115979 456043 116045 456044
rect 114323 445772 114389 445773
rect 114323 445708 114324 445772
rect 114388 445708 114389 445772
rect 114323 445707 114389 445708
rect 113035 392052 113101 392053
rect 113035 391988 113036 392052
rect 113100 391988 113101 392052
rect 113035 391987 113101 391988
rect 111747 389060 111813 389061
rect 111747 388996 111748 389060
rect 111812 388996 111813 389060
rect 111747 388995 111813 388996
rect 110643 367708 110709 367709
rect 110643 367644 110644 367708
rect 110708 367644 110709 367708
rect 110643 367643 110709 367644
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 329592 110414 362898
rect 113038 353701 113098 391987
rect 113514 367174 114134 388356
rect 114326 386341 114386 445707
rect 115982 390421 116042 456043
rect 117234 446407 117854 478338
rect 118555 445772 118621 445773
rect 118555 445708 118556 445772
rect 118620 445708 118621 445772
rect 118555 445707 118621 445708
rect 115979 390420 116045 390421
rect 115979 390356 115980 390420
rect 116044 390356 116045 390420
rect 115979 390355 116045 390356
rect 114323 386340 114389 386341
rect 114323 386276 114324 386340
rect 114388 386276 114389 386340
rect 114323 386275 114389 386276
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113035 353700 113101 353701
rect 113035 353636 113036 353700
rect 113100 353636 113101 353700
rect 113035 353635 113101 353636
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 329592 114134 330618
rect 117234 370894 117854 388356
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 118558 365669 118618 445707
rect 119478 441630 119538 580211
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120211 462908 120277 462909
rect 120211 462844 120212 462908
rect 120276 462844 120277 462908
rect 120211 462843 120277 462844
rect 119843 444684 119909 444685
rect 119843 444620 119844 444684
rect 119908 444620 119909 444684
rect 119843 444619 119909 444620
rect 119846 443730 119906 444619
rect 119846 443670 120090 443730
rect 120030 442781 120090 443670
rect 120027 442780 120093 442781
rect 120027 442716 120028 442780
rect 120092 442716 120093 442780
rect 120027 442715 120093 442716
rect 120214 441630 120274 462843
rect 120954 446407 121574 482058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 122603 469844 122669 469845
rect 122603 469780 122604 469844
rect 122668 469780 122669 469844
rect 122603 469779 122669 469780
rect 121683 451892 121749 451893
rect 121683 451828 121684 451892
rect 121748 451828 121749 451892
rect 121683 451827 121749 451828
rect 119478 441570 119906 441630
rect 120214 441570 120642 441630
rect 119846 432170 119906 441570
rect 120395 434756 120461 434757
rect 120395 434692 120396 434756
rect 120460 434692 120461 434756
rect 120395 434691 120461 434692
rect 119846 432110 120274 432170
rect 120214 431493 120274 432110
rect 120211 431492 120277 431493
rect 120211 431428 120212 431492
rect 120276 431428 120277 431492
rect 120211 431427 120277 431428
rect 120398 427830 120458 434691
rect 120030 427770 120458 427830
rect 119058 417454 119378 417486
rect 119058 417218 119100 417454
rect 119336 417218 119378 417454
rect 119058 417134 119378 417218
rect 119058 416898 119100 417134
rect 119336 416898 119378 417134
rect 119058 416866 119378 416898
rect 118555 365668 118621 365669
rect 118555 365604 118556 365668
rect 118620 365604 118621 365668
rect 118555 365603 118621 365604
rect 120030 360365 120090 427770
rect 120582 412650 120642 441570
rect 120214 412590 120642 412650
rect 120214 390421 120274 412590
rect 121686 403749 121746 451827
rect 122606 437490 122666 469779
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 123339 447676 123405 447677
rect 123339 447612 123340 447676
rect 123404 447612 123405 447676
rect 123339 447611 123405 447612
rect 123342 444277 123402 447611
rect 123339 444276 123405 444277
rect 123339 444212 123340 444276
rect 123404 444212 123405 444276
rect 123339 444211 123405 444212
rect 122606 437430 122850 437490
rect 122790 435301 122850 437430
rect 122787 435300 122853 435301
rect 122787 435236 122788 435300
rect 122852 435236 122853 435300
rect 122787 435235 122853 435236
rect 122603 425644 122669 425645
rect 122603 425580 122604 425644
rect 122668 425580 122669 425644
rect 122603 425579 122669 425580
rect 121683 403748 121749 403749
rect 121683 403684 121684 403748
rect 121748 403684 121749 403748
rect 121683 403683 121749 403684
rect 120211 390420 120277 390421
rect 120211 390356 120212 390420
rect 120276 390356 120277 390420
rect 120211 390355 120277 390356
rect 120954 374614 121574 388356
rect 122606 387157 122666 425579
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 122603 387156 122669 387157
rect 122603 387092 122604 387156
rect 122668 387092 122669 387156
rect 122603 387091 122669 387092
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120027 360364 120093 360365
rect 120027 360300 120028 360364
rect 120092 360300 120093 360364
rect 120027 360299 120093 360300
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 329592 117854 334338
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 329592 121574 338058
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 329592 128414 344898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 329592 132134 348618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 143579 442372 143645 442373
rect 143579 442308 143580 442372
rect 143644 442308 143645 442372
rect 143579 442307 143645 442308
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 140819 401708 140885 401709
rect 140819 401644 140820 401708
rect 140884 401644 140885 401708
rect 140819 401643 140885 401644
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 137139 388788 137205 388789
rect 137139 388724 137140 388788
rect 137204 388724 137205 388788
rect 137139 388723 137205 388724
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 136035 355468 136101 355469
rect 136035 355404 136036 355468
rect 136100 355404 136101 355468
rect 136035 355403 136101 355404
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 133091 345268 133157 345269
rect 133091 345204 133092 345268
rect 133156 345204 133157 345268
rect 133091 345203 133157 345204
rect 133094 329901 133154 345203
rect 133091 329900 133157 329901
rect 133091 329836 133092 329900
rect 133156 329836 133157 329900
rect 133091 329835 133157 329836
rect 135234 329592 135854 352338
rect 133091 328540 133157 328541
rect 133091 328476 133092 328540
rect 133156 328476 133157 328540
rect 133091 328475 133157 328476
rect 84699 327724 84765 327725
rect 84699 327660 84700 327724
rect 84764 327660 84765 327724
rect 84699 327659 84765 327660
rect 77155 327180 77221 327181
rect 77155 327116 77156 327180
rect 77220 327116 77221 327180
rect 77155 327115 77221 327116
rect 83963 327180 84029 327181
rect 83963 327116 83964 327180
rect 84028 327116 84029 327180
rect 83963 327115 84029 327116
rect 69430 296670 69674 296730
rect 69430 295493 69490 296670
rect 69427 295492 69493 295493
rect 69427 295428 69428 295492
rect 69492 295428 69493 295492
rect 69427 295427 69493 295428
rect 72978 291454 73298 291486
rect 72978 291218 73020 291454
rect 73256 291218 73298 291454
rect 72978 291134 73298 291218
rect 72978 290898 73020 291134
rect 73256 290898 73298 291134
rect 72978 290866 73298 290898
rect 67771 279444 67837 279445
rect 67771 279380 67772 279444
rect 67836 279380 67837 279444
rect 67771 279379 67837 279380
rect 67590 277350 67834 277410
rect 67774 268837 67834 277350
rect 67771 268836 67837 268837
rect 67771 268772 67772 268836
rect 67836 268772 67837 268836
rect 67771 268771 67837 268772
rect 67955 267748 68021 267749
rect 67955 267684 67956 267748
rect 68020 267684 68021 267748
rect 67955 267683 68021 267684
rect 66667 266932 66733 266933
rect 66667 266868 66668 266932
rect 66732 266868 66733 266932
rect 66667 266867 66733 266868
rect 66670 208997 66730 266867
rect 67403 251972 67469 251973
rect 67403 251908 67404 251972
rect 67468 251908 67469 251972
rect 67403 251907 67469 251908
rect 67406 241365 67466 251907
rect 67771 243540 67837 243541
rect 67771 243476 67772 243540
rect 67836 243476 67837 243540
rect 67771 243475 67837 243476
rect 67403 241364 67469 241365
rect 67403 241300 67404 241364
rect 67468 241300 67469 241364
rect 67403 241299 67469 241300
rect 66954 212614 67574 239592
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66667 208996 66733 208997
rect 66667 208932 66668 208996
rect 66732 208932 66733 208996
rect 66667 208931 66733 208932
rect 66954 176600 67574 212058
rect 66954 68614 67574 93100
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 66115 26892 66181 26893
rect 66115 26828 66116 26892
rect 66180 26828 66181 26892
rect 66115 26827 66181 26828
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 67774 19957 67834 243475
rect 67958 235925 68018 267683
rect 72978 255454 73298 255486
rect 72978 255218 73020 255454
rect 73256 255218 73298 255454
rect 72978 255134 73298 255218
rect 72978 254898 73020 255134
rect 73256 254898 73298 255134
rect 72978 254866 73298 254898
rect 69427 254012 69493 254013
rect 69427 253948 69428 254012
rect 69492 253948 69493 254012
rect 69427 253947 69493 253948
rect 69430 248430 69490 253947
rect 69246 248370 69490 248430
rect 69246 245170 69306 248370
rect 69430 246470 69858 246530
rect 69430 245989 69490 246470
rect 69427 245988 69493 245989
rect 69427 245924 69428 245988
rect 69492 245924 69493 245988
rect 69427 245923 69493 245924
rect 69246 245110 69490 245170
rect 69243 244356 69309 244357
rect 69243 244292 69244 244356
rect 69308 244292 69309 244356
rect 69243 244291 69309 244292
rect 69246 241773 69306 244291
rect 69430 243810 69490 245110
rect 69430 243750 69674 243810
rect 69243 241772 69309 241773
rect 69243 241708 69244 241772
rect 69308 241708 69309 241772
rect 69243 241707 69309 241708
rect 67955 235924 68021 235925
rect 67955 235860 67956 235924
rect 68020 235860 68021 235924
rect 67955 235859 68021 235860
rect 69614 204237 69674 243750
rect 69798 222189 69858 246470
rect 69795 222188 69861 222189
rect 69795 222124 69796 222188
rect 69860 222124 69861 222188
rect 69795 222123 69861 222124
rect 73794 219454 74414 239592
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 69611 204236 69677 204237
rect 69611 204172 69612 204236
rect 69676 204172 69677 204236
rect 69611 204171 69677 204172
rect 73794 183454 74414 218898
rect 77158 218653 77218 327115
rect 77514 223174 78134 239592
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77155 218652 77221 218653
rect 77155 218588 77156 218652
rect 77220 218588 77221 218652
rect 77155 218587 77221 218588
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 176600 74414 182898
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 176600 78134 186618
rect 81234 226894 81854 239592
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 83966 192541 84026 327115
rect 84702 227493 84762 327659
rect 88338 309454 88658 309486
rect 88338 309218 88380 309454
rect 88616 309218 88658 309454
rect 88338 309134 88658 309218
rect 88338 308898 88380 309134
rect 88616 308898 88658 309134
rect 88338 308866 88658 308898
rect 119058 309454 119378 309486
rect 119058 309218 119100 309454
rect 119336 309218 119378 309454
rect 119058 309134 119378 309218
rect 119058 308898 119100 309134
rect 119336 308898 119378 309134
rect 119058 308866 119378 308898
rect 103698 291454 104018 291486
rect 103698 291218 103740 291454
rect 103976 291218 104018 291454
rect 103698 291134 104018 291218
rect 103698 290898 103740 291134
rect 103976 290898 104018 291134
rect 103698 290866 104018 290898
rect 88338 273454 88658 273486
rect 88338 273218 88380 273454
rect 88616 273218 88658 273454
rect 88338 273134 88658 273218
rect 88338 272898 88380 273134
rect 88616 272898 88658 273134
rect 88338 272866 88658 272898
rect 119058 273454 119378 273486
rect 119058 273218 119100 273454
rect 119336 273218 119378 273454
rect 119058 273134 119378 273218
rect 119058 272898 119100 273134
rect 119336 272898 119378 273134
rect 119058 272866 119378 272898
rect 103698 255454 104018 255486
rect 103698 255218 103740 255454
rect 103976 255218 104018 255454
rect 103698 255134 104018 255218
rect 103698 254898 103740 255134
rect 103976 254898 104018 255134
rect 103698 254866 104018 254898
rect 84954 230614 85574 239592
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84699 227492 84765 227493
rect 84699 227428 84700 227492
rect 84764 227428 84765 227492
rect 84699 227427 84765 227428
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 83963 192540 84029 192541
rect 83963 192476 83964 192540
rect 84028 192476 84029 192540
rect 83963 192475 84029 192476
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 176600 81854 190338
rect 84954 176600 85574 194058
rect 91794 237454 92414 239592
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 95514 205174 96134 239592
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 176600 96134 204618
rect 99234 208894 99854 239592
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 97027 177988 97093 177989
rect 97027 177924 97028 177988
rect 97092 177924 97093 177988
rect 97027 177923 97093 177924
rect 97030 175130 97090 177923
rect 98315 176900 98381 176901
rect 98315 176836 98316 176900
rect 98380 176836 98381 176900
rect 98315 176835 98381 176836
rect 96960 175070 97090 175130
rect 98318 175130 98378 176835
rect 99234 176600 99854 208338
rect 102954 212614 103574 239592
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 100707 177580 100773 177581
rect 100707 177516 100708 177580
rect 100772 177516 100773 177580
rect 100707 177515 100773 177516
rect 99419 176492 99485 176493
rect 99419 176428 99420 176492
rect 99484 176428 99485 176492
rect 99419 176427 99485 176428
rect 99422 175130 99482 176427
rect 98318 175070 98380 175130
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 177515
rect 101995 176764 102061 176765
rect 101995 176700 101996 176764
rect 102060 176700 102061 176764
rect 101995 176699 102061 176700
rect 101998 175130 102058 176699
rect 102954 176600 103574 212058
rect 109794 219454 110414 239592
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 104571 177580 104637 177581
rect 104571 177516 104572 177580
rect 104636 177516 104637 177580
rect 104571 177515 104637 177516
rect 105675 177580 105741 177581
rect 105675 177516 105676 177580
rect 105740 177516 105741 177580
rect 105675 177515 105741 177516
rect 106963 177580 107029 177581
rect 106963 177516 106964 177580
rect 107028 177516 107029 177580
rect 106963 177515 107029 177516
rect 103283 176492 103349 176493
rect 103283 176428 103284 176492
rect 103348 176428 103349 176492
rect 103283 176427 103349 176428
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176427
rect 104574 175130 104634 177515
rect 105678 175130 105738 177515
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 105738 175130
rect 106966 175130 107026 177515
rect 108067 177036 108133 177037
rect 108067 176972 108068 177036
rect 108132 176972 108133 177036
rect 108067 176971 108133 176972
rect 108070 175130 108130 176971
rect 109794 176600 110414 182898
rect 113514 223174 114134 239592
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 110643 178260 110709 178261
rect 110643 178196 110644 178260
rect 110708 178196 110709 178260
rect 110643 178195 110709 178196
rect 109539 175404 109605 175405
rect 109539 175340 109540 175404
rect 109604 175340 109605 175404
rect 109539 175339 109605 175340
rect 109542 175130 109602 175339
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109472 175070 109602 175130
rect 110646 175130 110706 178195
rect 113219 177580 113285 177581
rect 113219 177516 113220 177580
rect 113284 177516 113285 177580
rect 113219 177515 113285 177516
rect 112115 177172 112181 177173
rect 112115 177108 112116 177172
rect 112180 177108 112181 177172
rect 112115 177107 112181 177108
rect 112118 175130 112178 177107
rect 113222 175130 113282 177515
rect 113514 176600 114134 186618
rect 117234 226894 117854 239592
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 116899 177580 116965 177581
rect 116899 177516 116900 177580
rect 116964 177516 116965 177580
rect 116899 177515 116965 177516
rect 115795 176764 115861 176765
rect 115795 176700 115796 176764
rect 115860 176700 115861 176764
rect 115795 176699 115861 176700
rect 114323 175676 114389 175677
rect 114323 175612 114324 175676
rect 114388 175612 114389 175676
rect 114323 175611 114389 175612
rect 110646 175070 110756 175130
rect 109472 174494 109532 175070
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 113144 175070 113282 175130
rect 114326 175130 114386 175611
rect 115798 175130 115858 176699
rect 114326 175070 114428 175130
rect 112056 174494 112116 175070
rect 113144 174494 113204 175070
rect 114368 174494 114428 175070
rect 115728 175070 115858 175130
rect 116902 175130 116962 177515
rect 117234 176600 117854 190338
rect 120954 230614 121574 239592
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 119475 177580 119541 177581
rect 119475 177516 119476 177580
rect 119540 177516 119541 177580
rect 119475 177515 119541 177516
rect 120763 177580 120829 177581
rect 120763 177516 120764 177580
rect 120828 177516 120829 177580
rect 120763 177515 120829 177516
rect 118371 177172 118437 177173
rect 118371 177108 118372 177172
rect 118436 177108 118437 177172
rect 118371 177107 118437 177108
rect 118374 175130 118434 177107
rect 119478 175130 119538 177515
rect 120766 175130 120826 177515
rect 120954 176600 121574 194058
rect 127794 237454 128414 239592
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 125731 177580 125797 177581
rect 125731 177516 125732 177580
rect 125796 177516 125797 177580
rect 125731 177515 125797 177516
rect 124443 176764 124509 176765
rect 124443 176700 124444 176764
rect 124508 176700 124509 176764
rect 124443 176699 124509 176700
rect 121867 175540 121933 175541
rect 121867 175476 121868 175540
rect 121932 175476 121933 175540
rect 121867 175475 121933 175476
rect 121870 175130 121930 175475
rect 124446 175130 124506 176699
rect 125734 175130 125794 177515
rect 127019 176764 127085 176765
rect 127019 176700 127020 176764
rect 127084 176700 127085 176764
rect 127019 176699 127085 176700
rect 127022 175130 127082 176699
rect 127794 176600 128414 200898
rect 131514 205174 132134 239592
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 129411 177580 129477 177581
rect 129411 177516 129412 177580
rect 129476 177516 129477 177580
rect 129411 177515 129477 177516
rect 116902 175070 117012 175130
rect 115728 174494 115788 175070
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 119400 175070 119538 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 129414 175130 129474 177515
rect 131514 176600 132134 204618
rect 133094 189957 133154 328475
rect 134418 291454 134738 291486
rect 134418 291218 134460 291454
rect 134696 291218 134738 291454
rect 134418 291134 134738 291218
rect 134418 290898 134460 291134
rect 134696 290898 134738 291134
rect 134418 290866 134738 290898
rect 134418 255454 134738 255486
rect 134418 255218 134460 255454
rect 134696 255218 134738 255454
rect 134418 255134 134738 255218
rect 134418 254898 134460 255134
rect 134696 254898 134738 255134
rect 134418 254866 134738 254898
rect 136038 242045 136098 355403
rect 136035 242044 136101 242045
rect 136035 241980 136036 242044
rect 136100 241980 136101 242044
rect 136035 241979 136101 241980
rect 135234 208894 135854 239592
rect 137142 237285 137202 388723
rect 138059 366348 138125 366349
rect 138059 366284 138060 366348
rect 138124 366284 138125 366348
rect 138059 366283 138125 366284
rect 138062 242045 138122 366283
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 329592 139574 356058
rect 139715 349892 139781 349893
rect 139715 349828 139716 349892
rect 139780 349828 139781 349892
rect 139715 349827 139781 349828
rect 138059 242044 138125 242045
rect 138059 241980 138060 242044
rect 138124 241980 138125 242044
rect 138059 241979 138125 241980
rect 137139 237284 137205 237285
rect 137139 237220 137140 237284
rect 137204 237220 137205 237284
rect 137139 237219 137205 237220
rect 137142 237013 137202 237219
rect 137139 237012 137205 237013
rect 137139 236948 137140 237012
rect 137204 236948 137205 237012
rect 137139 236947 137205 236948
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 133091 189956 133157 189957
rect 133091 189892 133092 189956
rect 133156 189892 133157 189956
rect 133091 189891 133157 189892
rect 132355 176764 132421 176765
rect 132355 176700 132356 176764
rect 132420 176700 132421 176764
rect 132355 176699 132421 176700
rect 134379 176764 134445 176765
rect 134379 176700 134380 176764
rect 134444 176700 134445 176764
rect 134379 176699 134445 176700
rect 130699 175812 130765 175813
rect 130699 175748 130700 175812
rect 130764 175748 130765 175812
rect 130699 175747 130765 175748
rect 130702 175130 130762 175747
rect 132358 175130 132418 176699
rect 134382 175130 134442 176699
rect 135234 176600 135854 208338
rect 138954 212614 139574 239592
rect 139718 234021 139778 349827
rect 139715 234020 139781 234021
rect 139715 233956 139716 234020
rect 139780 233956 139781 234020
rect 139715 233955 139781 233956
rect 140822 224773 140882 401643
rect 143395 327044 143461 327045
rect 143395 326980 143396 327044
rect 143460 326980 143461 327044
rect 143395 326979 143461 326980
rect 140819 224772 140885 224773
rect 140819 224708 140820 224772
rect 140884 224708 140885 224772
rect 140819 224707 140885 224708
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 136035 176764 136101 176765
rect 136035 176700 136036 176764
rect 136100 176700 136101 176764
rect 136035 176699 136101 176700
rect 136038 175130 136098 176699
rect 138954 176600 139574 212058
rect 143398 189821 143458 326979
rect 143582 232933 143642 442307
rect 145794 435454 146414 470898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 148179 455564 148245 455565
rect 148179 455500 148180 455564
rect 148244 455500 148245 455564
rect 148179 455499 148245 455500
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 329592 146414 362898
rect 148182 241501 148242 455499
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 151859 355604 151925 355605
rect 151859 355540 151860 355604
rect 151924 355540 151925 355604
rect 151859 355539 151925 355540
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 329592 150134 330618
rect 150387 327588 150453 327589
rect 150387 327524 150388 327588
rect 150452 327524 150453 327588
rect 150387 327523 150453 327524
rect 149778 309454 150098 309486
rect 149778 309218 149820 309454
rect 150056 309218 150098 309454
rect 149778 309134 150098 309218
rect 149778 308898 149820 309134
rect 150056 308898 150098 309134
rect 149778 308866 150098 308898
rect 149778 273454 150098 273486
rect 149778 273218 149820 273454
rect 150056 273218 150098 273454
rect 149778 273134 150098 273218
rect 149778 272898 149820 273134
rect 150056 272898 150098 273134
rect 149778 272866 150098 272898
rect 148179 241500 148245 241501
rect 148179 241436 148180 241500
rect 148244 241436 148245 241500
rect 148179 241435 148245 241436
rect 143579 232932 143645 232933
rect 143579 232868 143580 232932
rect 143644 232868 143645 232932
rect 143579 232867 143645 232868
rect 145794 219454 146414 239592
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 143395 189820 143461 189821
rect 143395 189756 143396 189820
rect 143460 189756 143461 189820
rect 143395 189755 143461 189756
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 149514 223174 150134 239592
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 150390 197981 150450 327523
rect 151862 241909 151922 355539
rect 153234 334894 153854 370338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 159219 586532 159285 586533
rect 159219 586468 159220 586532
rect 159284 586468 159285 586532
rect 159219 586467 159285 586468
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156459 360908 156525 360909
rect 156459 360844 156460 360908
rect 156524 360844 156525 360908
rect 156459 360843 156525 360844
rect 155171 341188 155237 341189
rect 155171 341124 155172 341188
rect 155236 341124 155237 341188
rect 155171 341123 155237 341124
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 329592 153854 334338
rect 154067 330172 154133 330173
rect 154067 330108 154068 330172
rect 154132 330108 154133 330172
rect 154067 330107 154133 330108
rect 154070 324730 154130 330107
rect 154251 327724 154317 327725
rect 154251 327660 154252 327724
rect 154316 327660 154317 327724
rect 154251 327659 154317 327660
rect 154254 325277 154314 327659
rect 154251 325276 154317 325277
rect 154251 325212 154252 325276
rect 154316 325212 154317 325276
rect 154251 325211 154317 325212
rect 154070 324670 154314 324730
rect 154254 323645 154314 324670
rect 154251 323644 154317 323645
rect 154251 323580 154252 323644
rect 154316 323580 154317 323644
rect 154251 323579 154317 323580
rect 155174 320789 155234 341123
rect 155723 327588 155789 327589
rect 155723 327524 155724 327588
rect 155788 327524 155789 327588
rect 155723 327523 155789 327524
rect 155726 325005 155786 327523
rect 155723 325004 155789 325005
rect 155723 324940 155724 325004
rect 155788 324940 155789 325004
rect 155723 324939 155789 324940
rect 155171 320788 155237 320789
rect 155171 320724 155172 320788
rect 155236 320724 155237 320788
rect 155171 320723 155237 320724
rect 156462 318749 156522 360843
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156459 318748 156525 318749
rect 156459 318684 156460 318748
rect 156524 318684 156525 318748
rect 156459 318683 156525 318684
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 154619 260812 154685 260813
rect 154619 260748 154620 260812
rect 154684 260748 154685 260812
rect 154619 260747 154685 260748
rect 154251 244628 154317 244629
rect 154251 244564 154252 244628
rect 154316 244564 154317 244628
rect 154251 244563 154317 244564
rect 151859 241908 151925 241909
rect 151859 241844 151860 241908
rect 151924 241844 151925 241908
rect 151859 241843 151925 241844
rect 153234 226894 153854 239592
rect 154254 238770 154314 244563
rect 154070 238710 154314 238770
rect 154070 230349 154130 238710
rect 154622 231437 154682 260747
rect 155171 243540 155237 243541
rect 155171 243476 155172 243540
rect 155236 243476 155237 243540
rect 155171 243475 155237 243476
rect 154619 231436 154685 231437
rect 154619 231372 154620 231436
rect 154684 231372 154685 231436
rect 154619 231371 154685 231372
rect 154067 230348 154133 230349
rect 154067 230284 154068 230348
rect 154132 230284 154133 230348
rect 154067 230283 154133 230284
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 150387 197980 150453 197981
rect 150387 197916 150388 197980
rect 150452 197916 150453 197980
rect 150387 197915 150453 197916
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 148179 177580 148245 177581
rect 148179 177516 148180 177580
rect 148244 177516 148245 177580
rect 148179 177515 148245 177516
rect 129414 175070 129524 175130
rect 118312 174494 118372 175070
rect 119400 174494 119460 175070
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123069 174996 123135 174997
rect 123069 174932 123070 174996
rect 123134 174932 123135 174996
rect 123069 174931 123135 174932
rect 123072 174494 123132 174931
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128101 174860 128167 174861
rect 128101 174796 128102 174860
rect 128166 174796 128167 174860
rect 128101 174795 128167 174796
rect 128104 174494 128164 174795
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 132048 175070 132418 175130
rect 133136 175070 133338 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 133278 174725 133338 175070
rect 134360 175070 134442 175130
rect 135720 175070 136098 175130
rect 148182 175130 148242 177515
rect 149514 176600 150134 186618
rect 153234 190894 153854 226338
rect 154622 206277 154682 231371
rect 155174 228989 155234 243475
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 155171 228988 155237 228989
rect 155171 228924 155172 228988
rect 155236 228924 155237 228988
rect 155171 228923 155237 228924
rect 154619 206276 154685 206277
rect 154619 206212 154620 206276
rect 154684 206212 154685 206276
rect 154619 206211 154685 206212
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 176600 153854 190338
rect 156954 194614 157574 230058
rect 159222 197981 159282 586467
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 160691 448628 160757 448629
rect 160691 448564 160692 448628
rect 160756 448564 160757 448628
rect 160691 448563 160757 448564
rect 160694 303789 160754 448563
rect 163794 417454 164414 452898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 165659 441692 165725 441693
rect 165659 441628 165660 441692
rect 165724 441628 165725 441692
rect 165659 441627 165725 441628
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 161979 323236 162045 323237
rect 161979 323172 161980 323236
rect 162044 323172 162045 323236
rect 161979 323171 162045 323172
rect 160691 303788 160757 303789
rect 160691 303724 160692 303788
rect 160756 303724 160757 303788
rect 160691 303723 160757 303724
rect 161982 302837 162042 323171
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 161979 302836 162045 302837
rect 161979 302772 161980 302836
rect 162044 302772 162045 302836
rect 161979 302771 162045 302772
rect 161979 293588 162045 293589
rect 161979 293524 161980 293588
rect 162044 293524 162045 293588
rect 161979 293523 162045 293524
rect 161982 206277 162042 293523
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 161979 206276 162045 206277
rect 161979 206212 161980 206276
rect 162044 206212 162045 206276
rect 161979 206211 162045 206212
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 159219 197980 159285 197981
rect 159219 197916 159220 197980
rect 159284 197916 159285 197980
rect 159219 197915 159285 197916
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 176600 157574 194058
rect 158851 176764 158917 176765
rect 158851 176700 158852 176764
rect 158916 176700 158917 176764
rect 158851 176699 158917 176700
rect 158854 175130 158914 176699
rect 163794 176600 164414 200898
rect 164739 175676 164805 175677
rect 164739 175612 164740 175676
rect 164804 175612 164805 175676
rect 164739 175611 164805 175612
rect 148182 175070 148292 175130
rect 133275 174724 133341 174725
rect 133275 174660 133276 174724
rect 133340 174660 133341 174724
rect 133275 174659 133341 174660
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 69072 165454 69420 165486
rect 69072 165218 69128 165454
rect 69364 165218 69420 165454
rect 69072 165134 69420 165218
rect 69072 164898 69128 165134
rect 69364 164898 69420 165134
rect 69072 164866 69420 164898
rect 164136 165454 164484 165486
rect 164136 165218 164192 165454
rect 164428 165218 164484 165454
rect 164136 165134 164484 165218
rect 164136 164898 164192 165134
rect 164428 164898 164484 165134
rect 164136 164866 164484 164898
rect 164742 164389 164802 175611
rect 164739 164388 164805 164389
rect 164739 164324 164740 164388
rect 164804 164324 164805 164388
rect 164739 164323 164805 164324
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 69072 129454 69420 129486
rect 69072 129218 69128 129454
rect 69364 129218 69420 129454
rect 69072 129134 69420 129218
rect 69072 128898 69128 129134
rect 69364 128898 69420 129134
rect 69072 128866 69420 128898
rect 164136 129454 164484 129486
rect 164136 129218 164192 129454
rect 164428 129218 164484 129454
rect 164136 129134 164484 129218
rect 164136 128898 164192 129134
rect 164428 128898 164484 129134
rect 164136 128866 164484 128898
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 85536 94890 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 85536 94830 85866 94890
rect 86624 94830 86786 94890
rect 87984 94830 88074 94890
rect 73794 75454 74414 93100
rect 74766 91221 74826 94830
rect 74763 91220 74829 91221
rect 74763 91156 74764 91220
rect 74828 91156 74829 91220
rect 74763 91155 74829 91156
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 67771 19956 67837 19957
rect 67771 19892 67772 19956
rect 67836 19892 67837 19956
rect 67771 19891 67837 19892
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 93100
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 93100
rect 84334 91765 84394 94830
rect 84331 91764 84397 91765
rect 84331 91700 84332 91764
rect 84396 91700 84397 91764
rect 84331 91699 84397 91700
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 93100
rect 85806 91221 85866 94830
rect 86726 92445 86786 94830
rect 86723 92444 86789 92445
rect 86723 92380 86724 92444
rect 86788 92380 86789 92444
rect 86723 92379 86789 92380
rect 88014 91221 88074 94830
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 88934 92445 88994 94830
rect 88931 92444 88997 92445
rect 88931 92380 88932 92444
rect 88996 92380 88997 92444
rect 88931 92379 88997 92380
rect 90222 91221 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 94920 94890 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 94920 94830 95066 94890
rect 96008 94830 96354 94890
rect 91326 91221 91386 94830
rect 85803 91220 85869 91221
rect 85803 91156 85804 91220
rect 85868 91156 85869 91220
rect 85803 91155 85869 91156
rect 88011 91220 88077 91221
rect 88011 91156 88012 91220
rect 88076 91156 88077 91220
rect 88011 91155 88077 91156
rect 90219 91220 90285 91221
rect 90219 91156 90220 91220
rect 90284 91156 90285 91220
rect 90219 91155 90285 91156
rect 91323 91220 91389 91221
rect 91323 91156 91324 91220
rect 91388 91156 91389 91220
rect 91323 91155 91389 91156
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 93100
rect 92614 91221 92674 94830
rect 93902 91357 93962 94830
rect 93899 91356 93965 91357
rect 93899 91292 93900 91356
rect 93964 91292 93965 91356
rect 93899 91291 93965 91292
rect 95006 91221 95066 94830
rect 92611 91220 92677 91221
rect 92611 91156 92612 91220
rect 92676 91156 92677 91220
rect 92611 91155 92677 91156
rect 95003 91220 95069 91221
rect 95003 91156 95004 91220
rect 95068 91156 95069 91220
rect 95003 91155 95069 91156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 93100
rect 96294 91221 96354 94830
rect 96662 94830 96748 94890
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 99544 94890 99604 95200
rect 100632 94890 100692 95200
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 99136 94830 99298 94890
rect 99544 94830 99666 94890
rect 96662 93941 96722 94830
rect 96659 93940 96725 93941
rect 96659 93876 96660 93940
rect 96724 93876 96725 93940
rect 96659 93875 96725 93876
rect 97214 91221 97274 94830
rect 98134 91221 98194 94830
rect 98502 91493 98562 94830
rect 99238 93805 99298 94830
rect 99235 93804 99301 93805
rect 99235 93740 99236 93804
rect 99300 93740 99301 93804
rect 99235 93739 99301 93740
rect 99606 93669 99666 94830
rect 100526 94830 100692 94890
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 100954 94890
rect 99603 93668 99669 93669
rect 99603 93604 99604 93668
rect 99668 93604 99669 93668
rect 99603 93603 99669 93604
rect 98499 91492 98565 91493
rect 98499 91428 98500 91492
rect 98564 91428 98565 91492
rect 98499 91427 98565 91428
rect 96291 91220 96357 91221
rect 96291 91156 96292 91220
rect 96356 91156 96357 91220
rect 96291 91155 96357 91156
rect 97211 91220 97277 91221
rect 97211 91156 97212 91220
rect 97276 91156 97277 91220
rect 97211 91155 97277 91156
rect 98131 91220 98197 91221
rect 98131 91156 98132 91220
rect 98196 91156 98197 91220
rect 98131 91155 98197 91156
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 93100
rect 100526 91221 100586 94830
rect 100894 91221 100954 94830
rect 101814 94830 101916 94890
rect 101992 94890 102052 95200
rect 102944 94890 103004 95200
rect 103216 94890 103276 95200
rect 104304 94890 104364 95200
rect 101992 94830 102058 94890
rect 101814 91357 101874 94830
rect 101998 91493 102058 94830
rect 102550 94830 103004 94890
rect 103102 94830 103276 94890
rect 104206 94830 104364 94890
rect 104440 94890 104500 95200
rect 105392 94890 105452 95200
rect 105664 94890 105724 95200
rect 106480 94890 106540 95200
rect 104440 94830 104634 94890
rect 105392 94830 105554 94890
rect 105664 94830 105738 94890
rect 101995 91492 102061 91493
rect 101995 91428 101996 91492
rect 102060 91428 102061 91492
rect 101995 91427 102061 91428
rect 101811 91356 101877 91357
rect 101811 91292 101812 91356
rect 101876 91292 101877 91356
rect 101811 91291 101877 91292
rect 102550 91221 102610 94830
rect 103102 93870 103162 94830
rect 102734 93810 103162 93870
rect 102734 91221 102794 93810
rect 100523 91220 100589 91221
rect 100523 91156 100524 91220
rect 100588 91156 100589 91220
rect 100523 91155 100589 91156
rect 100891 91220 100957 91221
rect 100891 91156 100892 91220
rect 100956 91156 100957 91220
rect 100891 91155 100957 91156
rect 102547 91220 102613 91221
rect 102547 91156 102548 91220
rect 102612 91156 102613 91220
rect 102547 91155 102613 91156
rect 102731 91220 102797 91221
rect 102731 91156 102732 91220
rect 102796 91156 102797 91220
rect 102731 91155 102797 91156
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 93100
rect 104206 91221 104266 94830
rect 104574 91221 104634 94830
rect 105494 91221 105554 94830
rect 105678 91901 105738 94830
rect 106414 94830 106540 94890
rect 106616 94890 106676 95200
rect 107704 94890 107764 95200
rect 108112 94890 108172 95200
rect 106616 94830 106842 94890
rect 105675 91900 105741 91901
rect 105675 91836 105676 91900
rect 105740 91836 105741 91900
rect 105675 91835 105741 91836
rect 106414 91765 106474 94830
rect 106411 91764 106477 91765
rect 106411 91700 106412 91764
rect 106476 91700 106477 91764
rect 106411 91699 106477 91700
rect 106782 91629 106842 94830
rect 107702 94830 107764 94890
rect 108070 94830 108172 94890
rect 109064 94890 109124 95200
rect 109472 94890 109532 95200
rect 110152 94890 110212 95200
rect 110696 94890 110756 95200
rect 111240 94890 111300 95200
rect 109064 94830 109234 94890
rect 109472 94830 109602 94890
rect 106779 91628 106845 91629
rect 106779 91564 106780 91628
rect 106844 91564 106845 91628
rect 106779 91563 106845 91564
rect 107702 91357 107762 94830
rect 107699 91356 107765 91357
rect 107699 91292 107700 91356
rect 107764 91292 107765 91356
rect 107699 91291 107765 91292
rect 108070 91221 108130 94830
rect 109174 92445 109234 94830
rect 109171 92444 109237 92445
rect 109171 92380 109172 92444
rect 109236 92380 109237 92444
rect 109171 92379 109237 92380
rect 109542 91221 109602 94830
rect 110094 94830 110212 94890
rect 110646 94830 110756 94890
rect 111198 94830 111300 94890
rect 111920 94890 111980 95200
rect 112328 94890 112388 95200
rect 113144 95029 113204 95200
rect 113141 95028 113207 95029
rect 113141 94964 113142 95028
rect 113206 94964 113207 95028
rect 113141 94963 113207 94964
rect 113688 94890 113748 95200
rect 114368 94890 114428 95200
rect 114507 95028 114573 95029
rect 114507 94964 114508 95028
rect 114572 94964 114573 95028
rect 114507 94963 114573 94964
rect 111920 94830 111994 94890
rect 110094 93261 110154 94830
rect 110091 93260 110157 93261
rect 110091 93196 110092 93260
rect 110156 93196 110157 93260
rect 110091 93195 110157 93196
rect 104203 91220 104269 91221
rect 104203 91156 104204 91220
rect 104268 91156 104269 91220
rect 104203 91155 104269 91156
rect 104571 91220 104637 91221
rect 104571 91156 104572 91220
rect 104636 91156 104637 91220
rect 104571 91155 104637 91156
rect 105491 91220 105557 91221
rect 105491 91156 105492 91220
rect 105556 91156 105557 91220
rect 105491 91155 105557 91156
rect 108067 91220 108133 91221
rect 108067 91156 108068 91220
rect 108132 91156 108133 91220
rect 108067 91155 108133 91156
rect 109539 91220 109605 91221
rect 109539 91156 109540 91220
rect 109604 91156 109605 91220
rect 109539 91155 109605 91156
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 93100
rect 110646 91221 110706 94830
rect 111198 92445 111258 94830
rect 111195 92444 111261 92445
rect 111195 92380 111196 92444
rect 111260 92380 111261 92444
rect 111195 92379 111261 92380
rect 111934 91221 111994 94830
rect 112302 94830 112388 94890
rect 113222 94830 113748 94890
rect 114326 94830 114428 94890
rect 112302 91221 112362 94830
rect 113222 91221 113282 94830
rect 110643 91220 110709 91221
rect 110643 91156 110644 91220
rect 110708 91156 110709 91220
rect 110643 91155 110709 91156
rect 111931 91220 111997 91221
rect 111931 91156 111932 91220
rect 111996 91156 111997 91220
rect 111931 91155 111997 91156
rect 112299 91220 112365 91221
rect 112299 91156 112300 91220
rect 112364 91156 112365 91220
rect 112299 91155 112365 91156
rect 113219 91220 113285 91221
rect 113219 91156 113220 91220
rect 113284 91156 113285 91220
rect 113219 91155 113285 91156
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 79174 114134 93100
rect 114326 91221 114386 94830
rect 114510 92445 114570 94963
rect 114776 94890 114836 95200
rect 115456 94890 115516 95200
rect 115864 94890 115924 95200
rect 114776 94830 114938 94890
rect 114507 92444 114573 92445
rect 114507 92380 114508 92444
rect 114572 92380 114573 92444
rect 114507 92379 114573 92380
rect 114878 91765 114938 94830
rect 115430 94830 115516 94890
rect 115798 94830 115924 94890
rect 116680 94890 116740 95200
rect 117088 94890 117148 95200
rect 116680 94830 116778 94890
rect 114875 91764 114941 91765
rect 114875 91700 114876 91764
rect 114940 91700 114941 91764
rect 114875 91699 114941 91700
rect 115430 91357 115490 94830
rect 115427 91356 115493 91357
rect 115427 91292 115428 91356
rect 115492 91292 115493 91356
rect 115427 91291 115493 91292
rect 115798 91221 115858 94830
rect 116718 91765 116778 94830
rect 117086 94830 117148 94890
rect 117904 94890 117964 95200
rect 118176 94890 118236 95200
rect 119400 94890 119460 95200
rect 117904 94830 118066 94890
rect 118176 94830 118250 94890
rect 116715 91764 116781 91765
rect 116715 91700 116716 91764
rect 116780 91700 116781 91764
rect 116715 91699 116781 91700
rect 117086 91221 117146 94830
rect 114323 91220 114389 91221
rect 114323 91156 114324 91220
rect 114388 91156 114389 91220
rect 114323 91155 114389 91156
rect 115795 91220 115861 91221
rect 115795 91156 115796 91220
rect 115860 91156 115861 91220
rect 115795 91155 115861 91156
rect 117083 91220 117149 91221
rect 117083 91156 117084 91220
rect 117148 91156 117149 91220
rect 117083 91155 117149 91156
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 82894 117854 93100
rect 118006 91357 118066 94830
rect 118003 91356 118069 91357
rect 118003 91292 118004 91356
rect 118068 91292 118069 91356
rect 118003 91291 118069 91292
rect 118190 91221 118250 94830
rect 119294 94830 119460 94890
rect 119536 94890 119596 95200
rect 120216 94890 120276 95200
rect 120624 94890 120684 95200
rect 121712 94890 121772 95200
rect 119536 94830 119722 94890
rect 119294 91221 119354 94830
rect 119662 93533 119722 94830
rect 120214 94830 120276 94890
rect 120582 94830 120684 94890
rect 121686 94830 121772 94890
rect 121984 94890 122044 95200
rect 122800 94890 122860 95200
rect 123208 94890 123268 95200
rect 121984 94830 122114 94890
rect 122800 94830 123034 94890
rect 119659 93532 119725 93533
rect 119659 93468 119660 93532
rect 119724 93468 119725 93532
rect 119659 93467 119725 93468
rect 120214 92173 120274 94830
rect 120211 92172 120277 92173
rect 120211 92108 120212 92172
rect 120276 92108 120277 92172
rect 120211 92107 120277 92108
rect 120582 91221 120642 94830
rect 121686 93533 121746 94830
rect 121683 93532 121749 93533
rect 121683 93468 121684 93532
rect 121748 93468 121749 93532
rect 121683 93467 121749 93468
rect 118187 91220 118253 91221
rect 118187 91156 118188 91220
rect 118252 91156 118253 91220
rect 118187 91155 118253 91156
rect 119291 91220 119357 91221
rect 119291 91156 119292 91220
rect 119356 91156 119357 91220
rect 119291 91155 119357 91156
rect 120579 91220 120645 91221
rect 120579 91156 120580 91220
rect 120644 91156 120645 91220
rect 120579 91155 120645 91156
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 86614 121574 93100
rect 122054 91221 122114 94830
rect 122974 93870 123034 94830
rect 122606 93810 123034 93870
rect 123158 94830 123268 94890
rect 122606 91490 122666 93810
rect 122606 91430 122850 91490
rect 122790 91357 122850 91430
rect 122787 91356 122853 91357
rect 122787 91292 122788 91356
rect 122852 91292 122853 91356
rect 122787 91291 122853 91292
rect 123158 91221 123218 94830
rect 124024 94757 124084 95200
rect 124432 94890 124492 95200
rect 125384 94890 125444 95200
rect 124432 94830 124506 94890
rect 124021 94756 124087 94757
rect 124021 94692 124022 94756
rect 124086 94692 124087 94756
rect 124021 94691 124087 94692
rect 124446 91221 124506 94830
rect 125366 94830 125444 94890
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125794 94890
rect 125366 91357 125426 94830
rect 125734 91629 125794 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 126608 94830 126714 94890
rect 125731 91628 125797 91629
rect 125731 91564 125732 91628
rect 125796 91564 125797 91628
rect 125731 91563 125797 91564
rect 126470 91357 126530 94830
rect 125363 91356 125429 91357
rect 125363 91292 125364 91356
rect 125428 91292 125429 91356
rect 125363 91291 125429 91292
rect 126467 91356 126533 91357
rect 126467 91292 126468 91356
rect 126532 91292 126533 91356
rect 126467 91291 126533 91292
rect 126654 91221 126714 94830
rect 127574 94830 128164 94890
rect 129328 94890 129388 95200
rect 130688 94890 130748 95200
rect 131912 94890 131972 95200
rect 133136 94890 133196 95200
rect 129328 94830 129474 94890
rect 130688 94830 130762 94890
rect 131912 94830 132050 94890
rect 127574 91221 127634 94830
rect 122051 91220 122117 91221
rect 122051 91156 122052 91220
rect 122116 91156 122117 91220
rect 122051 91155 122117 91156
rect 123155 91220 123221 91221
rect 123155 91156 123156 91220
rect 123220 91156 123221 91220
rect 123155 91155 123221 91156
rect 124443 91220 124509 91221
rect 124443 91156 124444 91220
rect 124508 91156 124509 91220
rect 124443 91155 124509 91156
rect 126651 91220 126717 91221
rect 126651 91156 126652 91220
rect 126716 91156 126717 91220
rect 126651 91155 126717 91156
rect 127571 91220 127637 91221
rect 127571 91156 127572 91220
rect 127636 91156 127637 91220
rect 127571 91155 127637 91156
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 93100
rect 129414 91221 129474 94830
rect 130702 92037 130762 94830
rect 131990 94077 132050 94830
rect 133094 94830 133196 94890
rect 134360 94890 134420 95200
rect 135584 94890 135644 95200
rect 151307 95028 151373 95029
rect 151307 94964 151308 95028
rect 151372 94964 151373 95028
rect 151307 94963 151373 94964
rect 134360 94830 134442 94890
rect 135584 94830 136098 94890
rect 131987 94076 132053 94077
rect 131987 94012 131988 94076
rect 132052 94012 132053 94076
rect 131987 94011 132053 94012
rect 130699 92036 130765 92037
rect 130699 91972 130700 92036
rect 130764 91972 130765 92036
rect 130699 91971 130765 91972
rect 129411 91220 129477 91221
rect 129411 91156 129412 91220
rect 129476 91156 129477 91220
rect 129411 91155 129477 91156
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 61174 132134 93100
rect 133094 91221 133154 94830
rect 134382 91221 134442 94830
rect 133091 91220 133157 91221
rect 133091 91156 133092 91220
rect 133156 91156 133157 91220
rect 133091 91155 133157 91156
rect 134379 91220 134445 91221
rect 134379 91156 134380 91220
rect 134444 91156 134445 91220
rect 134379 91155 134445 91156
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 64894 135854 93100
rect 136038 92445 136098 94830
rect 136035 92444 136101 92445
rect 136035 92380 136036 92444
rect 136100 92380 136101 92444
rect 136035 92379 136101 92380
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 93100
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 79174 150134 93100
rect 151310 92445 151370 94963
rect 151496 94890 151556 95200
rect 151494 94830 151556 94890
rect 151632 94890 151692 95200
rect 151768 95029 151828 95200
rect 151765 95028 151831 95029
rect 151765 94964 151766 95028
rect 151830 94964 151831 95028
rect 151765 94963 151831 94964
rect 151904 94890 151964 95200
rect 151632 94830 151738 94890
rect 151307 92444 151373 92445
rect 151307 92380 151308 92444
rect 151372 92380 151373 92444
rect 151307 92379 151373 92380
rect 151494 91221 151554 94830
rect 151678 91357 151738 94830
rect 151862 94830 151964 94890
rect 151675 91356 151741 91357
rect 151675 91292 151676 91356
rect 151740 91292 151741 91356
rect 151675 91291 151741 91292
rect 151862 91221 151922 94830
rect 151491 91220 151557 91221
rect 151491 91156 151492 91220
rect 151556 91156 151557 91220
rect 151491 91155 151557 91156
rect 151859 91220 151925 91221
rect 151859 91156 151860 91220
rect 151924 91156 151925 91220
rect 151859 91155 151925 91156
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 82894 153854 93100
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 86614 157574 93100
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 93100
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 165662 10301 165722 441627
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 172467 449988 172533 449989
rect 172467 449924 172468 449988
rect 172532 449924 172533 449988
rect 172467 449923 172533 449924
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 170259 320380 170325 320381
rect 170259 320316 170260 320380
rect 170324 320316 170325 320380
rect 170259 320315 170325 320316
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 168419 197980 168485 197981
rect 168419 197916 168420 197980
rect 168484 197916 168485 197980
rect 168419 197915 168485 197916
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 166211 97204 166277 97205
rect 166211 97140 166212 97204
rect 166276 97140 166277 97204
rect 166211 97139 166277 97140
rect 167514 97174 168134 132618
rect 166214 84013 166274 97139
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 166211 84012 166277 84013
rect 166211 83948 166212 84012
rect 166276 83948 166277 84012
rect 166211 83947 166277 83948
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 165659 10300 165725 10301
rect 165659 10236 165660 10300
rect 165724 10236 165725 10300
rect 165659 10235 165725 10236
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 -3226 168134 24618
rect 168422 4861 168482 197915
rect 170262 8941 170322 320315
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 172470 241773 172530 449923
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 184059 364580 184125 364581
rect 184059 364516 184060 364580
rect 184124 364516 184125 364580
rect 184059 364515 184125 364516
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 180011 296036 180077 296037
rect 180011 295972 180012 296036
rect 180076 295972 180077 296036
rect 180011 295971 180077 295972
rect 178539 292636 178605 292637
rect 178539 292572 178540 292636
rect 178604 292572 178605 292636
rect 178539 292571 178605 292572
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 172467 241772 172533 241773
rect 172467 241708 172468 241772
rect 172532 241708 172533 241772
rect 172467 241707 172533 241708
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 170259 8940 170325 8941
rect 170259 8876 170260 8940
rect 170324 8876 170325 8940
rect 170259 8875 170325 8876
rect 168419 4860 168485 4861
rect 168419 4796 168420 4860
rect 168484 4796 168485 4860
rect 168419 4795 168485 4796
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 212614 175574 248058
rect 178542 216477 178602 292571
rect 180014 237285 180074 295971
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 180011 237284 180077 237285
rect 180011 237220 180012 237284
rect 180076 237220 180077 237284
rect 180011 237219 180077 237220
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 178539 216476 178605 216477
rect 178539 216412 178540 216476
rect 178604 216412 178605 216476
rect 178539 216411 178605 216412
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 184062 142765 184122 364515
rect 185514 331174 186134 366618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 188291 349212 188357 349213
rect 188291 349148 188292 349212
rect 188356 349148 188357 349212
rect 188291 349147 188357 349148
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 186819 301068 186885 301069
rect 186819 301004 186820 301068
rect 186884 301004 186885 301068
rect 186819 301003 186885 301004
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 186267 236604 186333 236605
rect 186267 236540 186268 236604
rect 186332 236540 186333 236604
rect 186267 236539 186333 236540
rect 186270 235653 186330 236539
rect 186267 235652 186333 235653
rect 186267 235588 186268 235652
rect 186332 235588 186333 235652
rect 186267 235587 186333 235588
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 184059 142764 184125 142765
rect 184059 142700 184060 142764
rect 184124 142700 184125 142764
rect 184059 142699 184125 142700
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 186822 14517 186882 301003
rect 188294 192677 188354 349147
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203011 345676 203077 345677
rect 203011 345612 203012 345676
rect 203076 345612 203077 345676
rect 203011 345611 203077 345612
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 203014 345133 203074 345611
rect 203011 345132 203077 345133
rect 203011 345068 203012 345132
rect 203076 345068 203077 345132
rect 203011 345067 203077 345068
rect 196571 330308 196637 330309
rect 196571 330244 196572 330308
rect 196636 330244 196637 330308
rect 196571 330243 196637 330244
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 191051 287332 191117 287333
rect 191051 287268 191052 287332
rect 191116 287268 191117 287332
rect 191051 287267 191117 287268
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 188291 192676 188357 192677
rect 188291 192612 188292 192676
rect 188356 192612 188357 192676
rect 188291 192611 188357 192612
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 186819 14516 186885 14517
rect 186819 14452 186820 14516
rect 186884 14452 186885 14516
rect 186819 14451 186885 14452
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 191054 10301 191114 287267
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 195835 241500 195901 241501
rect 195835 241436 195836 241500
rect 195900 241436 195901 241500
rect 195835 241435 195901 241436
rect 195838 240685 195898 241435
rect 195835 240684 195901 240685
rect 195835 240620 195836 240684
rect 195900 240620 195901 240684
rect 195835 240619 195901 240620
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 195838 229805 195898 240619
rect 195835 229804 195901 229805
rect 195835 229740 195836 229804
rect 195900 229740 195901 229804
rect 195835 229739 195901 229740
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 196574 97205 196634 330243
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 286182 200414 308898
rect 197307 284748 197373 284749
rect 197307 284684 197308 284748
rect 197372 284684 197373 284748
rect 197307 284683 197373 284684
rect 197310 280941 197370 284683
rect 197307 280940 197373 280941
rect 197307 280876 197308 280940
rect 197372 280876 197373 280940
rect 197307 280875 197373 280876
rect 197123 267204 197189 267205
rect 197123 267140 197124 267204
rect 197188 267140 197189 267204
rect 197123 267139 197189 267140
rect 197126 231573 197186 267139
rect 199883 265300 199949 265301
rect 199883 265236 199884 265300
rect 199948 265236 199949 265300
rect 199883 265235 199949 265236
rect 199515 248436 199581 248437
rect 199515 248372 199516 248436
rect 199580 248372 199581 248436
rect 199515 248371 199581 248372
rect 197123 231572 197189 231573
rect 197123 231508 197124 231572
rect 197188 231508 197189 231572
rect 197123 231507 197189 231508
rect 199518 223005 199578 248371
rect 199886 240277 199946 265235
rect 200067 248436 200133 248437
rect 200067 248372 200068 248436
rect 200132 248372 200133 248436
rect 200067 248371 200133 248372
rect 200070 247621 200130 248371
rect 200067 247620 200133 247621
rect 200067 247556 200068 247620
rect 200132 247556 200133 247620
rect 200067 247555 200133 247556
rect 199883 240276 199949 240277
rect 199883 240212 199884 240276
rect 199948 240212 199949 240276
rect 199883 240211 199949 240212
rect 203014 238645 203074 345067
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 286182 204134 312618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 207979 365804 208045 365805
rect 207979 365740 207980 365804
rect 208044 365740 208045 365804
rect 207979 365739 208045 365740
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 286182 207854 316338
rect 205403 283932 205469 283933
rect 205403 283868 205404 283932
rect 205468 283868 205469 283932
rect 205403 283867 205469 283868
rect 204408 255454 204728 255486
rect 204408 255218 204450 255454
rect 204686 255218 204728 255454
rect 204408 255134 204728 255218
rect 204408 254898 204450 255134
rect 204686 254898 204728 255134
rect 204408 254866 204728 254898
rect 203011 238644 203077 238645
rect 203011 238580 203012 238644
rect 203076 238580 203077 238644
rect 203011 238579 203077 238580
rect 199794 237454 200414 238182
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199515 223004 199581 223005
rect 199515 222940 199516 223004
rect 199580 222940 199581 223004
rect 199515 222939 199581 222940
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 196571 97204 196637 97205
rect 196571 97140 196572 97204
rect 196636 97140 196637 97204
rect 196571 97139 196637 97140
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 191051 10300 191117 10301
rect 191051 10236 191052 10300
rect 191116 10236 191117 10300
rect 191051 10235 191117 10236
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 205174 204134 238182
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 205406 93669 205466 283867
rect 207234 208894 207854 238182
rect 207982 237285 208042 365739
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 212579 339692 212645 339693
rect 212579 339628 212580 339692
rect 212644 339628 212645 339692
rect 212579 339627 212645 339628
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 286182 211574 320058
rect 212395 283932 212461 283933
rect 212395 283868 212396 283932
rect 212460 283868 212461 283932
rect 212395 283867 212461 283868
rect 207979 237284 208045 237285
rect 207979 237220 207980 237284
rect 208044 237220 208045 237284
rect 207979 237219 208045 237220
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 205403 93668 205469 93669
rect 205403 93604 205404 93668
rect 205468 93604 205469 93668
rect 205403 93603 205469 93604
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 212614 211574 238182
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 212398 133109 212458 283867
rect 212582 238645 212642 339627
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 218651 303788 218717 303789
rect 218651 303724 218652 303788
rect 218716 303724 218717 303788
rect 218651 303723 218717 303724
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 286182 218414 290898
rect 217547 284340 217613 284341
rect 217547 284276 217548 284340
rect 217612 284276 217613 284340
rect 217547 284275 217613 284276
rect 216443 284068 216509 284069
rect 216443 284004 216444 284068
rect 216508 284004 216509 284068
rect 216443 284003 216509 284004
rect 214419 283932 214485 283933
rect 214419 283868 214420 283932
rect 214484 283868 214485 283932
rect 214419 283867 214485 283868
rect 215523 283932 215589 283933
rect 215523 283868 215524 283932
rect 215588 283868 215589 283932
rect 215523 283867 215589 283868
rect 212579 238644 212645 238645
rect 212579 238580 212580 238644
rect 212644 238580 212645 238644
rect 212579 238579 212645 238580
rect 212579 237420 212645 237421
rect 212579 237356 212580 237420
rect 212644 237356 212645 237420
rect 212579 237355 212645 237356
rect 212582 204237 212642 237355
rect 214422 207093 214482 283867
rect 215526 233885 215586 283867
rect 215523 233884 215589 233885
rect 215523 233820 215524 233884
rect 215588 233820 215589 233884
rect 215523 233819 215589 233820
rect 214419 207092 214485 207093
rect 214419 207028 214420 207092
rect 214484 207028 214485 207092
rect 214419 207027 214485 207028
rect 212579 204236 212645 204237
rect 212579 204172 212580 204236
rect 212644 204172 212645 204236
rect 212579 204171 212645 204172
rect 213131 204236 213197 204237
rect 213131 204172 213132 204236
rect 213196 204172 213197 204236
rect 213131 204171 213197 204172
rect 213134 141405 213194 204171
rect 216446 181389 216506 284003
rect 217550 222325 217610 284275
rect 218654 238509 218714 303723
rect 221514 295174 222134 330618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 222331 315348 222397 315349
rect 222331 315284 222332 315348
rect 222396 315284 222397 315348
rect 222331 315283 222397 315284
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 286182 222134 294618
rect 219768 273454 220088 273486
rect 219768 273218 219810 273454
rect 220046 273218 220088 273454
rect 219768 273134 220088 273218
rect 219768 272898 219810 273134
rect 220046 272898 220088 273134
rect 219768 272866 220088 272898
rect 222334 238645 222394 315283
rect 225234 298894 225854 334338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 233739 361724 233805 361725
rect 233739 361660 233740 361724
rect 233804 361660 233805 361724
rect 233739 361659 233805 361660
rect 231899 351932 231965 351933
rect 231899 351868 231900 351932
rect 231964 351868 231965 351932
rect 231899 351867 231965 351868
rect 229691 350844 229757 350845
rect 229691 350780 229692 350844
rect 229756 350780 229757 350844
rect 229691 350779 229757 350780
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 227851 302836 227917 302837
rect 227851 302772 227852 302836
rect 227916 302772 227917 302836
rect 227851 302771 227917 302772
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 223619 291956 223685 291957
rect 223619 291892 223620 291956
rect 223684 291892 223685 291956
rect 223619 291891 223685 291892
rect 223622 285701 223682 291891
rect 225234 286182 225854 298338
rect 223803 285836 223869 285837
rect 223803 285772 223804 285836
rect 223868 285772 223869 285836
rect 223803 285771 223869 285772
rect 223619 285700 223685 285701
rect 223619 285636 223620 285700
rect 223684 285636 223685 285700
rect 223619 285635 223685 285636
rect 223806 277410 223866 285771
rect 224907 284340 224973 284341
rect 224907 284276 224908 284340
rect 224972 284276 224973 284340
rect 224907 284275 224973 284276
rect 223622 277350 223866 277410
rect 222331 238644 222397 238645
rect 222331 238580 222332 238644
rect 222396 238580 222397 238644
rect 222331 238579 222397 238580
rect 218651 238508 218717 238509
rect 218651 238444 218652 238508
rect 218716 238444 218717 238508
rect 218651 238443 218717 238444
rect 217547 222324 217613 222325
rect 217547 222260 217548 222324
rect 217612 222260 217613 222324
rect 217547 222259 217613 222260
rect 217794 219454 218414 238182
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 216443 181388 216509 181389
rect 216443 181324 216444 181388
rect 216508 181324 216509 181388
rect 216443 181323 216509 181324
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 213131 141404 213197 141405
rect 213131 141340 213132 141404
rect 213196 141340 213197 141404
rect 213131 141339 213197 141340
rect 212395 133108 212461 133109
rect 212395 133044 212396 133108
rect 212460 133044 212461 133108
rect 212395 133043 212461 133044
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 223174 222134 238182
rect 223622 238101 223682 277350
rect 224910 240141 224970 284275
rect 227483 283932 227549 283933
rect 227483 283868 227484 283932
rect 227548 283868 227549 283932
rect 227483 283867 227549 283868
rect 224907 240140 224973 240141
rect 224907 240076 224908 240140
rect 224972 240076 224973 240140
rect 224907 240075 224973 240076
rect 223619 238100 223685 238101
rect 223619 238036 223620 238100
rect 223684 238036 223685 238100
rect 223619 238035 223685 238036
rect 223622 237285 223682 238035
rect 223619 237284 223685 237285
rect 223619 237220 223620 237284
rect 223684 237220 223685 237284
rect 223619 237219 223685 237220
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 226894 225854 238182
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 227486 95165 227546 283867
rect 227854 240141 227914 302771
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 286182 229574 302058
rect 227851 240140 227917 240141
rect 227851 240076 227852 240140
rect 227916 240076 227917 240140
rect 227851 240075 227917 240076
rect 229694 238645 229754 350779
rect 230979 339556 231045 339557
rect 230979 339492 230980 339556
rect 231044 339492 231045 339556
rect 230979 339491 231045 339492
rect 229691 238644 229757 238645
rect 229691 238580 229692 238644
rect 229756 238580 229757 238644
rect 229691 238579 229757 238580
rect 230982 238237 231042 339491
rect 231902 240141 231962 351867
rect 231899 240140 231965 240141
rect 231899 240076 231900 240140
rect 231964 240076 231965 240140
rect 231899 240075 231965 240076
rect 233742 238645 233802 361659
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 286182 236414 308898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 240731 342276 240797 342277
rect 240731 342212 240732 342276
rect 240796 342212 240797 342276
rect 240731 342211 240797 342212
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 237419 297396 237485 297397
rect 237419 297332 237420 297396
rect 237484 297332 237485 297396
rect 237419 297331 237485 297332
rect 237235 283932 237301 283933
rect 237235 283868 237236 283932
rect 237300 283868 237301 283932
rect 237235 283867 237301 283868
rect 235128 255454 235448 255486
rect 235128 255218 235170 255454
rect 235406 255218 235448 255454
rect 235128 255134 235448 255218
rect 235128 254898 235170 255134
rect 235406 254898 235448 255134
rect 235128 254866 235448 254898
rect 233739 238644 233805 238645
rect 233739 238580 233740 238644
rect 233804 238580 233805 238644
rect 233739 238579 233805 238580
rect 230979 238236 231045 238237
rect 228954 230614 229574 238182
rect 230979 238172 230980 238236
rect 231044 238172 231045 238236
rect 230979 238171 231045 238172
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 227483 95164 227549 95165
rect 227483 95100 227484 95164
rect 227548 95100 227549 95164
rect 227483 95099 227549 95100
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 237454 236414 238182
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 237238 185741 237298 283867
rect 237422 240141 237482 297331
rect 239514 286182 240134 312618
rect 238523 284340 238589 284341
rect 238523 284276 238524 284340
rect 238588 284276 238589 284340
rect 238523 284275 238589 284276
rect 237419 240140 237485 240141
rect 237419 240076 237420 240140
rect 237484 240076 237485 240140
rect 237419 240075 237485 240076
rect 237235 185740 237301 185741
rect 237235 185676 237236 185740
rect 237300 185676 237301 185740
rect 237235 185675 237301 185676
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 238526 93125 238586 284275
rect 240734 248430 240794 342211
rect 243234 316894 243854 352338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 248459 360364 248525 360365
rect 248459 360300 248460 360364
rect 248524 360300 248525 360364
rect 248459 360299 248525 360300
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 244227 340916 244293 340917
rect 244227 340852 244228 340916
rect 244292 340852 244293 340916
rect 244227 340851 244293 340852
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 242939 293180 243005 293181
rect 242939 293116 242940 293180
rect 243004 293116 243005 293180
rect 242939 293115 243005 293116
rect 242942 285290 243002 293115
rect 243234 286182 243854 316338
rect 244230 306390 244290 340851
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 244230 306330 244474 306390
rect 242942 285230 244290 285290
rect 244230 284205 244290 285230
rect 244227 284204 244293 284205
rect 244227 284140 244228 284204
rect 244292 284140 244293 284204
rect 244227 284139 244293 284140
rect 244227 284068 244293 284069
rect 244227 284004 244228 284068
rect 244292 284004 244293 284068
rect 244227 284003 244293 284004
rect 244230 267069 244290 284003
rect 244414 281077 244474 306330
rect 246954 284614 247574 320058
rect 245699 284612 245765 284613
rect 245699 284548 245700 284612
rect 245764 284548 245765 284612
rect 245699 284547 245765 284548
rect 245702 282165 245762 284547
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 245699 282164 245765 282165
rect 245699 282100 245700 282164
rect 245764 282100 245765 282164
rect 245699 282099 245765 282100
rect 244411 281076 244477 281077
rect 244411 281012 244412 281076
rect 244476 281012 244477 281076
rect 244411 281011 244477 281012
rect 244227 267068 244293 267069
rect 244227 267004 244228 267068
rect 244292 267004 244293 267068
rect 244227 267003 244293 267004
rect 246954 248614 247574 284058
rect 248462 275365 248522 360299
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 248459 275364 248525 275365
rect 248459 275300 248460 275364
rect 248524 275300 248525 275364
rect 248459 275299 248525 275300
rect 240734 248370 241346 248430
rect 241286 238645 241346 248370
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 243491 246260 243557 246261
rect 243491 246196 243492 246260
rect 243556 246196 243557 246260
rect 243491 246195 243557 246196
rect 243494 238770 243554 246195
rect 245883 242996 245949 242997
rect 245883 242932 245884 242996
rect 245948 242932 245949 242996
rect 245883 242931 245949 242932
rect 245699 240276 245765 240277
rect 245699 240212 245700 240276
rect 245764 240212 245765 240276
rect 245699 240211 245765 240212
rect 242942 238710 243554 238770
rect 241283 238644 241349 238645
rect 241283 238580 241284 238644
rect 241348 238580 241349 238644
rect 241283 238579 241349 238580
rect 239514 205174 240134 238182
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 169174 240134 204618
rect 241286 194173 241346 238579
rect 242942 195941 243002 238710
rect 243234 208894 243854 238182
rect 245702 227493 245762 240211
rect 245886 230485 245946 242931
rect 245883 230484 245949 230485
rect 245883 230420 245884 230484
rect 245948 230420 245949 230484
rect 245883 230419 245949 230420
rect 245699 227492 245765 227493
rect 245699 227428 245700 227492
rect 245764 227428 245765 227492
rect 245699 227427 245765 227428
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 242939 195940 243005 195941
rect 242939 195876 242940 195940
rect 243004 195876 243005 195940
rect 242939 195875 243005 195876
rect 241283 194172 241349 194173
rect 241283 194108 241284 194172
rect 241348 194108 241349 194172
rect 241283 194107 241349 194108
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 238523 93124 238589 93125
rect 238523 93060 238524 93124
rect 238588 93060 238589 93124
rect 238523 93059 238589 93060
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 176614 247574 212058
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 178000 254414 182898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 258395 307868 258461 307869
rect 258395 307804 258396 307868
rect 258460 307804 258461 307868
rect 258395 307803 258461 307804
rect 258398 296730 258458 307803
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 178000 258134 186618
rect 258214 296670 258458 296730
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 258214 177581 258274 296670
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 178000 261854 190338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 270723 310724 270789 310725
rect 270723 310660 270724 310724
rect 270788 310660 270789 310724
rect 270723 310659 270789 310660
rect 269067 309364 269133 309365
rect 269067 309300 269068 309364
rect 269132 309300 269133 309364
rect 269067 309299 269133 309300
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 263915 178260 263981 178261
rect 263915 178196 263916 178260
rect 263980 178196 263981 178260
rect 263915 178195 263981 178196
rect 258211 177580 258277 177581
rect 258211 177516 258212 177580
rect 258276 177516 258277 177580
rect 258211 177515 258277 177516
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 263918 171150 263978 178195
rect 264954 178000 265574 194058
rect 265755 194036 265821 194037
rect 265755 193972 265756 194036
rect 265820 193972 265821 194036
rect 265755 193971 265821 193972
rect 265019 176764 265085 176765
rect 265019 176700 265020 176764
rect 265084 176700 265085 176764
rect 265019 176699 265085 176700
rect 263918 171090 264162 171150
rect 256207 165454 256527 165486
rect 256207 165218 256249 165454
rect 256485 165218 256527 165454
rect 256207 165134 256527 165218
rect 256207 164898 256249 165134
rect 256485 164898 256527 165134
rect 256207 164866 256527 164898
rect 259471 165454 259791 165486
rect 259471 165218 259513 165454
rect 259749 165218 259791 165454
rect 259471 165134 259791 165218
rect 259471 164898 259513 165134
rect 259749 164898 259791 165134
rect 259471 164866 259791 164898
rect 264102 151061 264162 171090
rect 265022 165613 265082 176699
rect 265019 165612 265085 165613
rect 265019 165548 265020 165612
rect 265084 165548 265085 165612
rect 265019 165547 265085 165548
rect 265571 164932 265637 164933
rect 265571 164868 265572 164932
rect 265636 164868 265637 164932
rect 265571 164867 265637 164868
rect 265019 154460 265085 154461
rect 265019 154396 265020 154460
rect 265084 154396 265085 154460
rect 265019 154395 265085 154396
rect 264099 151060 264165 151061
rect 264099 150996 264100 151060
rect 264164 150996 264165 151060
rect 264099 150995 264165 150996
rect 264099 150516 264165 150517
rect 264099 150452 264100 150516
rect 264164 150452 264165 150516
rect 264099 150451 264165 150452
rect 254575 147454 254895 147486
rect 254575 147218 254617 147454
rect 254853 147218 254895 147454
rect 254575 147134 254895 147218
rect 254575 146898 254617 147134
rect 254853 146898 254895 147134
rect 254575 146866 254895 146898
rect 257839 147454 258159 147486
rect 257839 147218 257881 147454
rect 258117 147218 258159 147454
rect 257839 147134 258159 147218
rect 257839 146898 257881 147134
rect 258117 146898 258159 147134
rect 257839 146866 258159 146898
rect 261103 147454 261423 147486
rect 261103 147218 261145 147454
rect 261381 147218 261423 147454
rect 261103 147134 261423 147218
rect 261103 146898 261145 147134
rect 261381 146898 261423 147134
rect 261103 146866 261423 146898
rect 264102 145349 264162 150451
rect 264099 145348 264165 145349
rect 264099 145284 264100 145348
rect 264164 145284 264165 145348
rect 264099 145283 264165 145284
rect 265022 142493 265082 154395
rect 265019 142492 265085 142493
rect 265019 142428 265020 142492
rect 265084 142428 265085 142492
rect 265019 142427 265085 142428
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 256207 129454 256527 129486
rect 256207 129218 256249 129454
rect 256485 129218 256527 129454
rect 256207 129134 256527 129218
rect 256207 128898 256249 129134
rect 256485 128898 256527 129134
rect 256207 128866 256527 128898
rect 259471 129454 259791 129486
rect 259471 129218 259513 129454
rect 259749 129218 259791 129454
rect 259471 129134 259791 129218
rect 259471 128898 259513 129134
rect 259749 128898 259791 129134
rect 259471 128866 259791 128898
rect 264099 113796 264165 113797
rect 264099 113732 264100 113796
rect 264164 113732 264165 113796
rect 264099 113731 264165 113732
rect 264102 113190 264162 113731
rect 264102 113130 264530 113190
rect 254575 111454 254895 111486
rect 254575 111218 254617 111454
rect 254853 111218 254895 111454
rect 254575 111134 254895 111218
rect 254575 110898 254617 111134
rect 254853 110898 254895 111134
rect 254575 110866 254895 110898
rect 257839 111454 258159 111486
rect 257839 111218 257881 111454
rect 258117 111218 258159 111454
rect 257839 111134 258159 111218
rect 257839 110898 257881 111134
rect 258117 110898 258159 111134
rect 257839 110866 258159 110898
rect 261103 111454 261423 111486
rect 261103 111218 261145 111454
rect 261381 111218 261423 111454
rect 261103 111134 261423 111218
rect 261103 110898 261145 111134
rect 261381 110898 261423 111134
rect 261103 110866 261423 110898
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 264099 99108 264165 99109
rect 264099 99044 264100 99108
rect 264164 99044 264165 99108
rect 264099 99043 264165 99044
rect 264102 98970 264162 99043
rect 263918 98910 264162 98970
rect 252507 97204 252573 97205
rect 252507 97140 252508 97204
rect 252572 97140 252573 97204
rect 252507 97139 252573 97140
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 252510 3501 252570 97139
rect 257846 96870 259562 96930
rect 257846 95981 257906 96870
rect 257843 95980 257909 95981
rect 257843 95916 257844 95980
rect 257908 95916 257909 95980
rect 257843 95915 257909 95916
rect 259315 95844 259381 95845
rect 259315 95780 259316 95844
rect 259380 95780 259381 95844
rect 259315 95779 259381 95780
rect 253794 75454 254414 94000
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 252507 3500 252573 3501
rect 252507 3436 252508 3500
rect 252572 3436 252573 3500
rect 252507 3435 252573 3436
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 79174 258134 94000
rect 259318 88229 259378 95779
rect 259315 88228 259381 88229
rect 259315 88164 259316 88228
rect 259380 88164 259381 88228
rect 259315 88163 259381 88164
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 259502 63613 259562 96870
rect 260971 95980 261037 95981
rect 260971 95916 260972 95980
rect 261036 95916 261037 95980
rect 260971 95915 261037 95916
rect 259499 63612 259565 63613
rect 259499 63548 259500 63612
rect 259564 63548 259565 63612
rect 259499 63547 259565 63548
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 260974 18597 261034 95915
rect 261234 82894 261854 94000
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 260971 18596 261037 18597
rect 260971 18532 260972 18596
rect 261036 18532 261037 18596
rect 260971 18531 261037 18532
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 46338
rect 263918 35189 263978 98910
rect 264470 98290 264530 113130
rect 265574 98973 265634 164867
rect 265758 154325 265818 193971
rect 266307 193220 266373 193221
rect 266307 193156 266308 193220
rect 266372 193156 266373 193220
rect 266307 193155 266373 193156
rect 266310 159085 266370 193155
rect 267779 185876 267845 185877
rect 267779 185812 267780 185876
rect 267844 185812 267845 185876
rect 267779 185811 267845 185812
rect 266859 172548 266925 172549
rect 266859 172484 266860 172548
rect 266924 172484 266925 172548
rect 266859 172483 266925 172484
rect 266307 159084 266373 159085
rect 266307 159020 266308 159084
rect 266372 159020 266373 159084
rect 266307 159019 266373 159020
rect 266862 156229 266922 172483
rect 267782 160173 267842 185811
rect 267963 180844 268029 180845
rect 267963 180780 267964 180844
rect 268028 180780 268029 180844
rect 267963 180779 268029 180780
rect 267966 172549 268026 180779
rect 267963 172548 268029 172549
rect 267963 172484 267964 172548
rect 268028 172484 268029 172548
rect 267963 172483 268029 172484
rect 268331 166292 268397 166293
rect 268331 166228 268332 166292
rect 268396 166228 268397 166292
rect 268331 166227 268397 166228
rect 267779 160172 267845 160173
rect 267779 160108 267780 160172
rect 267844 160108 267845 160172
rect 267779 160107 267845 160108
rect 267043 156636 267109 156637
rect 267043 156572 267044 156636
rect 267108 156572 267109 156636
rect 267043 156571 267109 156572
rect 266859 156228 266925 156229
rect 266859 156164 266860 156228
rect 266924 156164 266925 156228
rect 266859 156163 266925 156164
rect 265755 154324 265821 154325
rect 265755 154260 265756 154324
rect 265820 154260 265821 154324
rect 265755 154259 265821 154260
rect 266859 151196 266925 151197
rect 266859 151132 266860 151196
rect 266924 151132 266925 151196
rect 266859 151131 266925 151132
rect 265755 132836 265821 132837
rect 265755 132772 265756 132836
rect 265820 132772 265821 132836
rect 265755 132771 265821 132772
rect 265571 98972 265637 98973
rect 265571 98908 265572 98972
rect 265636 98908 265637 98972
rect 265571 98907 265637 98908
rect 264102 98230 264530 98290
rect 264102 50285 264162 98230
rect 264954 86614 265574 94000
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 265758 51781 265818 132771
rect 266862 123589 266922 151131
rect 267046 147797 267106 156571
rect 268334 151333 268394 166227
rect 269070 163845 269130 309299
rect 270539 290052 270605 290053
rect 270539 289988 270540 290052
rect 270604 289988 270605 290052
rect 270539 289987 270605 289988
rect 269251 213892 269317 213893
rect 269251 213828 269252 213892
rect 269316 213828 269317 213892
rect 269251 213827 269317 213828
rect 269254 169149 269314 213827
rect 269251 169148 269317 169149
rect 269251 169084 269252 169148
rect 269316 169084 269317 169148
rect 269251 169083 269317 169084
rect 270355 166564 270421 166565
rect 270355 166500 270356 166564
rect 270420 166500 270421 166564
rect 270355 166499 270421 166500
rect 269067 163844 269133 163845
rect 269067 163780 269068 163844
rect 269132 163780 269133 163844
rect 269067 163779 269133 163780
rect 269619 163436 269685 163437
rect 269619 163372 269620 163436
rect 269684 163372 269685 163436
rect 269619 163371 269685 163372
rect 268515 156908 268581 156909
rect 268515 156844 268516 156908
rect 268580 156844 268581 156908
rect 268515 156843 268581 156844
rect 268331 151332 268397 151333
rect 268331 151268 268332 151332
rect 268396 151268 268397 151332
rect 268331 151267 268397 151268
rect 267043 147796 267109 147797
rect 267043 147732 267044 147796
rect 267108 147732 267109 147796
rect 267043 147731 267109 147732
rect 268518 145893 268578 156843
rect 268699 149972 268765 149973
rect 268699 149908 268700 149972
rect 268764 149908 268765 149972
rect 268699 149907 268765 149908
rect 268515 145892 268581 145893
rect 268515 145828 268516 145892
rect 268580 145828 268581 145892
rect 268515 145827 268581 145828
rect 268331 145756 268397 145757
rect 268331 145692 268332 145756
rect 268396 145692 268397 145756
rect 268331 145691 268397 145692
rect 267227 142764 267293 142765
rect 267227 142700 267228 142764
rect 267292 142700 267293 142764
rect 267227 142699 267293 142700
rect 267230 124541 267290 142699
rect 267227 124540 267293 124541
rect 267227 124476 267228 124540
rect 267292 124476 267293 124540
rect 267227 124475 267293 124476
rect 266859 123588 266925 123589
rect 266859 123524 266860 123588
rect 266924 123524 266925 123588
rect 266859 123523 266925 123524
rect 266859 122092 266925 122093
rect 266859 122028 266860 122092
rect 266924 122028 266925 122092
rect 266859 122027 266925 122028
rect 266307 118012 266373 118013
rect 266307 117948 266308 118012
rect 266372 117948 266373 118012
rect 266307 117947 266373 117948
rect 266310 106181 266370 117947
rect 266307 106180 266373 106181
rect 266307 106116 266308 106180
rect 266372 106116 266373 106180
rect 266307 106115 266373 106116
rect 266862 57221 266922 122027
rect 267779 110532 267845 110533
rect 267779 110468 267780 110532
rect 267844 110468 267845 110532
rect 267779 110467 267845 110468
rect 267043 105500 267109 105501
rect 267043 105436 267044 105500
rect 267108 105436 267109 105500
rect 267043 105435 267109 105436
rect 267046 73949 267106 105435
rect 267782 87685 267842 110467
rect 268334 104685 268394 145691
rect 268702 112029 268762 149907
rect 269622 128213 269682 163371
rect 270358 157453 270418 166499
rect 270355 157452 270421 157453
rect 270355 157388 270356 157452
rect 270420 157388 270421 157452
rect 270355 157387 270421 157388
rect 269803 151060 269869 151061
rect 269803 150996 269804 151060
rect 269868 150996 269869 151060
rect 269803 150995 269869 150996
rect 269806 140725 269866 150995
rect 269803 140724 269869 140725
rect 269803 140660 269804 140724
rect 269868 140660 269869 140724
rect 269803 140659 269869 140660
rect 270355 140044 270421 140045
rect 270355 139980 270356 140044
rect 270420 139980 270421 140044
rect 270355 139979 270421 139980
rect 269803 138684 269869 138685
rect 269803 138620 269804 138684
rect 269868 138620 269869 138684
rect 269803 138619 269869 138620
rect 269619 128212 269685 128213
rect 269619 128148 269620 128212
rect 269684 128148 269685 128212
rect 269619 128147 269685 128148
rect 269806 121277 269866 138619
rect 270358 138277 270418 139979
rect 270355 138276 270421 138277
rect 270355 138212 270356 138276
rect 270420 138212 270421 138276
rect 270355 138211 270421 138212
rect 270542 137869 270602 289987
rect 270726 162757 270786 310659
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 277163 346492 277229 346493
rect 277163 346428 277164 346492
rect 277228 346428 277229 346492
rect 277163 346427 277229 346428
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 273299 296852 273365 296853
rect 273299 296788 273300 296852
rect 273364 296788 273365 296852
rect 273299 296787 273365 296788
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 272563 188460 272629 188461
rect 272563 188396 272564 188460
rect 272628 188396 272629 188460
rect 272563 188395 272629 188396
rect 272566 165613 272626 188395
rect 272563 165612 272629 165613
rect 272563 165548 272564 165612
rect 272628 165548 272629 165612
rect 272563 165547 272629 165548
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 270723 162756 270789 162757
rect 270723 162692 270724 162756
rect 270788 162692 270789 162756
rect 270723 162691 270789 162692
rect 271091 145892 271157 145893
rect 271091 145828 271092 145892
rect 271156 145828 271157 145892
rect 271091 145827 271157 145828
rect 270539 137868 270605 137869
rect 270539 137804 270540 137868
rect 270604 137804 270605 137868
rect 270539 137803 270605 137804
rect 270355 127124 270421 127125
rect 270355 127060 270356 127124
rect 270420 127060 270421 127124
rect 270355 127059 270421 127060
rect 269803 121276 269869 121277
rect 269803 121212 269804 121276
rect 269868 121212 269869 121276
rect 269803 121211 269869 121212
rect 269067 114748 269133 114749
rect 269067 114684 269068 114748
rect 269132 114684 269133 114748
rect 269067 114683 269133 114684
rect 268699 112028 268765 112029
rect 268699 111964 268700 112028
rect 268764 111964 268765 112028
rect 268699 111963 268765 111964
rect 268331 104684 268397 104685
rect 268331 104620 268332 104684
rect 268396 104620 268397 104684
rect 268331 104619 268397 104620
rect 269070 102509 269130 114683
rect 269619 109716 269685 109717
rect 269619 109652 269620 109716
rect 269684 109652 269685 109716
rect 269619 109651 269685 109652
rect 269067 102508 269133 102509
rect 269067 102444 269068 102508
rect 269132 102444 269133 102508
rect 269067 102443 269133 102444
rect 269067 102372 269133 102373
rect 269067 102308 269068 102372
rect 269132 102308 269133 102372
rect 269067 102307 269133 102308
rect 267963 102236 268029 102237
rect 267963 102172 267964 102236
rect 268028 102172 268029 102236
rect 267963 102171 268029 102172
rect 267779 87684 267845 87685
rect 267779 87620 267780 87684
rect 267844 87620 267845 87684
rect 267779 87619 267845 87620
rect 267966 86189 268026 102171
rect 267963 86188 268029 86189
rect 267963 86124 267964 86188
rect 268028 86124 268029 86188
rect 267963 86123 268029 86124
rect 267043 73948 267109 73949
rect 267043 73884 267044 73948
rect 267108 73884 267109 73948
rect 267043 73883 267109 73884
rect 266859 57220 266925 57221
rect 266859 57156 266860 57220
rect 266924 57156 266925 57220
rect 266859 57155 266925 57156
rect 269070 53141 269130 102307
rect 269622 74085 269682 109651
rect 270358 109173 270418 127059
rect 270355 109172 270421 109173
rect 270355 109108 270356 109172
rect 270420 109108 270421 109172
rect 270355 109107 270421 109108
rect 271094 104277 271154 145827
rect 271643 134468 271709 134469
rect 271643 134404 271644 134468
rect 271708 134404 271709 134468
rect 271643 134403 271709 134404
rect 271646 115837 271706 134403
rect 271794 129454 272414 164898
rect 273302 154869 273362 296787
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 273483 220284 273549 220285
rect 273483 220220 273484 220284
rect 273548 220220 273549 220284
rect 273483 220219 273549 220220
rect 273486 164253 273546 220219
rect 275514 205174 276134 240618
rect 276243 223548 276309 223549
rect 276243 223484 276244 223548
rect 276308 223484 276309 223548
rect 276243 223483 276309 223484
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275139 189684 275205 189685
rect 275139 189620 275140 189684
rect 275204 189620 275205 189684
rect 275139 189619 275205 189620
rect 273483 164252 273549 164253
rect 273483 164188 273484 164252
rect 273548 164188 273549 164252
rect 273483 164187 273549 164188
rect 274035 161532 274101 161533
rect 274035 161468 274036 161532
rect 274100 161468 274101 161532
rect 274035 161467 274101 161468
rect 273483 155956 273549 155957
rect 273483 155892 273484 155956
rect 273548 155892 273549 155956
rect 273483 155891 273549 155892
rect 273299 154868 273365 154869
rect 273299 154804 273300 154868
rect 273364 154804 273365 154868
rect 273299 154803 273365 154804
rect 272563 149836 272629 149837
rect 272563 149772 272564 149836
rect 272628 149772 272629 149836
rect 272563 149771 272629 149772
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271643 115836 271709 115837
rect 271643 115772 271644 115836
rect 271708 115772 271709 115836
rect 271643 115771 271709 115772
rect 271275 114884 271341 114885
rect 271275 114820 271276 114884
rect 271340 114820 271341 114884
rect 271275 114819 271341 114820
rect 271091 104276 271157 104277
rect 271091 104212 271092 104276
rect 271156 104212 271157 104276
rect 271091 104211 271157 104212
rect 270539 100876 270605 100877
rect 270539 100812 270540 100876
rect 270604 100812 270605 100876
rect 270539 100811 270605 100812
rect 270542 95981 270602 100811
rect 270723 96524 270789 96525
rect 270723 96460 270724 96524
rect 270788 96460 270789 96524
rect 270723 96459 270789 96460
rect 270539 95980 270605 95981
rect 270539 95916 270540 95980
rect 270604 95916 270605 95980
rect 270539 95915 270605 95916
rect 270726 82381 270786 96459
rect 270723 82380 270789 82381
rect 270723 82316 270724 82380
rect 270788 82316 270789 82380
rect 270723 82315 270789 82316
rect 271278 79525 271338 114819
rect 271794 93454 272414 128898
rect 272566 108901 272626 149771
rect 273486 140861 273546 155891
rect 273851 141404 273917 141405
rect 273851 141340 273852 141404
rect 273916 141340 273917 141404
rect 273851 141339 273917 141340
rect 273483 140860 273549 140861
rect 273483 140796 273484 140860
rect 273548 140796 273549 140860
rect 273483 140795 273549 140796
rect 273299 121684 273365 121685
rect 273299 121620 273300 121684
rect 273364 121620 273365 121684
rect 273299 121619 273365 121620
rect 273302 117877 273362 121619
rect 273299 117876 273365 117877
rect 273299 117812 273300 117876
rect 273364 117812 273365 117876
rect 273299 117811 273365 117812
rect 272563 108900 272629 108901
rect 272563 108836 272564 108900
rect 272628 108836 272629 108900
rect 272563 108835 272629 108836
rect 272563 104820 272629 104821
rect 272563 104756 272564 104820
rect 272628 104756 272629 104820
rect 272563 104755 272629 104756
rect 272566 101013 272626 104755
rect 272563 101012 272629 101013
rect 272563 100948 272564 101012
rect 272628 100948 272629 101012
rect 272563 100947 272629 100948
rect 273854 100061 273914 141339
rect 274038 123453 274098 161467
rect 274035 123452 274101 123453
rect 274035 123388 274036 123452
rect 274100 123388 274101 123452
rect 274035 123387 274101 123388
rect 274035 117876 274101 117877
rect 274035 117812 274036 117876
rect 274100 117812 274101 117876
rect 274035 117811 274101 117812
rect 273851 100060 273917 100061
rect 273851 99996 273852 100060
rect 273916 99996 273917 100060
rect 273851 99995 273917 99996
rect 273851 98836 273917 98837
rect 273851 98772 273852 98836
rect 273916 98772 273917 98836
rect 273851 98771 273917 98772
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271275 79524 271341 79525
rect 271275 79460 271276 79524
rect 271340 79460 271341 79524
rect 271275 79459 271341 79460
rect 269619 74084 269685 74085
rect 269619 74020 269620 74084
rect 269684 74020 269685 74084
rect 269619 74019 269685 74020
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 269067 53140 269133 53141
rect 269067 53076 269068 53140
rect 269132 53076 269133 53140
rect 269067 53075 269133 53076
rect 265755 51780 265821 51781
rect 265755 51716 265756 51780
rect 265820 51716 265821 51780
rect 265755 51715 265821 51716
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264099 50284 264165 50285
rect 264099 50220 264100 50284
rect 264164 50220 264165 50284
rect 264099 50219 264165 50220
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 263915 35188 263981 35189
rect 263915 35124 263916 35188
rect 263980 35124 263981 35188
rect 263915 35123 263981 35124
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 273854 21317 273914 98771
rect 274038 89181 274098 117811
rect 274035 89180 274101 89181
rect 274035 89116 274036 89180
rect 274100 89116 274101 89180
rect 274035 89115 274101 89116
rect 273851 21316 273917 21317
rect 273851 21252 273852 21316
rect 273916 21252 273917 21316
rect 273851 21251 273917 21252
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 275142 3365 275202 189619
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 276246 162485 276306 223483
rect 276611 215932 276677 215933
rect 276611 215868 276612 215932
rect 276676 215868 276677 215932
rect 276611 215867 276677 215868
rect 276614 176765 276674 215867
rect 276611 176764 276677 176765
rect 276611 176700 276612 176764
rect 276676 176700 276677 176764
rect 276611 176699 276677 176700
rect 276243 162484 276309 162485
rect 276243 162420 276244 162484
rect 276308 162420 276309 162484
rect 276243 162419 276309 162420
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 276243 118012 276309 118013
rect 276243 117948 276244 118012
rect 276308 117948 276309 118012
rect 276243 117947 276309 117948
rect 276246 97205 276306 117947
rect 276614 97341 276674 176699
rect 276795 152148 276861 152149
rect 276795 152084 276796 152148
rect 276860 152084 276861 152148
rect 276795 152083 276861 152084
rect 276798 118149 276858 152083
rect 276795 118148 276861 118149
rect 276795 118084 276796 118148
rect 276860 118084 276861 118148
rect 276795 118083 276861 118084
rect 276611 97340 276677 97341
rect 276611 97276 276612 97340
rect 276676 97276 276677 97340
rect 276611 97275 276677 97276
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 276243 97204 276309 97205
rect 276243 97140 276244 97204
rect 276308 97140 276309 97204
rect 276243 97139 276309 97140
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 276795 96660 276861 96661
rect 276795 96596 276796 96660
rect 276860 96596 276861 96660
rect 276795 96595 276861 96596
rect 276798 76533 276858 96595
rect 276795 76532 276861 76533
rect 276795 76468 276796 76532
rect 276860 76468 276861 76532
rect 276795 76467 276861 76468
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275139 3364 275205 3365
rect 275139 3300 275140 3364
rect 275204 3300 275205 3364
rect 275139 3299 275205 3300
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 -3226 276134 24618
rect 277166 4045 277226 346427
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 278819 229940 278885 229941
rect 278819 229876 278820 229940
rect 278884 229876 278885 229940
rect 278819 229875 278885 229876
rect 277531 210628 277597 210629
rect 277531 210564 277532 210628
rect 277596 210564 277597 210628
rect 277531 210563 277597 210564
rect 277534 140997 277594 210563
rect 278822 157453 278882 229875
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 287099 298484 287165 298485
rect 287099 298420 287100 298484
rect 287164 298420 287165 298484
rect 287099 298419 287165 298420
rect 284339 292772 284405 292773
rect 284339 292708 284340 292772
rect 284404 292708 284405 292772
rect 284339 292707 284405 292708
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 281763 199476 281829 199477
rect 281763 199412 281764 199476
rect 281828 199412 281829 199476
rect 281763 199411 281829 199412
rect 281579 192540 281645 192541
rect 281579 192476 281580 192540
rect 281644 192476 281645 192540
rect 281579 192475 281645 192476
rect 280291 190636 280357 190637
rect 280291 190572 280292 190636
rect 280356 190572 280357 190636
rect 280291 190571 280357 190572
rect 280294 180810 280354 190571
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 278819 157452 278885 157453
rect 278819 157388 278820 157452
rect 278884 157388 278885 157452
rect 278819 157387 278885 157388
rect 278819 144804 278885 144805
rect 278819 144740 278820 144804
rect 278884 144740 278885 144804
rect 278819 144739 278885 144740
rect 277531 140996 277597 140997
rect 277531 140932 277532 140996
rect 277596 140932 277597 140996
rect 277531 140931 277597 140932
rect 278635 135692 278701 135693
rect 278635 135628 278636 135692
rect 278700 135628 278701 135692
rect 278635 135627 278701 135628
rect 278638 134605 278698 135627
rect 278822 135285 278882 144739
rect 279234 136894 279854 172338
rect 280110 180750 280354 180810
rect 280110 153781 280170 180750
rect 280291 180028 280357 180029
rect 280291 179964 280292 180028
rect 280356 179964 280357 180028
rect 280291 179963 280357 179964
rect 280107 153780 280173 153781
rect 280107 153716 280108 153780
rect 280172 153716 280173 153780
rect 280107 153715 280173 153716
rect 280294 144805 280354 179963
rect 280659 153372 280725 153373
rect 280659 153308 280660 153372
rect 280724 153308 280725 153372
rect 280659 153307 280725 153308
rect 280291 144804 280357 144805
rect 280291 144740 280292 144804
rect 280356 144740 280357 144804
rect 280291 144739 280357 144740
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 278819 135284 278885 135285
rect 278819 135220 278820 135284
rect 278884 135220 278885 135284
rect 278819 135219 278885 135220
rect 278635 134604 278701 134605
rect 278635 134540 278636 134604
rect 278700 134540 278701 134604
rect 278635 134539 278701 134540
rect 277899 134196 277965 134197
rect 277899 134132 277900 134196
rect 277964 134132 277965 134196
rect 277899 134131 277965 134132
rect 277902 61437 277962 134131
rect 279003 120324 279069 120325
rect 279003 120260 279004 120324
rect 279068 120260 279069 120324
rect 279003 120259 279069 120260
rect 279006 95845 279066 120259
rect 279234 100894 279854 136338
rect 280662 111757 280722 153307
rect 280843 143172 280909 143173
rect 280843 143108 280844 143172
rect 280908 143108 280909 143172
rect 280843 143107 280909 143108
rect 280659 111756 280725 111757
rect 280659 111692 280660 111756
rect 280724 111692 280725 111756
rect 280659 111691 280725 111692
rect 280291 106180 280357 106181
rect 280291 106116 280292 106180
rect 280356 106116 280357 106180
rect 280291 106115 280357 106116
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279003 95844 279069 95845
rect 279003 95780 279004 95844
rect 279068 95780 279069 95844
rect 279003 95779 279069 95780
rect 279234 64894 279854 100338
rect 280294 69597 280354 106115
rect 280846 102101 280906 143107
rect 281582 136917 281642 192475
rect 281766 146437 281826 199411
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 281763 146436 281829 146437
rect 281763 146372 281764 146436
rect 281828 146372 281829 146436
rect 281763 146371 281829 146372
rect 282954 140614 283574 176058
rect 283787 162756 283853 162757
rect 283787 162692 283788 162756
rect 283852 162692 283853 162756
rect 283787 162691 283853 162692
rect 283790 149701 283850 162691
rect 283787 149700 283853 149701
rect 283787 149636 283788 149700
rect 283852 149636 283853 149700
rect 283787 149635 283853 149636
rect 284342 145621 284402 292707
rect 284523 210492 284589 210493
rect 284523 210428 284524 210492
rect 284588 210428 284589 210492
rect 284523 210427 284589 210428
rect 284526 150517 284586 210427
rect 285811 196756 285877 196757
rect 285811 196692 285812 196756
rect 285876 196692 285877 196756
rect 285811 196691 285877 196692
rect 285627 195396 285693 195397
rect 285627 195332 285628 195396
rect 285692 195332 285693 195396
rect 285627 195331 285693 195332
rect 284523 150516 284589 150517
rect 284523 150452 284524 150516
rect 284588 150452 284589 150516
rect 284523 150451 284589 150452
rect 285075 149292 285141 149293
rect 285075 149228 285076 149292
rect 285140 149228 285141 149292
rect 285075 149227 285141 149228
rect 284339 145620 284405 145621
rect 284339 145556 284340 145620
rect 284404 145556 284405 145620
rect 284339 145555 284405 145556
rect 283787 140996 283853 140997
rect 283787 140932 283788 140996
rect 283852 140932 283853 140996
rect 283787 140931 283853 140932
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282499 139772 282565 139773
rect 282499 139708 282500 139772
rect 282564 139708 282565 139772
rect 282499 139707 282565 139708
rect 281579 136916 281645 136917
rect 281579 136852 281580 136916
rect 281644 136852 281645 136916
rect 281579 136851 281645 136852
rect 282315 136916 282381 136917
rect 282315 136852 282316 136916
rect 282380 136852 282381 136916
rect 282315 136851 282381 136852
rect 282318 135010 282378 136851
rect 282134 134950 282378 135010
rect 280843 102100 280909 102101
rect 280843 102036 280844 102100
rect 280908 102036 280909 102100
rect 280843 102035 280909 102036
rect 280291 69596 280357 69597
rect 280291 69532 280292 69596
rect 280356 69532 280357 69596
rect 280291 69531 280357 69532
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 277899 61436 277965 61437
rect 277899 61372 277900 61436
rect 277964 61372 277965 61436
rect 277899 61371 277965 61372
rect 279234 28894 279854 64338
rect 282134 58717 282194 134950
rect 282502 131749 282562 139707
rect 282499 131748 282565 131749
rect 282499 131684 282500 131748
rect 282564 131684 282565 131748
rect 282499 131683 282565 131684
rect 282315 128348 282381 128349
rect 282315 128284 282316 128348
rect 282380 128284 282381 128348
rect 282315 128283 282381 128284
rect 282318 122229 282378 128283
rect 282315 122228 282381 122229
rect 282315 122164 282316 122228
rect 282380 122164 282381 122228
rect 282315 122163 282381 122164
rect 282315 119508 282381 119509
rect 282315 119444 282316 119508
rect 282380 119444 282381 119508
rect 282315 119443 282381 119444
rect 282318 76669 282378 119443
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282315 76668 282381 76669
rect 282315 76604 282316 76668
rect 282380 76604 282381 76668
rect 282315 76603 282381 76604
rect 282954 68614 283574 104058
rect 283790 98701 283850 140931
rect 284891 135420 284957 135421
rect 284891 135356 284892 135420
rect 284956 135356 284957 135420
rect 284891 135355 284957 135356
rect 284339 101012 284405 101013
rect 284339 100948 284340 101012
rect 284404 100948 284405 101012
rect 284339 100947 284405 100948
rect 283787 98700 283853 98701
rect 283787 98636 283788 98700
rect 283852 98636 283853 98700
rect 283787 98635 283853 98636
rect 283971 98020 284037 98021
rect 283971 97956 283972 98020
rect 284036 97956 284037 98020
rect 283971 97955 284037 97956
rect 283974 83469 284034 97955
rect 283971 83468 284037 83469
rect 283971 83404 283972 83468
rect 284036 83404 284037 83468
rect 283971 83403 284037 83404
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282131 58716 282197 58717
rect 282131 58652 282132 58716
rect 282196 58652 282197 58716
rect 282131 58651 282197 58652
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 277163 4044 277229 4045
rect 277163 3980 277164 4044
rect 277228 3980 277229 4044
rect 277163 3979 277229 3980
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 68058
rect 284342 44845 284402 100947
rect 284339 44844 284405 44845
rect 284339 44780 284340 44844
rect 284404 44780 284405 44844
rect 284339 44779 284405 44780
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 284894 17237 284954 135355
rect 285078 107541 285138 149227
rect 285630 139501 285690 195331
rect 285814 151061 285874 196691
rect 285811 151060 285877 151061
rect 285811 150996 285812 151060
rect 285876 150996 285877 151060
rect 285811 150995 285877 150996
rect 286179 142220 286245 142221
rect 286179 142156 286180 142220
rect 286244 142156 286245 142220
rect 286179 142155 286245 142156
rect 285627 139500 285693 139501
rect 285627 139436 285628 139500
rect 285692 139436 285693 139500
rect 285627 139435 285693 139436
rect 285627 112028 285693 112029
rect 285627 111964 285628 112028
rect 285692 111964 285693 112028
rect 285627 111963 285693 111964
rect 285075 107540 285141 107541
rect 285075 107476 285076 107540
rect 285140 107476 285141 107540
rect 285075 107475 285141 107476
rect 284891 17236 284957 17237
rect 284891 17172 284892 17236
rect 284956 17172 284957 17236
rect 284891 17171 284957 17172
rect 285630 15877 285690 111963
rect 286182 101421 286242 142155
rect 287102 137053 287162 298419
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 288939 185604 289005 185605
rect 288939 185540 288940 185604
rect 289004 185540 289005 185604
rect 288939 185539 289005 185540
rect 288387 157452 288453 157453
rect 288387 157388 288388 157452
rect 288452 157388 288453 157452
rect 288387 157387 288453 157388
rect 288203 140452 288269 140453
rect 288203 140388 288204 140452
rect 288268 140388 288269 140452
rect 288203 140387 288269 140388
rect 287099 137052 287165 137053
rect 287099 136988 287100 137052
rect 287164 136988 287165 137052
rect 287099 136987 287165 136988
rect 287835 134876 287901 134877
rect 287835 134812 287836 134876
rect 287900 134812 287901 134876
rect 287835 134811 287901 134812
rect 286547 130388 286613 130389
rect 286547 130324 286548 130388
rect 286612 130324 286613 130388
rect 286547 130323 286613 130324
rect 286550 115837 286610 130323
rect 287651 128484 287717 128485
rect 287651 128420 287652 128484
rect 287716 128420 287717 128484
rect 287651 128419 287717 128420
rect 286547 115836 286613 115837
rect 286547 115772 286548 115836
rect 286612 115772 286613 115836
rect 286547 115771 286613 115772
rect 287099 112028 287165 112029
rect 287099 111964 287100 112028
rect 287164 111964 287165 112028
rect 287099 111963 287165 111964
rect 286179 101420 286245 101421
rect 286179 101356 286180 101420
rect 286244 101356 286245 101420
rect 286179 101355 286245 101356
rect 286179 99788 286245 99789
rect 286179 99724 286180 99788
rect 286244 99724 286245 99788
rect 286179 99723 286245 99724
rect 286182 48925 286242 99723
rect 287102 54501 287162 111963
rect 287099 54500 287165 54501
rect 287099 54436 287100 54500
rect 287164 54436 287165 54500
rect 287099 54435 287165 54436
rect 286179 48924 286245 48925
rect 286179 48860 286180 48924
rect 286244 48860 286245 48924
rect 286179 48859 286245 48860
rect 287654 37909 287714 128419
rect 287838 113253 287898 134811
rect 288206 134469 288266 140387
rect 288390 138413 288450 157387
rect 288387 138412 288453 138413
rect 288387 138348 288388 138412
rect 288452 138348 288453 138412
rect 288387 138347 288453 138348
rect 288203 134468 288269 134469
rect 288203 134404 288204 134468
rect 288268 134404 288269 134468
rect 288203 134403 288269 134404
rect 287835 113252 287901 113253
rect 287835 113188 287836 113252
rect 287900 113188 287901 113252
rect 287835 113187 287901 113188
rect 287651 37908 287717 37909
rect 287651 37844 287652 37908
rect 287716 37844 287717 37908
rect 287651 37843 287717 37844
rect 285627 15876 285693 15877
rect 285627 15812 285628 15876
rect 285692 15812 285693 15876
rect 285627 15811 285693 15812
rect 288942 3501 289002 185539
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 178000 290414 182898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 290595 178124 290661 178125
rect 290595 178060 290596 178124
rect 290660 178060 290661 178124
rect 290595 178059 290661 178060
rect 290598 138005 290658 178059
rect 293514 178000 294134 186618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 306419 287740 306485 287741
rect 306419 287676 306420 287740
rect 306484 287676 306485 287740
rect 306419 287675 306485 287676
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 298139 244900 298205 244901
rect 298139 244836 298140 244900
rect 298204 244836 298205 244900
rect 298139 244835 298205 244836
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 178000 297854 190338
rect 298142 175949 298202 244835
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 302187 216748 302253 216749
rect 302187 216684 302188 216748
rect 302252 216684 302253 216748
rect 302187 216683 302253 216684
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 178000 301574 194058
rect 301819 180028 301885 180029
rect 301819 179964 301820 180028
rect 301884 179964 301885 180028
rect 301819 179963 301885 179964
rect 301267 177444 301333 177445
rect 301267 177380 301268 177444
rect 301332 177380 301333 177444
rect 301267 177379 301333 177380
rect 298139 175948 298205 175949
rect 298139 175884 298140 175948
rect 298204 175884 298205 175948
rect 298139 175883 298205 175884
rect 301270 173773 301330 177379
rect 301267 173772 301333 173773
rect 301267 173708 301268 173772
rect 301332 173708 301333 173772
rect 301267 173707 301333 173708
rect 294207 165454 294527 165486
rect 294207 165218 294249 165454
rect 294485 165218 294527 165454
rect 294207 165134 294527 165218
rect 294207 164898 294249 165134
rect 294485 164898 294527 165134
rect 294207 164866 294527 164898
rect 297471 165454 297791 165486
rect 297471 165218 297513 165454
rect 297749 165218 297791 165454
rect 297471 165134 297791 165218
rect 297471 164898 297513 165134
rect 297749 164898 297791 165134
rect 297471 164866 297791 164898
rect 292575 147454 292895 147486
rect 292575 147218 292617 147454
rect 292853 147218 292895 147454
rect 292575 147134 292895 147218
rect 292575 146898 292617 147134
rect 292853 146898 292895 147134
rect 292575 146866 292895 146898
rect 295839 147454 296159 147486
rect 295839 147218 295881 147454
rect 296117 147218 296159 147454
rect 295839 147134 296159 147218
rect 295839 146898 295881 147134
rect 296117 146898 296159 147134
rect 295839 146866 296159 146898
rect 299103 147454 299423 147486
rect 299103 147218 299145 147454
rect 299381 147218 299423 147454
rect 299103 147134 299423 147218
rect 299103 146898 299145 147134
rect 299381 146898 299423 147134
rect 301822 147117 301882 179963
rect 301819 147116 301885 147117
rect 301819 147052 301820 147116
rect 301884 147052 301885 147116
rect 301819 147051 301885 147052
rect 299103 146866 299423 146898
rect 290595 138004 290661 138005
rect 290595 137940 290596 138004
rect 290660 137940 290661 138004
rect 290595 137939 290661 137940
rect 302190 136645 302250 216683
rect 304947 190500 305013 190501
rect 304947 190436 304948 190500
rect 305012 190436 305013 190500
rect 304947 190435 305013 190436
rect 302371 181388 302437 181389
rect 302371 181324 302372 181388
rect 302436 181324 302437 181388
rect 302371 181323 302437 181324
rect 302374 140453 302434 181323
rect 302371 140452 302437 140453
rect 302371 140388 302372 140452
rect 302436 140388 302437 140452
rect 302371 140387 302437 140388
rect 302187 136644 302253 136645
rect 302187 136580 302188 136644
rect 302252 136580 302253 136644
rect 302187 136579 302253 136580
rect 290227 133788 290293 133789
rect 290227 133724 290228 133788
rect 290292 133724 290293 133788
rect 290227 133723 290293 133724
rect 289123 131476 289189 131477
rect 289123 131412 289124 131476
rect 289188 131412 289189 131476
rect 289123 131411 289189 131412
rect 289126 64157 289186 131411
rect 289859 128892 289925 128893
rect 289859 128828 289860 128892
rect 289924 128828 289925 128892
rect 289859 128827 289925 128828
rect 289862 94893 289922 128827
rect 290230 122850 290290 133723
rect 294207 129454 294527 129486
rect 294207 129218 294249 129454
rect 294485 129218 294527 129454
rect 294207 129134 294527 129218
rect 294207 128898 294249 129134
rect 294485 128898 294527 129134
rect 294207 128866 294527 128898
rect 297471 129454 297791 129486
rect 297471 129218 297513 129454
rect 297749 129218 297791 129454
rect 297471 129134 297791 129218
rect 297471 128898 297513 129134
rect 297749 128898 297791 129134
rect 297471 128866 297791 128898
rect 290046 122790 290290 122850
rect 290046 113117 290106 122790
rect 304950 120733 305010 190435
rect 305131 180164 305197 180165
rect 305131 180100 305132 180164
rect 305196 180100 305197 180164
rect 305131 180099 305197 180100
rect 305134 167925 305194 180099
rect 305131 167924 305197 167925
rect 305131 167860 305132 167924
rect 305196 167860 305197 167924
rect 305131 167859 305197 167860
rect 306422 142765 306482 287675
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 310467 210356 310533 210357
rect 310467 210292 310468 210356
rect 310532 210292 310533 210356
rect 310467 210291 310533 210292
rect 309179 202332 309245 202333
rect 309179 202268 309180 202332
rect 309244 202268 309245 202332
rect 309179 202267 309245 202268
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 306603 176628 306669 176629
rect 306603 176564 306604 176628
rect 306668 176564 306669 176628
rect 306603 176563 306669 176564
rect 306606 164389 306666 176563
rect 307794 165454 308414 200898
rect 308627 178668 308693 178669
rect 308627 178604 308628 178668
rect 308692 178604 308693 178668
rect 308627 178603 308693 178604
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 306603 164388 306669 164389
rect 306603 164324 306604 164388
rect 306668 164324 306669 164388
rect 306603 164323 306669 164324
rect 306419 142764 306485 142765
rect 306419 142700 306420 142764
rect 306484 142700 306485 142764
rect 306419 142699 306485 142700
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 304947 120732 305013 120733
rect 304947 120668 304948 120732
rect 305012 120668 305013 120732
rect 304947 120667 305013 120668
rect 290043 113116 290109 113117
rect 290043 113052 290044 113116
rect 290108 113052 290109 113116
rect 290043 113051 290109 113052
rect 292575 111454 292895 111486
rect 292575 111218 292617 111454
rect 292853 111218 292895 111454
rect 292575 111134 292895 111218
rect 292575 110898 292617 111134
rect 292853 110898 292895 111134
rect 292575 110866 292895 110898
rect 295839 111454 296159 111486
rect 295839 111218 295881 111454
rect 296117 111218 296159 111454
rect 295839 111134 296159 111218
rect 295839 110898 295881 111134
rect 296117 110898 296159 111134
rect 295839 110866 296159 110898
rect 299103 111454 299423 111486
rect 299103 111218 299145 111454
rect 299381 111218 299423 111454
rect 299103 111134 299423 111218
rect 299103 110898 299145 111134
rect 299381 110898 299423 111134
rect 299103 110866 299423 110898
rect 303659 106180 303725 106181
rect 303659 106116 303660 106180
rect 303724 106116 303725 106180
rect 303659 106115 303725 106116
rect 290595 102780 290661 102781
rect 290595 102716 290596 102780
rect 290660 102716 290661 102780
rect 290595 102715 290661 102716
rect 289859 94892 289925 94893
rect 289859 94828 289860 94892
rect 289924 94828 289925 94892
rect 289859 94827 289925 94828
rect 289794 75454 290414 94000
rect 290598 80885 290658 102715
rect 290595 80884 290661 80885
rect 290595 80820 290596 80884
rect 290660 80820 290661 80884
rect 290595 80819 290661 80820
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289123 64156 289189 64157
rect 289123 64092 289124 64156
rect 289188 64092 289189 64156
rect 289123 64091 289189 64092
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 288939 3500 289005 3501
rect 288939 3436 288940 3500
rect 289004 3436 289005 3500
rect 288939 3435 289005 3436
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 79174 294134 94000
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 82894 297854 94000
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 86614 301574 94000
rect 303662 88229 303722 106115
rect 307794 93454 308414 128898
rect 308630 126853 308690 178603
rect 308627 126852 308693 126853
rect 308627 126788 308628 126852
rect 308692 126788 308693 126852
rect 308627 126787 308693 126788
rect 309182 109445 309242 202267
rect 309731 193900 309797 193901
rect 309731 193836 309732 193900
rect 309796 193836 309797 193900
rect 309731 193835 309797 193836
rect 309179 109444 309245 109445
rect 309179 109380 309180 109444
rect 309244 109380 309245 109444
rect 309179 109379 309245 109380
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 303659 88228 303725 88229
rect 303659 88164 303660 88228
rect 303724 88164 303725 88228
rect 303659 88163 303725 88164
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 309734 4045 309794 193835
rect 310470 116245 310530 210291
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 317459 358868 317525 358869
rect 317459 358804 317460 358868
rect 317524 358804 317525 358868
rect 317459 358803 317525 358804
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315987 306644 316053 306645
rect 315987 306580 315988 306644
rect 316052 306580 316053 306644
rect 315987 306579 316053 306580
rect 315990 306373 316050 306579
rect 315987 306372 316053 306373
rect 315987 306308 315988 306372
rect 316052 306308 316053 306372
rect 315987 306307 316053 306308
rect 316171 296852 316237 296853
rect 316171 296850 316172 296852
rect 315990 296790 316172 296850
rect 315990 296581 316050 296790
rect 316171 296788 316172 296790
rect 316236 296788 316237 296852
rect 316171 296787 316237 296788
rect 315987 296580 316053 296581
rect 315987 296516 315988 296580
rect 316052 296516 316053 296580
rect 315987 296515 316053 296516
rect 315987 287196 316053 287197
rect 315987 287132 315988 287196
rect 316052 287132 316053 287196
rect 315987 287131 316053 287132
rect 315990 287061 316050 287131
rect 315987 287060 316053 287061
rect 315987 286996 315988 287060
rect 316052 286996 316053 287060
rect 315987 286995 316053 286996
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 316171 277540 316237 277541
rect 316171 277476 316172 277540
rect 316236 277476 316237 277540
rect 316171 277475 316237 277476
rect 316174 277410 316234 277475
rect 315990 277405 316234 277410
rect 315987 277404 316234 277405
rect 315987 277340 315988 277404
rect 316052 277350 316234 277404
rect 316052 277340 316053 277350
rect 315987 277339 316053 277340
rect 316171 267884 316237 267885
rect 316171 267820 316172 267884
rect 316236 267820 316237 267884
rect 316171 267819 316237 267820
rect 316174 267749 316234 267819
rect 316171 267748 316237 267749
rect 316171 267684 316172 267748
rect 316236 267684 316237 267748
rect 316171 267683 316237 267684
rect 315987 248436 316053 248437
rect 315987 248372 315988 248436
rect 316052 248430 316053 248436
rect 316052 248372 316234 248430
rect 315987 248371 316234 248372
rect 315990 248370 316234 248371
rect 316174 248301 316234 248370
rect 316171 248300 316237 248301
rect 316171 248236 316172 248300
rect 316236 248236 316237 248300
rect 316171 248235 316237 248236
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315987 238780 316053 238781
rect 315987 238716 315988 238780
rect 316052 238716 316053 238780
rect 315987 238715 316053 238716
rect 315990 238645 316050 238715
rect 315987 238644 316053 238645
rect 315987 238580 315988 238644
rect 316052 238580 316053 238644
rect 315987 238579 316053 238580
rect 316171 229124 316237 229125
rect 316171 229060 316172 229124
rect 316236 229060 316237 229124
rect 316171 229059 316237 229060
rect 316174 228989 316234 229059
rect 316171 228988 316237 228989
rect 316171 228924 316172 228988
rect 316236 228924 316237 228988
rect 316171 228923 316237 228924
rect 315987 219468 316053 219469
rect 315987 219404 315988 219468
rect 316052 219404 316053 219468
rect 315987 219403 316053 219404
rect 315990 219197 316050 219403
rect 315987 219196 316053 219197
rect 315987 219132 315988 219196
rect 316052 219132 316053 219196
rect 315987 219131 316053 219132
rect 315987 209812 316053 209813
rect 315987 209748 315988 209812
rect 316052 209748 316053 209812
rect 315987 209747 316053 209748
rect 315990 209541 316050 209747
rect 315987 209540 316053 209541
rect 315987 209476 315988 209540
rect 316052 209476 316053 209540
rect 315987 209475 316053 209476
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 312307 189684 312373 189685
rect 312307 189620 312308 189684
rect 312372 189620 312373 189684
rect 312307 189619 312373 189620
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 310467 116244 310533 116245
rect 310467 116180 310468 116244
rect 310532 116180 310533 116244
rect 310467 116179 310533 116180
rect 311514 97174 312134 132618
rect 312310 109173 312370 189619
rect 313227 188324 313293 188325
rect 313227 188260 313228 188324
rect 313292 188260 313293 188324
rect 313227 188259 313293 188260
rect 312307 109172 312373 109173
rect 312307 109108 312308 109172
rect 312372 109108 312373 109172
rect 312307 109107 312373 109108
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 309731 4044 309797 4045
rect 309731 3980 309732 4044
rect 309796 3980 309797 4044
rect 309731 3979 309797 3980
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 -3226 312134 24618
rect 313230 3501 313290 188259
rect 315234 172894 315854 208338
rect 315987 200156 316053 200157
rect 315987 200092 315988 200156
rect 316052 200092 316053 200156
rect 315987 200091 316053 200092
rect 315990 199885 316050 200091
rect 315987 199884 316053 199885
rect 315987 199820 315988 199884
rect 316052 199820 316053 199884
rect 315987 199819 316053 199820
rect 315987 190500 316053 190501
rect 315987 190436 315988 190500
rect 316052 190436 316053 190500
rect 315987 190435 316053 190436
rect 315990 190365 316050 190435
rect 315987 190364 316053 190365
rect 315987 190300 315988 190364
rect 316052 190300 316053 190364
rect 315987 190299 316053 190300
rect 316171 188460 316237 188461
rect 316171 188396 316172 188460
rect 316236 188396 316237 188460
rect 316171 188395 316237 188396
rect 315987 180980 316053 180981
rect 315987 180916 315988 180980
rect 316052 180916 316053 180980
rect 315987 180915 316053 180916
rect 315990 180709 316050 180915
rect 315987 180708 316053 180709
rect 315987 180644 315988 180708
rect 316052 180644 316053 180708
rect 315987 180643 316053 180644
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315987 171324 316053 171325
rect 315987 171260 315988 171324
rect 316052 171260 316053 171324
rect 315987 171259 316053 171260
rect 315990 171053 316050 171259
rect 315987 171052 316053 171053
rect 315987 170988 315988 171052
rect 316052 170988 316053 171052
rect 315987 170987 316053 170988
rect 315987 161668 316053 161669
rect 315987 161604 315988 161668
rect 316052 161604 316053 161668
rect 315987 161603 316053 161604
rect 315990 161261 316050 161603
rect 315987 161260 316053 161261
rect 315987 161196 315988 161260
rect 316052 161196 316053 161260
rect 315987 161195 316053 161196
rect 315987 151876 316053 151877
rect 315987 151812 315988 151876
rect 316052 151812 316053 151876
rect 315987 151811 316053 151812
rect 315990 151605 316050 151811
rect 315987 151604 316053 151605
rect 315987 151540 315988 151604
rect 316052 151540 316053 151604
rect 315987 151539 316053 151540
rect 315987 142220 316053 142221
rect 315987 142156 315988 142220
rect 316052 142156 316053 142220
rect 315987 142155 316053 142156
rect 315990 142085 316050 142155
rect 315987 142084 316053 142085
rect 315987 142020 315988 142084
rect 316052 142020 316053 142084
rect 315987 142019 316053 142020
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315987 132700 316053 132701
rect 315987 132636 315988 132700
rect 316052 132636 316053 132700
rect 315987 132635 316053 132636
rect 315990 132429 316050 132635
rect 315987 132428 316053 132429
rect 315987 132364 315988 132428
rect 316052 132364 316053 132428
rect 315987 132363 316053 132364
rect 315987 123044 316053 123045
rect 315987 122980 315988 123044
rect 316052 122980 316053 123044
rect 315987 122979 316053 122980
rect 315990 122773 316050 122979
rect 315987 122772 316053 122773
rect 315987 122708 315988 122772
rect 316052 122708 316053 122772
rect 315987 122707 316053 122708
rect 316174 102237 316234 188395
rect 316171 102236 316237 102237
rect 316171 102172 316172 102236
rect 316236 102172 316237 102236
rect 316171 102171 316237 102172
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 313227 3500 313293 3501
rect 313227 3436 313228 3500
rect 313292 3436 313293 3500
rect 313227 3435 313293 3436
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 -5146 315854 28338
rect 317462 11661 317522 358803
rect 318954 356614 319574 392058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 322979 360228 323045 360229
rect 322979 360164 322980 360228
rect 323044 360164 323045 360228
rect 322979 360163 323045 360164
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 320219 316708 320285 316709
rect 320219 316644 320220 316708
rect 320284 316644 320285 316708
rect 320219 316643 320285 316644
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 317459 11660 317525 11661
rect 317459 11596 317460 11660
rect 317524 11596 317525 11660
rect 317459 11595 317525 11596
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 320222 3501 320282 316643
rect 322059 306508 322125 306509
rect 322059 306444 322060 306508
rect 322124 306444 322125 306508
rect 322059 306443 322125 306444
rect 322062 4861 322122 306443
rect 322059 4860 322125 4861
rect 322059 4796 322060 4860
rect 322124 4796 322125 4860
rect 322059 4795 322125 4796
rect 322982 3501 323042 360163
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 320219 3500 320285 3501
rect 320219 3436 320220 3500
rect 320284 3436 320285 3500
rect 320219 3435 320285 3436
rect 322979 3500 323045 3501
rect 322979 3436 322980 3500
rect 323044 3436 323045 3500
rect 322979 3435 323045 3436
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 72721 579218 72957 579454
rect 72721 578898 72957 579134
rect 75686 561218 75922 561454
rect 75686 560898 75922 561134
rect 72721 543218 72957 543454
rect 72721 542898 72957 543134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 78651 579218 78887 579454
rect 78651 578898 78887 579134
rect 84582 579218 84818 579454
rect 84582 578898 84818 579134
rect 81617 561218 81853 561454
rect 81617 560898 81853 561134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 78651 543218 78887 543454
rect 78651 542898 78887 543134
rect 84582 543218 84818 543454
rect 84582 542898 84818 543134
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 73020 435218 73256 435454
rect 73020 434898 73256 435134
rect 88380 417218 88616 417454
rect 88380 416898 88616 417134
rect 73020 399218 73256 399454
rect 73020 398898 73256 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 103740 435218 103976 435454
rect 103740 434898 103976 435134
rect 103740 399218 103976 399454
rect 103740 398898 103976 399134
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 119100 417218 119336 417454
rect 119100 416898 119336 417134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 73020 291218 73256 291454
rect 73020 290898 73256 291134
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73020 255218 73256 255454
rect 73020 254898 73256 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 88380 309218 88616 309454
rect 88380 308898 88616 309134
rect 119100 309218 119336 309454
rect 119100 308898 119336 309134
rect 103740 291218 103976 291454
rect 103740 290898 103976 291134
rect 88380 273218 88616 273454
rect 88380 272898 88616 273134
rect 119100 273218 119336 273454
rect 119100 272898 119336 273134
rect 103740 255218 103976 255454
rect 103740 254898 103976 255134
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 134460 291218 134696 291454
rect 134460 290898 134696 291134
rect 134460 255218 134696 255454
rect 134460 254898 134696 255134
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149820 309218 150056 309454
rect 149820 308898 150056 309134
rect 149820 273218 150056 273454
rect 149820 272898 150056 273134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 69128 165218 69364 165454
rect 69128 164898 69364 165134
rect 164192 165218 164428 165454
rect 164192 164898 164428 165134
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 69128 129218 69364 129454
rect 69128 128898 69364 129134
rect 164192 129218 164428 129454
rect 164192 128898 164428 129134
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 204450 255218 204686 255454
rect 204450 254898 204686 255134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 219810 273218 220046 273454
rect 219810 272898 220046 273134
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 235170 255218 235406 255454
rect 235170 254898 235406 255134
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 256249 165218 256485 165454
rect 256249 164898 256485 165134
rect 259513 165218 259749 165454
rect 259513 164898 259749 165134
rect 254617 147218 254853 147454
rect 254617 146898 254853 147134
rect 257881 147218 258117 147454
rect 257881 146898 258117 147134
rect 261145 147218 261381 147454
rect 261145 146898 261381 147134
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 256249 129218 256485 129454
rect 256249 128898 256485 129134
rect 259513 129218 259749 129454
rect 259513 128898 259749 129134
rect 254617 111218 254853 111454
rect 254617 110898 254853 111134
rect 257881 111218 258117 111454
rect 257881 110898 258117 111134
rect 261145 111218 261381 111454
rect 261145 110898 261381 111134
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 294249 165218 294485 165454
rect 294249 164898 294485 165134
rect 297513 165218 297749 165454
rect 297513 164898 297749 165134
rect 292617 147218 292853 147454
rect 292617 146898 292853 147134
rect 295881 147218 296117 147454
rect 295881 146898 296117 147134
rect 299145 147218 299381 147454
rect 299145 146898 299381 147134
rect 294249 129218 294485 129454
rect 294249 128898 294485 129134
rect 297513 129218 297749 129454
rect 297513 128898 297749 129134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 292617 111218 292853 111454
rect 292617 110898 292853 111134
rect 295881 111218 296117 111454
rect 295881 110898 296117 111134
rect 299145 111218 299381 111454
rect 299145 110898 299381 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 72721 579454
rect 72957 579218 78651 579454
rect 78887 579218 84582 579454
rect 84818 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 72721 579134
rect 72957 578898 78651 579134
rect 78887 578898 84582 579134
rect 84818 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 75686 561454
rect 75922 561218 81617 561454
rect 81853 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 75686 561134
rect 75922 560898 81617 561134
rect 81853 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 72721 543454
rect 72957 543218 78651 543454
rect 78887 543218 84582 543454
rect 84818 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 72721 543134
rect 72957 542898 78651 543134
rect 78887 542898 84582 543134
rect 84818 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73020 435454
rect 73256 435218 103740 435454
rect 103976 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73020 435134
rect 73256 434898 103740 435134
rect 103976 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 88380 417454
rect 88616 417218 119100 417454
rect 119336 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 88380 417134
rect 88616 416898 119100 417134
rect 119336 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73020 399454
rect 73256 399218 103740 399454
rect 103976 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73020 399134
rect 73256 398898 103740 399134
rect 103976 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 88380 309454
rect 88616 309218 119100 309454
rect 119336 309218 149820 309454
rect 150056 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 88380 309134
rect 88616 308898 119100 309134
rect 119336 308898 149820 309134
rect 150056 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73020 291454
rect 73256 291218 103740 291454
rect 103976 291218 134460 291454
rect 134696 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73020 291134
rect 73256 290898 103740 291134
rect 103976 290898 134460 291134
rect 134696 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 88380 273454
rect 88616 273218 119100 273454
rect 119336 273218 149820 273454
rect 150056 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 219810 273454
rect 220046 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 88380 273134
rect 88616 272898 119100 273134
rect 119336 272898 149820 273134
rect 150056 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 219810 273134
rect 220046 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73020 255454
rect 73256 255218 103740 255454
rect 103976 255218 134460 255454
rect 134696 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 204450 255454
rect 204686 255218 235170 255454
rect 235406 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73020 255134
rect 73256 254898 103740 255134
rect 103976 254898 134460 255134
rect 134696 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 204450 255134
rect 204686 254898 235170 255134
rect 235406 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 69128 165454
rect 69364 165218 164192 165454
rect 164428 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 256249 165454
rect 256485 165218 259513 165454
rect 259749 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 294249 165454
rect 294485 165218 297513 165454
rect 297749 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 69128 165134
rect 69364 164898 164192 165134
rect 164428 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 256249 165134
rect 256485 164898 259513 165134
rect 259749 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 294249 165134
rect 294485 164898 297513 165134
rect 297749 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 254617 147454
rect 254853 147218 257881 147454
rect 258117 147218 261145 147454
rect 261381 147218 292617 147454
rect 292853 147218 295881 147454
rect 296117 147218 299145 147454
rect 299381 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 254617 147134
rect 254853 146898 257881 147134
rect 258117 146898 261145 147134
rect 261381 146898 292617 147134
rect 292853 146898 295881 147134
rect 296117 146898 299145 147134
rect 299381 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 69128 129454
rect 69364 129218 164192 129454
rect 164428 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 256249 129454
rect 256485 129218 259513 129454
rect 259749 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 294249 129454
rect 294485 129218 297513 129454
rect 297749 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 69128 129134
rect 69364 128898 164192 129134
rect 164428 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 256249 129134
rect 256485 128898 259513 129134
rect 259749 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 294249 129134
rect 294485 128898 297513 129134
rect 297749 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 254617 111454
rect 254853 111218 257881 111454
rect 258117 111218 261145 111454
rect 261381 111218 292617 111454
rect 292853 111218 295881 111454
rect 296117 111218 299145 111454
rect 299381 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 254617 111134
rect 254853 110898 257881 111134
rect 258117 110898 261145 111134
rect 261381 110898 292617 111134
rect 292853 110898 295881 111134
rect 296117 110898 299145 111134
rect 299381 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use wrapped_spell  wrapped_spell_1
timestamp 1640163700
transform 1 0 68770 0 1 241592
box 0 0 86000 86000
use wrapped_ppm_decoder  wrapped_ppm_decoder_3
timestamp 1640163700
transform 1 0 68770 0 1 539166
box 0 0 20000 50000
use wrapped_ppm_coder  wrapped_ppm_coder_2
timestamp 1640163700
transform 1 0 68770 0 1 390356
box 0 0 51907 54051
use wrapped_function_generator  wrapped_function_generator_0
timestamp 1640163700
transform 1 0 200200 0 1 240182
box 0 0 44000 44000
use wb_openram_wrapper  wb_openram_wrapper
timestamp 1640163700
transform 1 0 252000 0 1 96000
box 0 144 12000 79688
use wb_bridge_2way  wb_bridge_2way
timestamp 1640163700
transform 1 0 290000 0 1 96000
box 0 0 12000 79688
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 1640163700
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 94000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 94000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 238182 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 176600 74414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 176600 110414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 176600 146414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 329592 74414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 329592 110414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 446407 74414 537166 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 591166 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 446407 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 329592 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 286182 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 178000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 178000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 94000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 94000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 238182 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 176600 78134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 176600 114134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 176600 150134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 329592 78134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 329592 114134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 446407 78134 537166 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 591166 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 446407 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 329592 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 286182 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 178000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 178000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 94000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 94000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 238182 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 176600 81854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 176600 117854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 176600 153854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 329592 81854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 329592 117854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 446407 81854 537166 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 591166 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 446407 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 329592 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 286182 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 178000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 178000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 94000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 94000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 238182 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 176600 85574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 176600 121574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 329592 85574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 329592 121574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 446407 85574 537166 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 591166 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 446407 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 176600 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 286182 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 178000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 178000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 238182 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 238182 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 176600 99854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 176600 135854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 329592 99854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 446407 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 329592 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 286182 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 286182 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 238182 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 176600 67574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 176600 103574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 176600 139574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 329592 67574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 329592 103574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 446407 67574 537166 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 591166 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 446407 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 329592 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 286182 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 238182 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 238182 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 176600 92414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 176600 128414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 329592 92414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 446407 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 329592 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 176600 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 286182 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 286182 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 238182 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 238182 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 176600 96134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 176600 132134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 329592 96134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 446407 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 329592 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 286182 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 286182 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
