magic
tech sky130A
magscale 1 2
timestamp 1640773853
<< metal1 >>
rect 62022 702992 62028 703044
rect 62080 703032 62086 703044
rect 267642 703032 267648 703044
rect 62080 703004 267648 703032
rect 62080 702992 62086 703004
rect 267642 702992 267648 703004
rect 267700 702992 267706 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 169754 702924 169760 702976
rect 169812 702964 169818 702976
rect 170306 702964 170312 702976
rect 169812 702936 170312 702964
rect 169812 702924 169818 702936
rect 170306 702924 170312 702936
rect 170364 702964 170370 702976
rect 281534 702964 281540 702976
rect 170364 702936 281540 702964
rect 170364 702924 170370 702936
rect 281534 702924 281540 702936
rect 281592 702924 281598 702976
rect 283834 702924 283840 702976
rect 283892 702964 283898 702976
rect 351914 702964 351920 702976
rect 283892 702936 351920 702964
rect 283892 702924 283898 702936
rect 351914 702924 351920 702936
rect 351972 702924 351978 702976
rect 202782 702856 202788 702908
rect 202840 702896 202846 702908
rect 273254 702896 273260 702908
rect 202840 702868 273260 702896
rect 202840 702856 202846 702868
rect 273254 702856 273260 702868
rect 273312 702856 273318 702908
rect 276014 702856 276020 702908
rect 276072 702896 276078 702908
rect 478506 702896 478512 702908
rect 276072 702868 478512 702896
rect 276072 702856 276078 702868
rect 478506 702856 478512 702868
rect 478564 702856 478570 702908
rect 130378 702788 130384 702840
rect 130436 702828 130442 702840
rect 218974 702828 218980 702840
rect 130436 702800 218980 702828
rect 130436 702788 130442 702800
rect 218974 702788 218980 702800
rect 219032 702788 219038 702840
rect 349798 702788 349804 702840
rect 349856 702828 349862 702840
rect 494790 702828 494796 702840
rect 349856 702800 494796 702828
rect 349856 702788 349862 702800
rect 494790 702788 494796 702800
rect 494848 702788 494854 702840
rect 233878 702720 233884 702772
rect 233936 702760 233942 702772
rect 397362 702760 397368 702772
rect 233936 702732 397368 702760
rect 233936 702720 233942 702732
rect 397362 702720 397368 702732
rect 397420 702720 397426 702772
rect 67634 702652 67640 702704
rect 67692 702692 67698 702704
rect 169754 702692 169760 702704
rect 67692 702664 169760 702692
rect 67692 702652 67698 702664
rect 169754 702652 169760 702664
rect 169812 702652 169818 702704
rect 197262 702652 197268 702704
rect 197320 702692 197326 702704
rect 364978 702692 364984 702704
rect 197320 702664 364984 702692
rect 197320 702652 197326 702664
rect 364978 702652 364984 702664
rect 365036 702652 365042 702704
rect 381538 702652 381544 702704
rect 381596 702692 381602 702704
rect 462314 702692 462320 702704
rect 381596 702664 462320 702692
rect 381596 702652 381602 702664
rect 462314 702652 462320 702664
rect 462372 702652 462378 702704
rect 24302 702584 24308 702636
rect 24360 702624 24366 702636
rect 79318 702624 79324 702636
rect 24360 702596 79324 702624
rect 24360 702584 24366 702596
rect 79318 702584 79324 702596
rect 79376 702584 79382 702636
rect 95142 702584 95148 702636
rect 95200 702624 95206 702636
rect 300118 702624 300124 702636
rect 95200 702596 300124 702624
rect 95200 702584 95206 702596
rect 300118 702584 300124 702596
rect 300176 702624 300182 702636
rect 356146 702624 356152 702636
rect 300176 702596 356152 702624
rect 300176 702584 300182 702596
rect 356146 702584 356152 702596
rect 356204 702584 356210 702636
rect 360838 702584 360844 702636
rect 360896 702624 360902 702636
rect 543458 702624 543464 702636
rect 360896 702596 543464 702624
rect 360896 702584 360902 702596
rect 543458 702584 543464 702596
rect 543516 702584 543522 702636
rect 88242 702516 88248 702568
rect 88300 702556 88306 702568
rect 235166 702556 235172 702568
rect 88300 702528 235172 702556
rect 88300 702516 88306 702528
rect 235166 702516 235172 702528
rect 235224 702516 235230 702568
rect 264238 702516 264244 702568
rect 264296 702556 264302 702568
rect 559650 702556 559656 702568
rect 264296 702528 559656 702556
rect 264296 702516 264302 702528
rect 559650 702516 559656 702528
rect 559708 702516 559714 702568
rect 8110 702448 8116 702500
rect 8168 702488 8174 702500
rect 88794 702488 88800 702500
rect 8168 702460 88800 702488
rect 8168 702448 8174 702460
rect 88794 702448 88800 702460
rect 88852 702448 88858 702500
rect 93762 702448 93768 702500
rect 93820 702488 93826 702500
rect 527174 702488 527180 702500
rect 93820 702460 527180 702488
rect 93820 702448 93826 702460
rect 527174 702448 527180 702460
rect 527232 702448 527238 702500
rect 75178 700272 75184 700324
rect 75236 700312 75242 700324
rect 105446 700312 105452 700324
rect 75236 700284 105452 700312
rect 75236 700272 75242 700284
rect 105446 700272 105452 700284
rect 105504 700272 105510 700324
rect 124858 700272 124864 700324
rect 124916 700312 124922 700324
rect 137830 700312 137836 700324
rect 124916 700284 137836 700312
rect 124916 700272 124922 700284
rect 137830 700272 137836 700284
rect 137888 700272 137894 700324
rect 327718 700272 327724 700324
rect 327776 700312 327782 700324
rect 348786 700312 348792 700324
rect 327776 700284 348792 700312
rect 327776 700272 327782 700284
rect 348786 700272 348792 700284
rect 348844 700272 348850 700324
rect 376110 700272 376116 700324
rect 376168 700312 376174 700324
rect 429838 700312 429844 700324
rect 376168 700284 429844 700312
rect 376168 700272 376174 700284
rect 429838 700272 429844 700284
rect 429896 700272 429902 700324
rect 66162 699660 66168 699712
rect 66220 699700 66226 699712
rect 72970 699700 72976 699712
rect 66220 699672 72976 699700
rect 66220 699660 66226 699672
rect 72970 699660 72976 699672
rect 73028 699660 73034 699712
rect 86862 699660 86868 699712
rect 86920 699700 86926 699712
rect 89162 699700 89168 699712
rect 86920 699672 89168 699700
rect 86920 699660 86926 699672
rect 89162 699660 89168 699672
rect 89220 699660 89226 699712
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 14458 670732 14464 670744
rect 3568 670704 14464 670732
rect 3568 670692 3574 670704
rect 14458 670692 14464 670704
rect 14516 670692 14522 670744
rect 2774 656956 2780 657008
rect 2832 656996 2838 657008
rect 4798 656996 4804 657008
rect 2832 656968 4804 656996
rect 2832 656956 2838 656968
rect 4798 656956 4804 656968
rect 4856 656956 4862 657008
rect 3510 632068 3516 632120
rect 3568 632108 3574 632120
rect 21358 632108 21364 632120
rect 3568 632080 21364 632108
rect 3568 632068 3574 632080
rect 21358 632068 21364 632080
rect 21416 632068 21422 632120
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 22738 618304 22744 618316
rect 3568 618276 22744 618304
rect 3568 618264 3574 618276
rect 22738 618264 22744 618276
rect 22796 618264 22802 618316
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 90358 605860 90364 605872
rect 3568 605832 90364 605860
rect 3568 605820 3574 605832
rect 90358 605820 90364 605832
rect 90416 605820 90422 605872
rect 67450 598952 67456 599004
rect 67508 598992 67514 599004
rect 259454 598992 259460 599004
rect 67508 598964 259460 598992
rect 67508 598952 67514 598964
rect 259454 598952 259460 598964
rect 259512 598952 259518 599004
rect 82814 597524 82820 597576
rect 82872 597564 82878 597576
rect 111150 597564 111156 597576
rect 82872 597536 111156 597564
rect 82872 597524 82878 597536
rect 111150 597524 111156 597536
rect 111208 597524 111214 597576
rect 79962 596776 79968 596828
rect 80020 596816 80026 596828
rect 86862 596816 86868 596828
rect 80020 596788 86868 596816
rect 80020 596776 80026 596788
rect 86862 596776 86868 596788
rect 86920 596816 86926 596828
rect 92474 596816 92480 596828
rect 86920 596788 92480 596816
rect 86920 596776 86926 596788
rect 92474 596776 92480 596788
rect 92532 596776 92538 596828
rect 70302 596164 70308 596216
rect 70360 596204 70366 596216
rect 349798 596204 349804 596216
rect 70360 596176 349804 596204
rect 70360 596164 70366 596176
rect 349798 596164 349804 596176
rect 349856 596164 349862 596216
rect 85942 594804 85948 594856
rect 86000 594844 86006 594856
rect 155218 594844 155224 594856
rect 86000 594816 155224 594844
rect 86000 594804 86006 594816
rect 155218 594804 155224 594816
rect 155276 594804 155282 594856
rect 40034 594056 40040 594108
rect 40092 594096 40098 594108
rect 89806 594096 89812 594108
rect 40092 594068 89812 594096
rect 40092 594056 40098 594068
rect 89806 594056 89812 594068
rect 89864 594056 89870 594108
rect 90358 593784 90364 593836
rect 90416 593824 90422 593836
rect 91186 593824 91192 593836
rect 90416 593796 91192 593824
rect 90416 593784 90422 593796
rect 91186 593784 91192 593796
rect 91244 593784 91250 593836
rect 88242 593376 88248 593428
rect 88300 593416 88306 593428
rect 113174 593416 113180 593428
rect 88300 593388 113180 593416
rect 88300 593376 88306 593388
rect 113174 593376 113180 593388
rect 113232 593376 113238 593428
rect 67358 592628 67364 592680
rect 67416 592668 67422 592680
rect 75178 592668 75184 592680
rect 67416 592640 75184 592668
rect 67416 592628 67422 592640
rect 75178 592628 75184 592640
rect 75236 592628 75242 592680
rect 75638 592084 75644 592136
rect 75696 592124 75702 592136
rect 96614 592124 96620 592136
rect 75696 592096 96620 592124
rect 75696 592084 75702 592096
rect 96614 592084 96620 592096
rect 96672 592084 96678 592136
rect 84102 592016 84108 592068
rect 84160 592056 84166 592068
rect 111794 592056 111800 592068
rect 84160 592028 111800 592056
rect 84160 592016 84166 592028
rect 111794 592016 111800 592028
rect 111852 592016 111858 592068
rect 79318 591472 79324 591524
rect 79376 591512 79382 591524
rect 80698 591512 80704 591524
rect 79376 591484 80704 591512
rect 79376 591472 79382 591484
rect 80698 591472 80704 591484
rect 80756 591472 80762 591524
rect 4798 591268 4804 591320
rect 4856 591308 4862 591320
rect 69106 591308 69112 591320
rect 4856 591280 69112 591308
rect 4856 591268 4862 591280
rect 69106 591268 69112 591280
rect 69164 591268 69170 591320
rect 72142 590792 72148 590844
rect 72200 590832 72206 590844
rect 79962 590832 79968 590844
rect 72200 590804 79968 590832
rect 72200 590792 72206 590804
rect 79962 590792 79968 590804
rect 80020 590792 80026 590844
rect 69106 590724 69112 590776
rect 69164 590764 69170 590776
rect 71682 590764 71688 590776
rect 69164 590736 71688 590764
rect 69164 590724 69170 590736
rect 71682 590724 71688 590736
rect 71740 590724 71746 590776
rect 78582 590724 78588 590776
rect 78640 590764 78646 590776
rect 93118 590764 93124 590776
rect 78640 590736 93124 590764
rect 78640 590724 78646 590736
rect 93118 590724 93124 590736
rect 93176 590724 93182 590776
rect 70118 590656 70124 590708
rect 70176 590696 70182 590708
rect 74442 590696 74448 590708
rect 70176 590668 74448 590696
rect 70176 590656 70182 590668
rect 74442 590656 74448 590668
rect 74500 590656 74506 590708
rect 85022 590656 85028 590708
rect 85080 590696 85086 590708
rect 88242 590696 88248 590708
rect 85080 590668 88248 590696
rect 85080 590656 85086 590668
rect 88242 590656 88248 590668
rect 88300 590656 88306 590708
rect 71682 589976 71688 590028
rect 71740 590016 71746 590028
rect 89070 590016 89076 590028
rect 71740 589988 89076 590016
rect 71740 589976 71746 589988
rect 89070 589976 89076 589988
rect 89128 589976 89134 590028
rect 74902 589908 74908 589960
rect 74960 589948 74966 589960
rect 75638 589948 75644 589960
rect 74960 589920 75644 589948
rect 74960 589908 74966 589920
rect 75638 589908 75644 589920
rect 75696 589908 75702 589960
rect 80698 589908 80704 589960
rect 80756 589948 80762 589960
rect 106918 589948 106924 589960
rect 80756 589920 106924 589948
rect 80756 589908 80762 589920
rect 106918 589908 106924 589920
rect 106976 589908 106982 589960
rect 7558 589296 7564 589348
rect 7616 589336 7622 589348
rect 74902 589336 74908 589348
rect 7616 589308 74908 589336
rect 7616 589296 7622 589308
rect 74902 589296 74908 589308
rect 74960 589296 74966 589348
rect 81894 588548 81900 588600
rect 81952 588588 81958 588600
rect 94498 588588 94504 588600
rect 81952 588560 94504 588588
rect 81952 588548 81958 588560
rect 94498 588548 94504 588560
rect 94556 588548 94562 588600
rect 76098 588412 76104 588464
rect 76156 588412 76162 588464
rect 76116 588180 76144 588412
rect 88978 588180 88984 588192
rect 76116 588152 88984 588180
rect 88978 588140 88984 588152
rect 89036 588140 89042 588192
rect 70366 587948 71774 587976
rect 55122 587868 55128 587920
rect 55180 587908 55186 587920
rect 66806 587908 66812 587920
rect 55180 587880 66812 587908
rect 55180 587868 55186 587880
rect 66806 587868 66812 587880
rect 66864 587868 66870 587920
rect 67542 587868 67548 587920
rect 67600 587908 67606 587920
rect 70366 587908 70394 587948
rect 67600 587880 70394 587908
rect 67600 587868 67606 587880
rect 71746 587704 71774 587948
rect 351914 587908 351920 587920
rect 80026 587880 351920 587908
rect 80026 587704 80054 587880
rect 351914 587868 351920 587880
rect 351972 587868 351978 587920
rect 71746 587676 80054 587704
rect 88794 587120 88800 587172
rect 88852 587160 88858 587172
rect 115198 587160 115204 587172
rect 88852 587132 115204 587160
rect 88852 587120 88858 587132
rect 115198 587120 115204 587132
rect 115256 587120 115262 587172
rect 88978 586576 88984 586628
rect 89036 586616 89042 586628
rect 98730 586616 98736 586628
rect 89036 586588 98736 586616
rect 89036 586576 89042 586588
rect 98730 586576 98736 586588
rect 98788 586576 98794 586628
rect 59078 586508 59084 586560
rect 59136 586548 59142 586560
rect 66254 586548 66260 586560
rect 59136 586520 66260 586548
rect 59136 586508 59142 586520
rect 66254 586508 66260 586520
rect 66312 586508 66318 586560
rect 57882 585148 57888 585200
rect 57940 585188 57946 585200
rect 66898 585188 66904 585200
rect 57940 585160 66904 585188
rect 57940 585148 57946 585160
rect 66898 585148 66904 585160
rect 66956 585148 66962 585200
rect 91278 584400 91284 584452
rect 91336 584440 91342 584452
rect 95142 584440 95148 584452
rect 91336 584412 95148 584440
rect 91336 584400 91342 584412
rect 95142 584400 95148 584412
rect 95200 584440 95206 584452
rect 128354 584440 128360 584452
rect 95200 584412 128360 584440
rect 95200 584400 95206 584412
rect 128354 584400 128360 584412
rect 128412 584400 128418 584452
rect 93762 583720 93768 583772
rect 93820 583760 93826 583772
rect 116578 583760 116584 583772
rect 93820 583732 116584 583760
rect 93820 583720 93854 583732
rect 116578 583720 116584 583732
rect 116636 583720 116642 583772
rect 91830 583652 91836 583704
rect 91888 583692 91894 583704
rect 93826 583692 93854 583720
rect 91888 583664 93854 583692
rect 91888 583652 91894 583664
rect 50890 582360 50896 582412
rect 50948 582400 50954 582412
rect 66806 582400 66812 582412
rect 50948 582372 66812 582400
rect 50948 582360 50954 582372
rect 66806 582360 66812 582372
rect 66864 582360 66870 582412
rect 64690 581000 64696 581052
rect 64748 581040 64754 581052
rect 66530 581040 66536 581052
rect 64748 581012 66536 581040
rect 64748 581000 64754 581012
rect 66530 581000 66536 581012
rect 66588 581000 66594 581052
rect 91278 581000 91284 581052
rect 91336 581040 91342 581052
rect 108298 581040 108304 581052
rect 91336 581012 108304 581040
rect 91336 581000 91342 581012
rect 108298 581000 108304 581012
rect 108356 581000 108362 581052
rect 3050 580728 3056 580780
rect 3108 580768 3114 580780
rect 7558 580768 7564 580780
rect 3108 580740 7564 580768
rect 3108 580728 3114 580740
rect 7558 580728 7564 580740
rect 7616 580728 7622 580780
rect 61930 579640 61936 579692
rect 61988 579680 61994 579692
rect 66806 579680 66812 579692
rect 61988 579652 66812 579680
rect 61988 579640 61994 579652
rect 66806 579640 66812 579652
rect 66864 579640 66870 579692
rect 91278 576852 91284 576904
rect 91336 576892 91342 576904
rect 111058 576892 111064 576904
rect 91336 576864 111064 576892
rect 91336 576852 91342 576864
rect 111058 576852 111064 576864
rect 111116 576852 111122 576904
rect 21358 576104 21364 576156
rect 21416 576144 21422 576156
rect 39942 576144 39948 576156
rect 21416 576116 39948 576144
rect 21416 576104 21422 576116
rect 39942 576104 39948 576116
rect 40000 576104 40006 576156
rect 91186 576104 91192 576156
rect 91244 576144 91250 576156
rect 122834 576144 122840 576156
rect 91244 576116 122840 576144
rect 91244 576104 91250 576116
rect 122834 576104 122840 576116
rect 122892 576104 122898 576156
rect 39942 575492 39948 575544
rect 40000 575532 40006 575544
rect 66806 575532 66812 575544
rect 40000 575504 66812 575532
rect 40000 575492 40006 575504
rect 66806 575492 66812 575504
rect 66864 575492 66870 575544
rect 93118 574744 93124 574796
rect 93176 574784 93182 574796
rect 103514 574784 103520 574796
rect 93176 574756 103520 574784
rect 93176 574744 93182 574756
rect 103514 574744 103520 574756
rect 103572 574744 103578 574796
rect 104158 574132 104164 574184
rect 104216 574172 104222 574184
rect 109678 574172 109684 574184
rect 104216 574144 109684 574172
rect 104216 574132 104222 574144
rect 109678 574132 109684 574144
rect 109736 574132 109742 574184
rect 61838 574064 61844 574116
rect 61896 574104 61902 574116
rect 67358 574104 67364 574116
rect 61896 574076 67364 574104
rect 61896 574064 61902 574076
rect 67358 574064 67364 574076
rect 67416 574064 67422 574116
rect 91738 574064 91744 574116
rect 91796 574104 91802 574116
rect 136634 574104 136640 574116
rect 91796 574076 136640 574104
rect 91796 574064 91802 574076
rect 136634 574064 136640 574076
rect 136692 574064 136698 574116
rect 91738 572704 91744 572756
rect 91796 572744 91802 572756
rect 112438 572744 112444 572756
rect 91796 572716 112444 572744
rect 91796 572704 91802 572716
rect 112438 572704 112444 572716
rect 112496 572704 112502 572756
rect 91186 571412 91192 571464
rect 91244 571452 91250 571464
rect 94590 571452 94596 571464
rect 91244 571424 94596 571452
rect 91244 571412 91250 571424
rect 94590 571412 94596 571424
rect 94648 571412 94654 571464
rect 63310 571344 63316 571396
rect 63368 571384 63374 571396
rect 66806 571384 66812 571396
rect 63368 571356 66812 571384
rect 63368 571344 63374 571356
rect 66806 571344 66812 571356
rect 66864 571344 66870 571396
rect 91738 571344 91744 571396
rect 91796 571384 91802 571396
rect 122190 571384 122196 571396
rect 91796 571356 122196 571384
rect 91796 571344 91802 571356
rect 122190 571344 122196 571356
rect 122248 571344 122254 571396
rect 174538 569916 174544 569968
rect 174596 569956 174602 569968
rect 341518 569956 341524 569968
rect 174596 569928 341524 569956
rect 174596 569916 174602 569928
rect 341518 569916 341524 569928
rect 341576 569916 341582 569968
rect 48130 569168 48136 569220
rect 48188 569208 48194 569220
rect 67082 569208 67088 569220
rect 48188 569180 67088 569208
rect 48188 569168 48194 569180
rect 67082 569168 67088 569180
rect 67140 569168 67146 569220
rect 177942 568556 177948 568608
rect 178000 568596 178006 568608
rect 320174 568596 320180 568608
rect 178000 568568 320180 568596
rect 178000 568556 178006 568568
rect 320174 568556 320180 568568
rect 320232 568556 320238 568608
rect 64782 567196 64788 567248
rect 64840 567236 64846 567248
rect 66806 567236 66812 567248
rect 64840 567208 66812 567236
rect 64840 567196 64846 567208
rect 66806 567196 66812 567208
rect 66864 567196 66870 567248
rect 89806 567196 89812 567248
rect 89864 567236 89870 567248
rect 133138 567236 133144 567248
rect 89864 567208 133144 567236
rect 89864 567196 89870 567208
rect 133138 567196 133144 567208
rect 133196 567196 133202 567248
rect 155862 567196 155868 567248
rect 155920 567236 155926 567248
rect 311894 567236 311900 567248
rect 155920 567208 311900 567236
rect 155920 567196 155926 567208
rect 311894 567196 311900 567208
rect 311952 567196 311958 567248
rect 94590 566448 94596 566500
rect 94648 566488 94654 566500
rect 138014 566488 138020 566500
rect 94648 566460 138020 566488
rect 94648 566448 94654 566460
rect 138014 566448 138020 566460
rect 138072 566448 138078 566500
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 43438 565876 43444 565888
rect 3292 565848 43444 565876
rect 3292 565836 3298 565848
rect 43438 565836 43444 565848
rect 43496 565836 43502 565888
rect 53650 565836 53656 565888
rect 53708 565876 53714 565888
rect 67634 565876 67640 565888
rect 53708 565848 67640 565876
rect 53708 565836 53714 565848
rect 67634 565836 67640 565848
rect 67692 565836 67698 565888
rect 91554 565836 91560 565888
rect 91612 565876 91618 565888
rect 116670 565876 116676 565888
rect 91612 565848 116676 565876
rect 91612 565836 91618 565848
rect 116670 565836 116676 565848
rect 116728 565836 116734 565888
rect 138014 565836 138020 565888
rect 138072 565876 138078 565888
rect 213914 565876 213920 565888
rect 138072 565848 213920 565876
rect 138072 565836 138078 565848
rect 213914 565836 213920 565848
rect 213972 565836 213978 565888
rect 93118 565088 93124 565140
rect 93176 565128 93182 565140
rect 133874 565128 133880 565140
rect 93176 565100 133880 565128
rect 93176 565088 93182 565100
rect 133874 565088 133880 565100
rect 133932 565128 133938 565140
rect 135162 565128 135168 565140
rect 133932 565100 135168 565128
rect 133932 565088 133938 565100
rect 135162 565088 135168 565100
rect 135220 565088 135226 565140
rect 55858 564408 55864 564460
rect 55916 564448 55922 564460
rect 66806 564448 66812 564460
rect 55916 564420 66812 564448
rect 55916 564408 55922 564420
rect 66806 564408 66812 564420
rect 66864 564408 66870 564460
rect 91554 564408 91560 564460
rect 91612 564448 91618 564460
rect 107010 564448 107016 564460
rect 91612 564420 107016 564448
rect 91612 564408 91618 564420
rect 107010 564408 107016 564420
rect 107068 564408 107074 564460
rect 135162 564408 135168 564460
rect 135220 564448 135226 564460
rect 291194 564448 291200 564460
rect 135220 564420 291200 564448
rect 135220 564408 135226 564420
rect 291194 564408 291200 564420
rect 291252 564408 291258 564460
rect 52270 563048 52276 563100
rect 52328 563088 52334 563100
rect 66806 563088 66812 563100
rect 52328 563060 66812 563088
rect 52328 563048 52334 563060
rect 66806 563048 66812 563060
rect 66864 563048 66870 563100
rect 91554 563048 91560 563100
rect 91612 563088 91618 563100
rect 106182 563088 106188 563100
rect 91612 563060 106188 563088
rect 91612 563048 91618 563060
rect 106182 563048 106188 563060
rect 106240 563048 106246 563100
rect 191098 563048 191104 563100
rect 191156 563088 191162 563100
rect 357434 563088 357440 563100
rect 191156 563060 357440 563088
rect 191156 563048 191162 563060
rect 357434 563048 357440 563060
rect 357492 563048 357498 563100
rect 106182 562300 106188 562352
rect 106240 562340 106246 562352
rect 197354 562340 197360 562352
rect 106240 562312 197360 562340
rect 106240 562300 106246 562312
rect 197354 562300 197360 562312
rect 197412 562300 197418 562352
rect 197354 561756 197360 561808
rect 197412 561796 197418 561808
rect 241514 561796 241520 561808
rect 197412 561768 241520 561796
rect 197412 561756 197418 561768
rect 241514 561756 241520 561768
rect 241572 561756 241578 561808
rect 37182 561688 37188 561740
rect 37240 561728 37246 561740
rect 66806 561728 66812 561740
rect 37240 561700 66812 561728
rect 37240 561688 37246 561700
rect 66806 561688 66812 561700
rect 66864 561688 66870 561740
rect 186958 561688 186964 561740
rect 187016 561728 187022 561740
rect 267734 561728 267740 561740
rect 187016 561700 267740 561728
rect 187016 561688 187022 561700
rect 267734 561688 267740 561700
rect 267792 561688 267798 561740
rect 263594 561620 263600 561672
rect 263652 561660 263658 561672
rect 264238 561660 264244 561672
rect 263652 561632 264244 561660
rect 263652 561620 263658 561632
rect 264238 561620 264244 561632
rect 264296 561620 264302 561672
rect 178678 560328 178684 560380
rect 178736 560368 178742 560380
rect 263594 560368 263600 560380
rect 178736 560340 263600 560368
rect 178736 560328 178742 560340
rect 263594 560328 263600 560340
rect 263652 560328 263658 560380
rect 41322 560260 41328 560312
rect 41380 560300 41386 560312
rect 66806 560300 66812 560312
rect 41380 560272 66812 560300
rect 41380 560260 41386 560272
rect 66806 560260 66812 560272
rect 66864 560260 66870 560312
rect 111150 560260 111156 560312
rect 111208 560300 111214 560312
rect 111702 560300 111708 560312
rect 111208 560272 111708 560300
rect 111208 560260 111214 560272
rect 111702 560260 111708 560272
rect 111760 560300 111766 560312
rect 358998 560300 359004 560312
rect 111760 560272 359004 560300
rect 111760 560260 111766 560272
rect 358998 560260 359004 560272
rect 359056 560260 359062 560312
rect 133138 560192 133144 560244
rect 133196 560232 133202 560244
rect 133782 560232 133788 560244
rect 133196 560204 133788 560232
rect 133196 560192 133202 560204
rect 133782 560192 133788 560204
rect 133840 560192 133846 560244
rect 133782 558968 133788 559020
rect 133840 559008 133846 559020
rect 209774 559008 209780 559020
rect 133840 558980 209780 559008
rect 133840 558968 133846 558980
rect 209774 558968 209780 558980
rect 209832 558968 209838 559020
rect 89622 558900 89628 558952
rect 89680 558940 89686 558952
rect 129734 558940 129740 558952
rect 89680 558912 129740 558940
rect 89680 558900 89686 558912
rect 129734 558900 129740 558912
rect 129792 558900 129798 558952
rect 195882 558900 195888 558952
rect 195940 558940 195946 558952
rect 288434 558940 288440 558952
rect 195940 558912 288440 558940
rect 195940 558900 195946 558912
rect 288434 558900 288440 558912
rect 288492 558900 288498 558952
rect 59170 558288 59176 558340
rect 59228 558328 59234 558340
rect 62022 558328 62028 558340
rect 59228 558300 62028 558328
rect 59228 558288 59234 558300
rect 62022 558288 62028 558300
rect 62080 558288 62086 558340
rect 97258 558152 97264 558204
rect 97316 558192 97322 558204
rect 118510 558192 118516 558204
rect 97316 558164 118516 558192
rect 97316 558152 97322 558164
rect 118510 558152 118516 558164
rect 118568 558152 118574 558204
rect 198642 558152 198648 558204
rect 198700 558192 198706 558204
rect 582466 558192 582472 558204
rect 198700 558164 582472 558192
rect 198700 558152 198706 558164
rect 582466 558152 582472 558164
rect 582524 558152 582530 558204
rect 62022 557540 62028 557592
rect 62080 557580 62086 557592
rect 66806 557580 66812 557592
rect 62080 557552 66812 557580
rect 62080 557540 62086 557552
rect 66806 557540 66812 557552
rect 66864 557540 66870 557592
rect 188338 557540 188344 557592
rect 188396 557580 188402 557592
rect 268378 557580 268384 557592
rect 188396 557552 268384 557580
rect 188396 557540 188402 557552
rect 268378 557540 268384 557552
rect 268436 557540 268442 557592
rect 91094 557472 91100 557524
rect 91152 557512 91158 557524
rect 91278 557512 91284 557524
rect 91152 557484 91284 557512
rect 91152 557472 91158 557484
rect 91278 557472 91284 557484
rect 91336 557472 91342 557524
rect 92290 556792 92296 556844
rect 92348 556832 92354 556844
rect 148410 556832 148416 556844
rect 92348 556804 148416 556832
rect 92348 556792 92354 556804
rect 148410 556792 148416 556804
rect 148468 556792 148474 556844
rect 180150 556248 180156 556300
rect 180208 556288 180214 556300
rect 248506 556288 248512 556300
rect 180208 556260 248512 556288
rect 180208 556248 180214 556260
rect 248506 556248 248512 556260
rect 248564 556248 248570 556300
rect 91094 556180 91100 556232
rect 91152 556220 91158 556232
rect 122098 556220 122104 556232
rect 91152 556192 122104 556220
rect 91152 556180 91158 556192
rect 122098 556180 122104 556192
rect 122156 556180 122162 556232
rect 155310 556180 155316 556232
rect 155368 556220 155374 556232
rect 207014 556220 207020 556232
rect 155368 556192 207020 556220
rect 155368 556180 155374 556192
rect 207014 556180 207020 556192
rect 207072 556220 207078 556232
rect 582466 556220 582472 556232
rect 207072 556192 582472 556220
rect 207072 556180 207078 556192
rect 582466 556180 582472 556192
rect 582524 556180 582530 556232
rect 190362 554820 190368 554872
rect 190420 554860 190426 554872
rect 235258 554860 235264 554872
rect 190420 554832 235264 554860
rect 190420 554820 190426 554832
rect 235258 554820 235264 554832
rect 235316 554820 235322 554872
rect 43990 554752 43996 554804
rect 44048 554792 44054 554804
rect 66806 554792 66812 554804
rect 44048 554764 66812 554792
rect 44048 554752 44054 554764
rect 66806 554752 66812 554764
rect 66864 554752 66870 554804
rect 91094 554752 91100 554804
rect 91152 554792 91158 554804
rect 106182 554792 106188 554804
rect 91152 554764 106188 554792
rect 91152 554752 91158 554764
rect 106182 554752 106188 554764
rect 106240 554792 106246 554804
rect 247034 554792 247040 554804
rect 106240 554764 247040 554792
rect 106240 554752 106246 554764
rect 247034 554752 247040 554764
rect 247092 554792 247098 554804
rect 580350 554792 580356 554804
rect 247092 554764 580356 554792
rect 247092 554752 247098 554764
rect 580350 554752 580356 554764
rect 580408 554752 580414 554804
rect 57790 554004 57796 554056
rect 57848 554044 57854 554056
rect 66622 554044 66628 554056
rect 57848 554016 66628 554044
rect 57848 554004 57854 554016
rect 66622 554004 66628 554016
rect 66680 554004 66686 554056
rect 2774 553800 2780 553852
rect 2832 553840 2838 553852
rect 4798 553840 4804 553852
rect 2832 553812 4804 553840
rect 2832 553800 2838 553812
rect 4798 553800 4804 553812
rect 4856 553800 4862 553852
rect 197170 553460 197176 553512
rect 197228 553500 197234 553512
rect 287054 553500 287060 553512
rect 197228 553472 287060 553500
rect 197228 553460 197234 553472
rect 287054 553460 287060 553472
rect 287112 553460 287118 553512
rect 118510 553392 118516 553444
rect 118568 553432 118574 553444
rect 212534 553432 212540 553444
rect 118568 553404 212540 553432
rect 118568 553392 118574 553404
rect 212534 553392 212540 553404
rect 212592 553392 212598 553444
rect 91094 552100 91100 552152
rect 91152 552140 91158 552152
rect 101398 552140 101404 552152
rect 91152 552112 101404 552140
rect 91152 552100 91158 552112
rect 101398 552100 101404 552112
rect 101456 552100 101462 552152
rect 184290 552100 184296 552152
rect 184348 552140 184354 552152
rect 226978 552140 226984 552152
rect 184348 552112 226984 552140
rect 184348 552100 184354 552112
rect 226978 552100 226984 552112
rect 227036 552100 227042 552152
rect 91370 552032 91376 552084
rect 91428 552072 91434 552084
rect 108390 552072 108396 552084
rect 91428 552044 108396 552072
rect 91428 552032 91434 552044
rect 108390 552032 108396 552044
rect 108448 552032 108454 552084
rect 192478 552032 192484 552084
rect 192536 552072 192542 552084
rect 270494 552072 270500 552084
rect 192536 552044 270500 552072
rect 192536 552032 192542 552044
rect 270494 552032 270500 552044
rect 270552 552032 270558 552084
rect 198826 551284 198832 551336
rect 198884 551324 198890 551336
rect 331214 551324 331220 551336
rect 198884 551296 331220 551324
rect 198884 551284 198890 551296
rect 331214 551284 331220 551296
rect 331272 551284 331278 551336
rect 182910 550672 182916 550724
rect 182968 550712 182974 550724
rect 238754 550712 238760 550724
rect 182968 550684 238760 550712
rect 182968 550672 182974 550684
rect 238754 550672 238760 550684
rect 238812 550672 238818 550724
rect 91094 550604 91100 550656
rect 91152 550644 91158 550656
rect 124214 550644 124220 550656
rect 91152 550616 124220 550644
rect 91152 550604 91158 550616
rect 124214 550604 124220 550616
rect 124272 550644 124278 550656
rect 187142 550644 187148 550656
rect 124272 550616 187148 550644
rect 124272 550604 124278 550616
rect 187142 550604 187148 550616
rect 187200 550604 187206 550656
rect 199838 549312 199844 549364
rect 199896 549352 199902 549364
rect 251818 549352 251824 549364
rect 199896 549324 251824 549352
rect 199896 549312 199902 549324
rect 251818 549312 251824 549324
rect 251876 549312 251882 549364
rect 60642 549244 60648 549296
rect 60700 549284 60706 549296
rect 66806 549284 66812 549296
rect 60700 549256 66812 549284
rect 60700 549244 60706 549256
rect 66806 549244 66812 549256
rect 66864 549244 66870 549296
rect 91094 549244 91100 549296
rect 91152 549284 91158 549296
rect 97902 549284 97908 549296
rect 91152 549256 97908 549284
rect 91152 549244 91158 549256
rect 97902 549244 97908 549256
rect 97960 549284 97966 549296
rect 278038 549284 278044 549296
rect 97960 549256 278044 549284
rect 97960 549244 97966 549256
rect 278038 549244 278044 549256
rect 278096 549244 278102 549296
rect 90450 549176 90456 549228
rect 90508 549216 90514 549228
rect 91278 549216 91284 549228
rect 90508 549188 91284 549216
rect 90508 549176 90514 549188
rect 91278 549176 91284 549188
rect 91336 549176 91342 549228
rect 193858 547952 193864 548004
rect 193916 547992 193922 548004
rect 237374 547992 237380 548004
rect 193916 547964 237380 547992
rect 193916 547952 193922 547964
rect 237374 547952 237380 547964
rect 237432 547952 237438 548004
rect 59262 547884 59268 547936
rect 59320 547924 59326 547936
rect 66806 547924 66812 547936
rect 59320 547896 66812 547924
rect 59320 547884 59326 547896
rect 66806 547884 66812 547896
rect 66864 547884 66870 547936
rect 91278 547884 91284 547936
rect 91336 547924 91342 547936
rect 95234 547924 95240 547936
rect 91336 547896 95240 547924
rect 91336 547884 91342 547896
rect 95234 547884 95240 547896
rect 95292 547884 95298 547936
rect 177850 547884 177856 547936
rect 177908 547924 177914 547936
rect 284294 547924 284300 547936
rect 177908 547896 284300 547924
rect 177908 547884 177914 547896
rect 284294 547884 284300 547896
rect 284352 547884 284358 547936
rect 95234 547136 95240 547188
rect 95292 547176 95298 547188
rect 245654 547176 245660 547188
rect 95292 547148 245660 547176
rect 95292 547136 95298 547148
rect 245654 547136 245660 547148
rect 245712 547136 245718 547188
rect 52362 546456 52368 546508
rect 52420 546496 52426 546508
rect 66806 546496 66812 546508
rect 52420 546468 66812 546496
rect 52420 546456 52426 546468
rect 66806 546456 66812 546468
rect 66864 546456 66870 546508
rect 185578 546456 185584 546508
rect 185636 546496 185642 546508
rect 229094 546496 229100 546508
rect 185636 546468 229100 546496
rect 185636 546456 185642 546468
rect 229094 546456 229100 546468
rect 229152 546456 229158 546508
rect 324314 545572 324320 545624
rect 324372 545612 324378 545624
rect 324866 545612 324872 545624
rect 324372 545584 324872 545612
rect 324372 545572 324378 545584
rect 324866 545572 324872 545584
rect 324924 545612 324930 545624
rect 327718 545612 327724 545624
rect 324924 545584 327724 545612
rect 324924 545572 324930 545584
rect 327718 545572 327724 545584
rect 327776 545572 327782 545624
rect 188430 545164 188436 545216
rect 188488 545204 188494 545216
rect 324314 545204 324320 545216
rect 188488 545176 324320 545204
rect 188488 545164 188494 545176
rect 324314 545164 324320 545176
rect 324372 545164 324378 545216
rect 327074 545164 327080 545216
rect 327132 545204 327138 545216
rect 367094 545204 367100 545216
rect 327132 545176 367100 545204
rect 327132 545164 327138 545176
rect 367094 545164 367100 545176
rect 367152 545164 367158 545216
rect 50982 545096 50988 545148
rect 51040 545136 51046 545148
rect 66806 545136 66812 545148
rect 51040 545108 66812 545136
rect 51040 545096 51046 545108
rect 66806 545096 66812 545108
rect 66864 545096 66870 545148
rect 91554 545096 91560 545148
rect 91612 545136 91618 545148
rect 97258 545136 97264 545148
rect 91612 545108 97264 545136
rect 91612 545096 91618 545108
rect 97258 545096 97264 545108
rect 97316 545096 97322 545148
rect 137922 545096 137928 545148
rect 137980 545136 137986 545148
rect 300026 545136 300032 545148
rect 137980 545108 300032 545136
rect 137980 545096 137986 545108
rect 300026 545096 300032 545108
rect 300084 545096 300090 545148
rect 309962 545096 309968 545148
rect 310020 545136 310026 545148
rect 360286 545136 360292 545148
rect 310020 545108 360292 545136
rect 310020 545096 310026 545108
rect 360286 545096 360292 545108
rect 360344 545096 360350 545148
rect 194502 543804 194508 543856
rect 194560 543844 194566 543856
rect 223666 543844 223672 543856
rect 194560 543816 223672 543844
rect 194560 543804 194566 543816
rect 223666 543804 223672 543816
rect 223724 543804 223730 543856
rect 55030 543736 55036 543788
rect 55088 543776 55094 543788
rect 66806 543776 66812 543788
rect 55088 543748 66812 543776
rect 55088 543736 55094 543748
rect 66806 543736 66812 543748
rect 66864 543736 66870 543788
rect 89622 543736 89628 543788
rect 89680 543776 89686 543788
rect 270678 543776 270684 543788
rect 89680 543748 270684 543776
rect 89680 543736 89686 543748
rect 270678 543736 270684 543748
rect 270736 543736 270742 543788
rect 316586 543736 316592 543788
rect 316644 543776 316650 543788
rect 363046 543776 363052 543788
rect 316644 543748 363052 543776
rect 316644 543736 316650 543748
rect 363046 543736 363052 543748
rect 363104 543736 363110 543788
rect 357342 543668 357348 543720
rect 357400 543708 357406 543720
rect 582926 543708 582932 543720
rect 357400 543680 582932 543708
rect 357400 543668 357406 543680
rect 582926 543668 582932 543680
rect 582984 543668 582990 543720
rect 3418 542988 3424 543040
rect 3476 543028 3482 543040
rect 34514 543028 34520 543040
rect 3476 543000 34520 543028
rect 3476 542988 3482 543000
rect 34514 542988 34520 543000
rect 34572 542988 34578 543040
rect 195330 542444 195336 542496
rect 195388 542484 195394 542496
rect 218698 542484 218704 542496
rect 195388 542456 218704 542484
rect 195388 542444 195394 542456
rect 218698 542444 218704 542456
rect 218756 542444 218762 542496
rect 255958 542444 255964 542496
rect 256016 542484 256022 542496
rect 257338 542484 257344 542496
rect 256016 542456 257344 542484
rect 256016 542444 256022 542456
rect 257338 542444 257344 542456
rect 257396 542484 257402 542496
rect 356054 542484 356060 542496
rect 257396 542456 356060 542484
rect 257396 542444 257402 542456
rect 356054 542444 356060 542456
rect 356112 542484 356118 542496
rect 357342 542484 357348 542496
rect 356112 542456 357348 542484
rect 356112 542444 356118 542456
rect 357342 542444 357348 542456
rect 357400 542444 357406 542496
rect 34514 542376 34520 542428
rect 34572 542416 34578 542428
rect 35802 542416 35808 542428
rect 34572 542388 35808 542416
rect 34572 542376 34578 542388
rect 35802 542376 35808 542388
rect 35860 542416 35866 542428
rect 66806 542416 66812 542428
rect 35860 542388 66812 542416
rect 35860 542376 35866 542388
rect 66806 542376 66812 542388
rect 66864 542376 66870 542428
rect 91554 542376 91560 542428
rect 91612 542416 91618 542428
rect 95970 542416 95976 542428
rect 91612 542388 95976 542416
rect 91612 542376 91618 542388
rect 95970 542376 95976 542388
rect 96028 542376 96034 542428
rect 129642 542376 129648 542428
rect 129700 542416 129706 542428
rect 266722 542416 266728 542428
rect 129700 542388 266728 542416
rect 129700 542376 129706 542388
rect 266722 542376 266728 542388
rect 266780 542376 266786 542428
rect 67358 541832 67364 541884
rect 67416 541872 67422 541884
rect 67542 541872 67548 541884
rect 67416 541844 67548 541872
rect 67416 541832 67422 541844
rect 67542 541832 67548 541844
rect 67600 541832 67606 541884
rect 14458 541628 14464 541680
rect 14516 541668 14522 541680
rect 66990 541668 66996 541680
rect 14516 541640 66996 541668
rect 14516 541628 14522 541640
rect 66990 541628 66996 541640
rect 67048 541668 67054 541680
rect 67266 541668 67272 541680
rect 67048 541640 67272 541668
rect 67048 541628 67054 541640
rect 67266 541628 67272 541640
rect 67324 541628 67330 541680
rect 261754 541628 261760 541680
rect 261812 541668 261818 541680
rect 360194 541668 360200 541680
rect 261812 541640 360200 541668
rect 261812 541628 261818 541640
rect 360194 541628 360200 541640
rect 360252 541628 360258 541680
rect 189718 541016 189724 541068
rect 189776 541056 189782 541068
rect 230474 541056 230480 541068
rect 189776 541028 230480 541056
rect 189776 541016 189782 541028
rect 230474 541016 230480 541028
rect 230532 541016 230538 541068
rect 91922 540948 91928 541000
rect 91980 540988 91986 541000
rect 92382 540988 92388 541000
rect 91980 540960 92388 540988
rect 91980 540948 91986 540960
rect 92382 540948 92388 540960
rect 92440 540988 92446 541000
rect 124858 540988 124864 541000
rect 92440 540960 124864 540988
rect 92440 540948 92446 540960
rect 124858 540948 124864 540960
rect 124916 540988 124922 541000
rect 258442 540988 258448 541000
rect 124916 540960 258448 540988
rect 124916 540948 124922 540960
rect 258442 540948 258448 540960
rect 258500 540948 258506 541000
rect 338298 540948 338304 541000
rect 338356 540988 338362 541000
rect 367370 540988 367376 541000
rect 338356 540960 367376 540988
rect 338356 540948 338362 540960
rect 367370 540948 367376 540960
rect 367428 540948 367434 541000
rect 4798 540200 4804 540252
rect 4856 540240 4862 540252
rect 4856 540212 64874 540240
rect 4856 540200 4862 540212
rect 64846 539764 64874 540212
rect 64846 539736 69980 539764
rect 65886 539656 65892 539708
rect 65944 539696 65950 539708
rect 65944 539668 69888 539696
rect 65944 539656 65950 539668
rect 69860 539572 69888 539668
rect 69952 539628 69980 539736
rect 84166 539736 93854 539764
rect 70394 539628 70400 539640
rect 69952 539600 70400 539628
rect 70394 539588 70400 539600
rect 70452 539588 70458 539640
rect 81342 539588 81348 539640
rect 81400 539628 81406 539640
rect 84166 539628 84194 539736
rect 88794 539696 88800 539708
rect 81400 539600 84194 539628
rect 85592 539668 88800 539696
rect 81400 539588 81406 539600
rect 85592 539572 85620 539668
rect 88794 539656 88800 539668
rect 88852 539656 88858 539708
rect 93826 539628 93854 539736
rect 195146 539656 195152 539708
rect 195204 539696 195210 539708
rect 215846 539696 215852 539708
rect 195204 539668 215852 539696
rect 195204 539656 195210 539668
rect 215846 539656 215852 539668
rect 215904 539656 215910 539708
rect 315390 539656 315396 539708
rect 315448 539696 315454 539708
rect 361574 539696 361580 539708
rect 315448 539668 361580 539696
rect 315448 539656 315454 539668
rect 361574 539656 361580 539668
rect 361632 539656 361638 539708
rect 250622 539628 250628 539640
rect 93826 539600 250628 539628
rect 250622 539588 250628 539600
rect 250680 539588 250686 539640
rect 323578 539588 323584 539640
rect 323636 539628 323642 539640
rect 379422 539628 379428 539640
rect 323636 539600 379428 539628
rect 323636 539588 323642 539600
rect 379422 539588 379428 539600
rect 379480 539588 379486 539640
rect 69842 539520 69848 539572
rect 69900 539520 69906 539572
rect 85574 539520 85580 539572
rect 85632 539520 85638 539572
rect 268378 539520 268384 539572
rect 268436 539560 268442 539572
rect 272334 539560 272340 539572
rect 268436 539532 272340 539560
rect 268436 539520 268442 539532
rect 272334 539520 272340 539532
rect 272392 539520 272398 539572
rect 273254 539520 273260 539572
rect 273312 539560 273318 539572
rect 275646 539560 275652 539572
rect 273312 539532 275652 539560
rect 273312 539520 273318 539532
rect 275646 539520 275652 539532
rect 275704 539520 275710 539572
rect 278038 539520 278044 539572
rect 278096 539560 278102 539572
rect 278958 539560 278964 539572
rect 278096 539532 278964 539560
rect 278096 539520 278102 539532
rect 278958 539520 278964 539532
rect 279016 539520 279022 539572
rect 341518 539520 341524 539572
rect 341576 539560 341582 539572
rect 343726 539560 343732 539572
rect 341576 539532 343732 539560
rect 341576 539520 341582 539532
rect 343726 539520 343732 539532
rect 343784 539520 343790 539572
rect 345382 539520 345388 539572
rect 345440 539560 345446 539572
rect 349982 539560 349988 539572
rect 345440 539532 349988 539560
rect 345440 539520 345446 539532
rect 349982 539520 349988 539532
rect 350040 539520 350046 539572
rect 66162 538976 66168 539028
rect 66220 539016 66226 539028
rect 72418 539016 72424 539028
rect 66220 538988 72424 539016
rect 66220 538976 66226 538988
rect 72418 538976 72424 538988
rect 72476 538976 72482 539028
rect 72436 538948 72464 538976
rect 76742 538948 76748 538960
rect 72436 538920 76748 538948
rect 76742 538908 76748 538920
rect 76800 538908 76806 538960
rect 171778 538908 171784 538960
rect 171836 538948 171842 538960
rect 195146 538948 195152 538960
rect 171836 538920 195152 538948
rect 171836 538908 171842 538920
rect 195146 538908 195152 538920
rect 195204 538908 195210 538960
rect 7558 538840 7564 538892
rect 7616 538880 7622 538892
rect 91094 538880 91100 538892
rect 7616 538852 91100 538880
rect 7616 538840 7622 538852
rect 91094 538840 91100 538852
rect 91152 538840 91158 538892
rect 169018 538840 169024 538892
rect 169076 538880 169082 538892
rect 195238 538880 195244 538892
rect 169076 538852 195244 538880
rect 169076 538840 169082 538852
rect 195238 538840 195244 538852
rect 195296 538840 195302 538892
rect 195238 538296 195244 538348
rect 195296 538336 195302 538348
rect 223206 538336 223212 538348
rect 195296 538308 223212 538336
rect 195296 538296 195302 538308
rect 223206 538296 223212 538308
rect 223264 538296 223270 538348
rect 347038 538296 347044 538348
rect 347096 538336 347102 538348
rect 358814 538336 358820 538348
rect 347096 538308 358820 538336
rect 347096 538296 347102 538308
rect 358814 538296 358820 538308
rect 358872 538296 358878 538348
rect 226242 538228 226248 538280
rect 226300 538268 226306 538280
rect 297174 538268 297180 538280
rect 226300 538240 297180 538268
rect 226300 538228 226306 538240
rect 297174 538228 297180 538240
rect 297232 538228 297238 538280
rect 350350 538228 350356 538280
rect 350408 538268 350414 538280
rect 369854 538268 369860 538280
rect 350408 538240 369860 538268
rect 350408 538228 350414 538240
rect 369854 538228 369860 538240
rect 369912 538228 369918 538280
rect 88610 538160 88616 538212
rect 88668 538200 88674 538212
rect 89622 538200 89628 538212
rect 88668 538172 89628 538200
rect 88668 538160 88674 538172
rect 89622 538160 89628 538172
rect 89680 538160 89686 538212
rect 379422 538160 379428 538212
rect 379480 538200 379486 538212
rect 580166 538200 580172 538212
rect 379480 538172 580172 538200
rect 379480 538160 379486 538172
rect 580166 538160 580172 538172
rect 580224 538160 580230 538212
rect 12342 537548 12348 537600
rect 12400 537588 12406 537600
rect 91186 537588 91192 537600
rect 12400 537560 91192 537588
rect 12400 537548 12406 537560
rect 91186 537548 91192 537560
rect 91244 537548 91250 537600
rect 67542 537480 67548 537532
rect 67600 537520 67606 537532
rect 154758 537520 154764 537532
rect 67600 537492 154764 537520
rect 67600 537480 67606 537492
rect 154758 537480 154764 537492
rect 154816 537480 154822 537532
rect 197538 536868 197544 536920
rect 197596 536908 197602 536920
rect 220814 536908 220820 536920
rect 197596 536880 220820 536908
rect 197596 536868 197602 536880
rect 220814 536868 220820 536880
rect 220872 536868 220878 536920
rect 330478 536868 330484 536920
rect 330536 536908 330542 536920
rect 364426 536908 364432 536920
rect 330536 536880 364432 536908
rect 330536 536868 330542 536880
rect 364426 536868 364432 536880
rect 364484 536868 364490 536920
rect 178770 536800 178776 536852
rect 178828 536840 178834 536852
rect 233878 536840 233884 536852
rect 178828 536812 233884 536840
rect 178828 536800 178834 536812
rect 233878 536800 233884 536812
rect 233936 536840 233942 536852
rect 234062 536840 234068 536852
rect 233936 536812 234068 536840
rect 233936 536800 233942 536812
rect 234062 536800 234068 536812
rect 234120 536800 234126 536852
rect 342070 536800 342076 536852
rect 342128 536840 342134 536852
rect 378134 536840 378140 536852
rect 342128 536812 378140 536840
rect 342128 536800 342134 536812
rect 378134 536800 378140 536812
rect 378192 536800 378198 536852
rect 43438 536732 43444 536784
rect 43496 536772 43502 536784
rect 69566 536772 69572 536784
rect 43496 536744 69572 536772
rect 43496 536732 43502 536744
rect 69566 536732 69572 536744
rect 69624 536732 69630 536784
rect 86862 536732 86868 536784
rect 86920 536772 86926 536784
rect 130378 536772 130384 536784
rect 86920 536744 130384 536772
rect 86920 536732 86926 536744
rect 130378 536732 130384 536744
rect 130436 536732 130442 536784
rect 68646 536664 68652 536716
rect 68704 536704 68710 536716
rect 81342 536704 81348 536716
rect 68704 536676 81348 536704
rect 68704 536664 68710 536676
rect 81342 536664 81348 536676
rect 81400 536664 81406 536716
rect 75178 536596 75184 536648
rect 75236 536636 75242 536648
rect 85574 536636 85580 536648
rect 75236 536608 85580 536636
rect 75236 536596 75242 536608
rect 85574 536596 85580 536608
rect 85632 536596 85638 536648
rect 84286 536460 84292 536512
rect 84344 536500 84350 536512
rect 89070 536500 89076 536512
rect 84344 536472 89076 536500
rect 84344 536460 84350 536472
rect 89070 536460 89076 536472
rect 89128 536460 89134 536512
rect 81526 535576 81532 535628
rect 81584 535616 81590 535628
rect 83458 535616 83464 535628
rect 81584 535588 83464 535616
rect 81584 535576 81590 535588
rect 83458 535576 83464 535588
rect 83516 535576 83522 535628
rect 170490 535508 170496 535560
rect 170548 535548 170554 535560
rect 313366 535548 313372 535560
rect 170548 535520 313372 535548
rect 170548 535508 170554 535520
rect 313366 535508 313372 535520
rect 313424 535508 313430 535560
rect 332410 535508 332416 535560
rect 332468 535548 332474 535560
rect 358906 535548 358912 535560
rect 332468 535520 358912 535548
rect 332468 535508 332474 535520
rect 358906 535508 358912 535520
rect 358964 535508 358970 535560
rect 89622 535440 89628 535492
rect 89680 535480 89686 535492
rect 90542 535480 90548 535492
rect 89680 535452 90548 535480
rect 89680 535440 89686 535452
rect 90542 535440 90548 535452
rect 90600 535440 90606 535492
rect 146938 535440 146944 535492
rect 146996 535480 147002 535492
rect 293494 535480 293500 535492
rect 146996 535452 293500 535480
rect 146996 535440 147002 535452
rect 293494 535440 293500 535452
rect 293552 535440 293558 535492
rect 302326 535440 302332 535492
rect 302384 535480 302390 535492
rect 582742 535480 582748 535492
rect 302384 535452 582748 535480
rect 302384 535440 302390 535452
rect 582742 535440 582748 535452
rect 582800 535440 582806 535492
rect 199654 535372 199660 535424
rect 199712 535412 199718 535424
rect 202046 535412 202052 535424
rect 199712 535384 202052 535412
rect 199712 535372 199718 535384
rect 202046 535372 202052 535384
rect 202104 535372 202110 535424
rect 226242 535276 226248 535288
rect 219406 535248 226248 535276
rect 196618 534760 196624 534812
rect 196676 534800 196682 534812
rect 219406 534800 219434 535248
rect 226242 535236 226248 535248
rect 226300 535236 226306 535288
rect 355594 535236 355600 535288
rect 355652 535276 355658 535288
rect 355652 535248 364334 535276
rect 355652 535236 355658 535248
rect 196676 534772 219434 534800
rect 364306 534800 364334 535248
rect 425054 534800 425060 534812
rect 364306 534772 425060 534800
rect 196676 534760 196682 534772
rect 425054 534760 425060 534772
rect 425112 534760 425118 534812
rect 78306 534692 78312 534744
rect 78364 534732 78370 534744
rect 135254 534732 135260 534744
rect 78364 534704 135260 534732
rect 78364 534692 78370 534704
rect 135254 534692 135260 534704
rect 135312 534732 135318 534744
rect 136174 534732 136180 534744
rect 135312 534704 136180 534732
rect 135312 534692 135318 534704
rect 136174 534692 136180 534704
rect 136232 534692 136238 534744
rect 151078 534692 151084 534744
rect 151136 534732 151142 534744
rect 198734 534732 198740 534744
rect 151136 534704 198740 534732
rect 151136 534692 151142 534704
rect 198734 534692 198740 534704
rect 198792 534692 198798 534744
rect 136174 534080 136180 534132
rect 136232 534120 136238 534132
rect 143442 534120 143448 534132
rect 136232 534092 143448 534120
rect 136232 534080 136238 534092
rect 143442 534080 143448 534092
rect 143500 534080 143506 534132
rect 41322 534012 41328 534064
rect 41380 534052 41386 534064
rect 191098 534052 191104 534064
rect 41380 534024 191104 534052
rect 41380 534012 41386 534024
rect 191098 534012 191104 534024
rect 191156 534012 191162 534064
rect 78674 533332 78680 533384
rect 78732 533372 78738 533384
rect 79502 533372 79508 533384
rect 78732 533344 79508 533372
rect 78732 533332 78738 533344
rect 79502 533332 79508 533344
rect 79560 533332 79566 533384
rect 143442 532652 143448 532704
rect 143500 532692 143506 532704
rect 197446 532692 197452 532704
rect 143500 532664 197452 532692
rect 143500 532652 143506 532664
rect 197446 532652 197452 532664
rect 197504 532652 197510 532704
rect 81066 532040 81072 532092
rect 81124 532080 81130 532092
rect 132494 532080 132500 532092
rect 81124 532052 132500 532080
rect 81124 532040 81130 532052
rect 132494 532040 132500 532052
rect 132552 532080 132558 532092
rect 133690 532080 133696 532092
rect 132552 532052 133696 532080
rect 132552 532040 132558 532052
rect 133690 532040 133696 532052
rect 133748 532040 133754 532092
rect 3418 531972 3424 532024
rect 3476 532012 3482 532024
rect 89714 532012 89720 532024
rect 3476 531984 89720 532012
rect 3476 531972 3482 531984
rect 89714 531972 89720 531984
rect 89772 531972 89778 532024
rect 358722 531972 358728 532024
rect 358780 532012 358786 532024
rect 358998 532012 359004 532024
rect 358780 531984 359004 532012
rect 358780 531972 358786 531984
rect 358998 531972 359004 531984
rect 359056 532012 359062 532024
rect 582926 532012 582932 532024
rect 359056 531984 582932 532012
rect 359056 531972 359062 531984
rect 582926 531972 582932 531984
rect 582984 531972 582990 532024
rect 133690 531292 133696 531344
rect 133748 531332 133754 531344
rect 144178 531332 144184 531344
rect 133748 531304 144184 531332
rect 133748 531292 133754 531304
rect 144178 531292 144184 531304
rect 144236 531292 144242 531344
rect 79318 531224 79324 531276
rect 79376 531264 79382 531276
rect 79962 531264 79968 531276
rect 79376 531236 79968 531264
rect 79376 531224 79382 531236
rect 79962 531224 79968 531236
rect 80020 531224 80026 531276
rect 180058 530612 180064 530664
rect 180116 530652 180122 530664
rect 197538 530652 197544 530664
rect 180116 530624 197544 530652
rect 180116 530612 180122 530624
rect 197538 530612 197544 530624
rect 197596 530612 197602 530664
rect 64690 530544 64696 530596
rect 64748 530584 64754 530596
rect 79318 530584 79324 530596
rect 64748 530556 79324 530584
rect 64748 530544 64754 530556
rect 79318 530544 79324 530556
rect 79376 530544 79382 530596
rect 153102 530544 153108 530596
rect 153160 530584 153166 530596
rect 199654 530584 199660 530596
rect 153160 530556 199660 530584
rect 153160 530544 153166 530556
rect 199654 530544 199660 530556
rect 199712 530544 199718 530596
rect 50982 529864 50988 529916
rect 51040 529904 51046 529916
rect 178678 529904 178684 529916
rect 51040 529876 178684 529904
rect 51040 529864 51046 529876
rect 178678 529864 178684 529876
rect 178736 529864 178742 529916
rect 154758 529796 154764 529848
rect 154816 529836 154822 529848
rect 197446 529836 197452 529848
rect 154816 529808 197452 529836
rect 154816 529796 154822 529808
rect 197446 529796 197452 529808
rect 197504 529796 197510 529848
rect 358722 528572 358728 528624
rect 358780 528612 358786 528624
rect 367278 528612 367284 528624
rect 358780 528584 367284 528612
rect 358780 528572 358786 528584
rect 367278 528572 367284 528584
rect 367336 528572 367342 528624
rect 187142 528504 187148 528556
rect 187200 528544 187206 528556
rect 197446 528544 197452 528556
rect 187200 528516 197452 528544
rect 187200 528504 187206 528516
rect 197446 528504 197452 528516
rect 197504 528504 197510 528556
rect 358722 527144 358728 527196
rect 358780 527184 358786 527196
rect 398834 527184 398840 527196
rect 358780 527156 398840 527184
rect 358780 527144 358786 527156
rect 398834 527144 398840 527156
rect 398892 527144 398898 527196
rect 70486 526532 70492 526584
rect 70544 526572 70550 526584
rect 71038 526572 71044 526584
rect 70544 526544 71044 526572
rect 70544 526532 70550 526544
rect 71038 526532 71044 526544
rect 71096 526532 71102 526584
rect 71038 525784 71044 525836
rect 71096 525824 71102 525836
rect 162210 525824 162216 525836
rect 71096 525796 162216 525824
rect 71096 525784 71102 525796
rect 162210 525784 162216 525796
rect 162268 525784 162274 525836
rect 61930 525104 61936 525156
rect 61988 525144 61994 525156
rect 77938 525144 77944 525156
rect 61988 525116 77944 525144
rect 61988 525104 61994 525116
rect 77938 525104 77944 525116
rect 77996 525104 78002 525156
rect 50890 525036 50896 525088
rect 50948 525076 50954 525088
rect 191098 525076 191104 525088
rect 50948 525048 191104 525076
rect 50948 525036 50954 525048
rect 191098 525036 191104 525048
rect 191156 525036 191162 525088
rect 358722 524424 358728 524476
rect 358780 524464 358786 524476
rect 371234 524464 371240 524476
rect 358780 524436 371240 524464
rect 358780 524424 358786 524436
rect 371234 524424 371240 524436
rect 371292 524424 371298 524476
rect 34422 523676 34428 523728
rect 34480 523716 34486 523728
rect 195330 523716 195336 523728
rect 34480 523688 195336 523716
rect 34480 523676 34486 523688
rect 195330 523676 195336 523688
rect 195388 523676 195394 523728
rect 60642 522928 60648 522980
rect 60700 522968 60706 522980
rect 185670 522968 185676 522980
rect 60700 522940 185676 522968
rect 60700 522928 60706 522940
rect 185670 522928 185676 522940
rect 185728 522928 185734 522980
rect 155218 521636 155224 521688
rect 155276 521676 155282 521688
rect 197446 521676 197452 521688
rect 155276 521648 197452 521676
rect 155276 521636 155282 521648
rect 197446 521636 197452 521648
rect 197504 521636 197510 521688
rect 167638 520956 167644 521008
rect 167696 520996 167702 521008
rect 197538 520996 197544 521008
rect 167696 520968 197544 520996
rect 167696 520956 167702 520968
rect 197538 520956 197544 520968
rect 197596 520956 197602 521008
rect 63402 520888 63408 520940
rect 63460 520928 63466 520940
rect 187050 520928 187056 520940
rect 63460 520900 187056 520928
rect 63460 520888 63466 520900
rect 187050 520888 187056 520900
rect 187108 520888 187114 520940
rect 358722 520888 358728 520940
rect 358780 520928 358786 520940
rect 395982 520928 395988 520940
rect 358780 520900 395988 520928
rect 358780 520888 358786 520900
rect 395982 520888 395988 520900
rect 396040 520888 396046 520940
rect 395982 520276 395988 520328
rect 396040 520316 396046 520328
rect 582374 520316 582380 520328
rect 396040 520288 582380 520316
rect 396040 520276 396046 520288
rect 582374 520276 582380 520288
rect 582432 520276 582438 520328
rect 53742 519528 53748 519580
rect 53800 519568 53806 519580
rect 196710 519568 196716 519580
rect 53800 519540 196716 519568
rect 53800 519528 53806 519540
rect 196710 519528 196716 519540
rect 196768 519528 196774 519580
rect 358630 518916 358636 518968
rect 358688 518956 358694 518968
rect 445754 518956 445760 518968
rect 358688 518928 445760 518956
rect 358688 518916 358694 518928
rect 445754 518916 445760 518928
rect 445812 518916 445818 518968
rect 52362 518848 52368 518900
rect 52420 518888 52426 518900
rect 188430 518888 188436 518900
rect 52420 518860 188436 518888
rect 52420 518848 52426 518860
rect 188430 518848 188436 518860
rect 188488 518848 188494 518900
rect 52178 517488 52184 517540
rect 52236 517528 52242 517540
rect 52362 517528 52368 517540
rect 52236 517500 52368 517528
rect 52236 517488 52242 517500
rect 52362 517488 52368 517500
rect 52420 517488 52426 517540
rect 162118 516128 162124 516180
rect 162176 516168 162182 516180
rect 197446 516168 197452 516180
rect 162176 516140 197452 516168
rect 162176 516128 162182 516140
rect 197446 516128 197452 516140
rect 197504 516128 197510 516180
rect 358722 516128 358728 516180
rect 358780 516168 358786 516180
rect 363598 516168 363604 516180
rect 358780 516140 363604 516168
rect 358780 516128 358786 516140
rect 363598 516128 363604 516140
rect 363656 516128 363662 516180
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 14458 514808 14464 514820
rect 3568 514780 14464 514808
rect 3568 514768 3574 514780
rect 14458 514768 14464 514780
rect 14516 514768 14522 514820
rect 162210 510552 162216 510604
rect 162268 510592 162274 510604
rect 197446 510592 197452 510604
rect 162268 510564 197452 510592
rect 162268 510552 162274 510564
rect 197446 510552 197452 510564
rect 197504 510552 197510 510604
rect 49602 508512 49608 508564
rect 49660 508552 49666 508564
rect 189718 508552 189724 508564
rect 49660 508524 189724 508552
rect 49660 508512 49666 508524
rect 189718 508512 189724 508524
rect 189776 508512 189782 508564
rect 134518 507084 134524 507136
rect 134576 507124 134582 507136
rect 193950 507124 193956 507136
rect 134576 507096 193956 507124
rect 134576 507084 134582 507096
rect 193950 507084 193956 507096
rect 194008 507084 194014 507136
rect 358722 506472 358728 506524
rect 358780 506512 358786 506524
rect 382274 506512 382280 506524
rect 358780 506484 382280 506512
rect 358780 506472 358786 506484
rect 382274 506472 382280 506484
rect 382332 506472 382338 506524
rect 358722 505112 358728 505164
rect 358780 505152 358786 505164
rect 434714 505152 434720 505164
rect 358780 505124 434720 505152
rect 358780 505112 358786 505124
rect 434714 505112 434720 505124
rect 434772 505112 434778 505164
rect 61930 504364 61936 504416
rect 61988 504404 61994 504416
rect 180150 504404 180156 504416
rect 61988 504376 180156 504404
rect 61988 504364 61994 504376
rect 180150 504364 180156 504376
rect 180208 504364 180214 504416
rect 173158 502936 173164 502988
rect 173216 502976 173222 502988
rect 197446 502976 197452 502988
rect 173216 502948 197452 502976
rect 173216 502936 173222 502948
rect 197446 502936 197452 502948
rect 197504 502936 197510 502988
rect 358722 502392 358728 502444
rect 358780 502432 358786 502444
rect 364334 502432 364340 502444
rect 358780 502404 364340 502432
rect 358780 502392 358786 502404
rect 364334 502392 364340 502404
rect 364392 502392 364398 502444
rect 187142 502324 187148 502376
rect 187200 502364 187206 502376
rect 197446 502364 197452 502376
rect 187200 502336 197452 502364
rect 187200 502324 187206 502336
rect 197446 502324 197452 502336
rect 197504 502324 197510 502376
rect 2774 501848 2780 501900
rect 2832 501888 2838 501900
rect 4798 501888 4804 501900
rect 2832 501860 4804 501888
rect 2832 501848 2838 501860
rect 4798 501848 4804 501860
rect 4856 501848 4862 501900
rect 144178 500896 144184 500948
rect 144236 500936 144242 500948
rect 197446 500936 197452 500948
rect 144236 500908 197452 500936
rect 144236 500896 144242 500908
rect 197446 500896 197452 500908
rect 197504 500896 197510 500948
rect 363598 497428 363604 497480
rect 363656 497468 363662 497480
rect 405734 497468 405740 497480
rect 363656 497440 405740 497468
rect 363656 497428 363662 497440
rect 405734 497428 405740 497440
rect 405792 497428 405798 497480
rect 358630 496748 358636 496800
rect 358688 496788 358694 496800
rect 360194 496788 360200 496800
rect 358688 496760 360200 496788
rect 358688 496748 358694 496760
rect 360194 496748 360200 496760
rect 360252 496788 360258 496800
rect 583018 496788 583024 496800
rect 360252 496760 583024 496788
rect 360252 496748 360258 496760
rect 583018 496748 583024 496760
rect 583076 496748 583082 496800
rect 178678 495456 178684 495508
rect 178736 495496 178742 495508
rect 197446 495496 197452 495508
rect 178736 495468 197452 495496
rect 178736 495456 178742 495468
rect 197446 495456 197452 495468
rect 197504 495456 197510 495508
rect 358722 494708 358728 494760
rect 358780 494748 358786 494760
rect 385034 494748 385040 494760
rect 358780 494720 385040 494748
rect 358780 494708 358786 494720
rect 385034 494708 385040 494720
rect 385092 494708 385098 494760
rect 398926 494708 398932 494760
rect 398984 494748 398990 494760
rect 412634 494748 412640 494760
rect 398984 494720 412640 494748
rect 398984 494708 398990 494720
rect 412634 494708 412640 494720
rect 412692 494708 412698 494760
rect 392210 493280 392216 493332
rect 392268 493320 392274 493332
rect 398926 493320 398932 493332
rect 392268 493292 398932 493320
rect 392268 493280 392274 493292
rect 398926 493280 398932 493292
rect 398984 493280 398990 493332
rect 148318 492668 148324 492720
rect 148376 492708 148382 492720
rect 197446 492708 197452 492720
rect 148376 492680 197452 492708
rect 148376 492668 148382 492680
rect 197446 492668 197452 492680
rect 197504 492668 197510 492720
rect 358722 492668 358728 492720
rect 358780 492708 358786 492720
rect 392210 492708 392216 492720
rect 358780 492680 392216 492708
rect 358780 492668 358786 492680
rect 392210 492668 392216 492680
rect 392268 492708 392274 492720
rect 392578 492708 392584 492720
rect 392268 492680 392584 492708
rect 392268 492668 392274 492680
rect 392578 492668 392584 492680
rect 392636 492668 392642 492720
rect 187050 489880 187056 489932
rect 187108 489920 187114 489932
rect 197446 489920 197452 489932
rect 187108 489892 197452 489920
rect 187108 489880 187114 489892
rect 197446 489880 197452 489892
rect 197504 489880 197510 489932
rect 148410 487772 148416 487824
rect 148468 487812 148474 487824
rect 185394 487812 185400 487824
rect 148468 487784 185400 487812
rect 148468 487772 148474 487784
rect 185394 487772 185400 487784
rect 185452 487772 185458 487824
rect 184934 487160 184940 487212
rect 184992 487200 184998 487212
rect 185394 487200 185400 487212
rect 184992 487172 185400 487200
rect 184992 487160 184998 487172
rect 185394 487160 185400 487172
rect 185452 487200 185458 487212
rect 197446 487200 197452 487212
rect 185452 487172 197452 487200
rect 185452 487160 185458 487172
rect 197446 487160 197452 487172
rect 197504 487160 197510 487212
rect 358722 487160 358728 487212
rect 358780 487200 358786 487212
rect 380894 487200 380900 487212
rect 358780 487172 380900 487200
rect 358780 487160 358786 487172
rect 380894 487160 380900 487172
rect 380952 487160 380958 487212
rect 358170 484372 358176 484424
rect 358228 484412 358234 484424
rect 410518 484412 410524 484424
rect 358228 484384 410524 484412
rect 358228 484372 358234 484384
rect 410518 484372 410524 484384
rect 410576 484372 410582 484424
rect 180150 483624 180156 483676
rect 180208 483664 180214 483676
rect 197446 483664 197452 483676
rect 180208 483636 197452 483664
rect 180208 483624 180214 483636
rect 197446 483624 197452 483636
rect 197504 483624 197510 483676
rect 357894 481652 357900 481704
rect 357952 481692 357958 481704
rect 367186 481692 367192 481704
rect 357952 481664 367192 481692
rect 357952 481652 357958 481664
rect 367186 481652 367192 481664
rect 367244 481652 367250 481704
rect 132402 480224 132408 480276
rect 132460 480264 132466 480276
rect 197446 480264 197452 480276
rect 132460 480236 197452 480264
rect 132460 480224 132466 480236
rect 197446 480224 197452 480236
rect 197504 480224 197510 480276
rect 127618 477504 127624 477556
rect 127676 477544 127682 477556
rect 182082 477544 182088 477556
rect 127676 477516 182088 477544
rect 127676 477504 127682 477516
rect 182082 477504 182088 477516
rect 182140 477544 182146 477556
rect 197446 477544 197452 477556
rect 182140 477516 197452 477544
rect 182140 477504 182146 477516
rect 197446 477504 197452 477516
rect 197504 477504 197510 477556
rect 357894 477504 357900 477556
rect 357952 477544 357958 477556
rect 365714 477544 365720 477556
rect 357952 477516 365720 477544
rect 357952 477504 357958 477516
rect 365714 477504 365720 477516
rect 365772 477504 365778 477556
rect 145558 474716 145564 474768
rect 145616 474756 145622 474768
rect 197446 474756 197452 474768
rect 145616 474728 197452 474756
rect 145616 474716 145622 474728
rect 197446 474716 197452 474728
rect 197504 474716 197510 474768
rect 358722 474716 358728 474768
rect 358780 474756 358786 474768
rect 368566 474756 368572 474768
rect 358780 474728 368572 474756
rect 358780 474716 358786 474728
rect 368566 474716 368572 474728
rect 368624 474716 368630 474768
rect 3510 473968 3516 474020
rect 3568 474008 3574 474020
rect 7558 474008 7564 474020
rect 3568 473980 7564 474008
rect 3568 473968 3574 473980
rect 7558 473968 7564 473980
rect 7616 474008 7622 474020
rect 15838 474008 15844 474020
rect 7616 473980 15844 474008
rect 7616 473968 7622 473980
rect 15838 473968 15844 473980
rect 15896 473968 15902 474020
rect 142798 473356 142804 473408
rect 142856 473396 142862 473408
rect 197446 473396 197452 473408
rect 142856 473368 197452 473396
rect 142856 473356 142862 473368
rect 197446 473356 197452 473368
rect 197504 473356 197510 473408
rect 358078 473288 358084 473340
rect 358136 473328 358142 473340
rect 360194 473328 360200 473340
rect 358136 473300 360200 473328
rect 358136 473288 358142 473300
rect 360194 473288 360200 473300
rect 360252 473288 360258 473340
rect 358722 471996 358728 472048
rect 358780 472036 358786 472048
rect 374086 472036 374092 472048
rect 358780 472008 374092 472036
rect 358780 471996 358786 472008
rect 374086 471996 374092 472008
rect 374144 471996 374150 472048
rect 358722 470568 358728 470620
rect 358780 470608 358786 470620
rect 371418 470608 371424 470620
rect 358780 470580 371424 470608
rect 358780 470568 358786 470580
rect 371418 470568 371424 470580
rect 371476 470568 371482 470620
rect 59078 468460 59084 468512
rect 59136 468500 59142 468512
rect 85574 468500 85580 468512
rect 59136 468472 85580 468500
rect 59136 468460 59142 468472
rect 85574 468460 85580 468472
rect 85632 468460 85638 468512
rect 165522 467848 165528 467900
rect 165580 467888 165586 467900
rect 197446 467888 197452 467900
rect 165580 467860 197452 467888
rect 165580 467848 165586 467860
rect 197446 467848 197452 467860
rect 197504 467848 197510 467900
rect 67818 467780 67824 467832
rect 67876 467820 67882 467832
rect 74534 467820 74540 467832
rect 67876 467792 74540 467820
rect 67876 467780 67882 467792
rect 74534 467780 74540 467792
rect 74592 467780 74598 467832
rect 156598 465672 156604 465724
rect 156656 465712 156662 465724
rect 197446 465712 197452 465724
rect 156656 465684 197452 465712
rect 156656 465672 156662 465684
rect 197446 465672 197452 465684
rect 197504 465672 197510 465724
rect 130562 465060 130568 465112
rect 130620 465100 130626 465112
rect 156598 465100 156604 465112
rect 130620 465072 156604 465100
rect 130620 465060 130626 465072
rect 156598 465060 156604 465072
rect 156656 465060 156662 465112
rect 358722 465060 358728 465112
rect 358780 465100 358786 465112
rect 379514 465100 379520 465112
rect 358780 465072 379520 465100
rect 358780 465060 358786 465072
rect 379514 465060 379520 465072
rect 379572 465100 379578 465112
rect 583294 465100 583300 465112
rect 379572 465072 583300 465100
rect 379572 465060 379578 465072
rect 583294 465060 583300 465072
rect 583352 465060 583358 465112
rect 106182 464312 106188 464364
rect 106240 464352 106246 464364
rect 120810 464352 120816 464364
rect 106240 464324 120816 464352
rect 106240 464312 106246 464324
rect 120810 464312 120816 464324
rect 120868 464312 120874 464364
rect 65978 462952 65984 463004
rect 66036 462992 66042 463004
rect 91554 462992 91560 463004
rect 66036 462964 91560 462992
rect 66036 462952 66042 462964
rect 91554 462952 91560 462964
rect 91612 462952 91618 463004
rect 107010 462952 107016 463004
rect 107068 462992 107074 463004
rect 122926 462992 122932 463004
rect 107068 462964 122932 462992
rect 107068 462952 107074 462964
rect 122926 462952 122932 462964
rect 122984 462952 122990 463004
rect 2774 462544 2780 462596
rect 2832 462584 2838 462596
rect 4798 462584 4804 462596
rect 2832 462556 4804 462584
rect 2832 462544 2838 462556
rect 4798 462544 4804 462556
rect 4856 462544 4862 462596
rect 187234 462340 187240 462392
rect 187292 462380 187298 462392
rect 197446 462380 197452 462392
rect 187292 462352 197452 462380
rect 187292 462340 187298 462352
rect 197446 462340 197452 462352
rect 197504 462340 197510 462392
rect 358630 462340 358636 462392
rect 358688 462380 358694 462392
rect 360378 462380 360384 462392
rect 358688 462352 360384 462380
rect 358688 462340 358694 462352
rect 360378 462340 360384 462352
rect 360436 462340 360442 462392
rect 63218 461592 63224 461644
rect 63276 461632 63282 461644
rect 78766 461632 78772 461644
rect 63276 461604 78772 461632
rect 63276 461592 63282 461604
rect 78766 461592 78772 461604
rect 78824 461592 78830 461644
rect 76006 461456 76012 461508
rect 76064 461496 76070 461508
rect 76558 461496 76564 461508
rect 76064 461468 76564 461496
rect 76064 461456 76070 461468
rect 76558 461456 76564 461468
rect 76616 461456 76622 461508
rect 76558 460912 76564 460964
rect 76616 460952 76622 460964
rect 179414 460952 179420 460964
rect 76616 460924 179420 460952
rect 76616 460912 76622 460924
rect 179414 460912 179420 460924
rect 179472 460912 179478 460964
rect 191742 460844 191748 460896
rect 191800 460884 191806 460896
rect 197446 460884 197452 460896
rect 191800 460856 197452 460884
rect 191800 460844 191806 460856
rect 197446 460844 197452 460856
rect 197504 460844 197510 460896
rect 52362 460164 52368 460216
rect 52420 460204 52426 460216
rect 90450 460204 90456 460216
rect 52420 460176 90456 460204
rect 52420 460164 52426 460176
rect 90450 460164 90456 460176
rect 90508 460164 90514 460216
rect 166258 460164 166264 460216
rect 166316 460204 166322 460216
rect 191742 460204 191748 460216
rect 166316 460176 191748 460204
rect 166316 460164 166322 460176
rect 191742 460164 191748 460176
rect 191800 460164 191806 460216
rect 372982 460164 372988 460216
rect 373040 460204 373046 460216
rect 582558 460204 582564 460216
rect 373040 460176 582564 460204
rect 373040 460164 373046 460176
rect 582558 460164 582564 460176
rect 582616 460164 582622 460216
rect 56502 459552 56508 459604
rect 56560 459592 56566 459604
rect 67726 459592 67732 459604
rect 56560 459564 67732 459592
rect 56560 459552 56566 459564
rect 67726 459552 67732 459564
rect 67784 459552 67790 459604
rect 91094 459552 91100 459604
rect 91152 459592 91158 459604
rect 91554 459592 91560 459604
rect 91152 459564 91560 459592
rect 91152 459552 91158 459564
rect 91554 459552 91560 459564
rect 91612 459592 91618 459604
rect 159358 459592 159364 459604
rect 91612 459564 159364 459592
rect 91612 459552 91618 459564
rect 159358 459552 159364 459564
rect 159416 459552 159422 459604
rect 358722 459552 358728 459604
rect 358780 459592 358786 459604
rect 372706 459592 372712 459604
rect 358780 459564 372712 459592
rect 358780 459552 358786 459564
rect 372706 459552 372712 459564
rect 372764 459592 372770 459604
rect 372982 459592 372988 459604
rect 372764 459564 372988 459592
rect 372764 459552 372770 459564
rect 372982 459552 372988 459564
rect 373040 459552 373046 459604
rect 67726 458804 67732 458856
rect 67784 458844 67790 458856
rect 81434 458844 81440 458856
rect 67784 458816 81440 458844
rect 67784 458804 67790 458816
rect 81434 458804 81440 458816
rect 81492 458804 81498 458856
rect 91738 458804 91744 458856
rect 91796 458844 91802 458856
rect 120626 458844 120632 458856
rect 91796 458816 120632 458844
rect 91796 458804 91802 458816
rect 120626 458804 120632 458816
rect 120684 458804 120690 458856
rect 55122 457444 55128 457496
rect 55180 457484 55186 457496
rect 87598 457484 87604 457496
rect 55180 457456 87604 457484
rect 55180 457444 55186 457456
rect 87598 457444 87604 457456
rect 87656 457444 87662 457496
rect 115198 457444 115204 457496
rect 115256 457484 115262 457496
rect 126974 457484 126980 457496
rect 115256 457456 126980 457484
rect 115256 457444 115262 457456
rect 126974 457444 126980 457456
rect 127032 457444 127038 457496
rect 69014 456764 69020 456816
rect 69072 456804 69078 456816
rect 69842 456804 69848 456816
rect 69072 456776 69848 456804
rect 69072 456764 69078 456776
rect 69842 456764 69848 456776
rect 69900 456804 69906 456816
rect 157978 456804 157984 456816
rect 69900 456776 157984 456804
rect 69900 456764 69906 456776
rect 157978 456764 157984 456776
rect 158036 456764 158042 456816
rect 62022 456016 62028 456068
rect 62080 456056 62086 456068
rect 78674 456056 78680 456068
rect 62080 456028 78680 456056
rect 62080 456016 62086 456028
rect 78674 456016 78680 456028
rect 78732 456016 78738 456068
rect 108298 456016 108304 456068
rect 108356 456056 108362 456068
rect 127710 456056 127716 456068
rect 108356 456028 127716 456056
rect 108356 456016 108362 456028
rect 127710 456016 127716 456028
rect 127768 456016 127774 456068
rect 88334 455404 88340 455456
rect 88392 455444 88398 455456
rect 88978 455444 88984 455456
rect 88392 455416 88984 455444
rect 88392 455404 88398 455416
rect 88978 455404 88984 455416
rect 89036 455444 89042 455456
rect 125594 455444 125600 455456
rect 89036 455416 125600 455444
rect 89036 455404 89042 455416
rect 125594 455404 125600 455416
rect 125652 455404 125658 455456
rect 191282 455404 191288 455456
rect 191340 455444 191346 455456
rect 197446 455444 197452 455456
rect 191340 455416 197452 455444
rect 191340 455404 191346 455416
rect 197446 455404 197452 455416
rect 197504 455404 197510 455456
rect 358722 455404 358728 455456
rect 358780 455444 358786 455456
rect 376754 455444 376760 455456
rect 358780 455416 376760 455444
rect 358780 455404 358786 455416
rect 376754 455404 376760 455416
rect 376812 455444 376818 455456
rect 582374 455444 582380 455456
rect 376812 455416 582380 455444
rect 376812 455404 376818 455416
rect 582374 455404 582380 455416
rect 582432 455404 582438 455456
rect 14458 455336 14464 455388
rect 14516 455376 14522 455388
rect 111794 455376 111800 455388
rect 14516 455348 111800 455376
rect 14516 455336 14522 455348
rect 111794 455336 111800 455348
rect 111852 455336 111858 455388
rect 77294 455268 77300 455320
rect 77352 455308 77358 455320
rect 77938 455308 77944 455320
rect 77352 455280 77944 455308
rect 77352 455268 77358 455280
rect 77938 455268 77944 455280
rect 77996 455268 78002 455320
rect 63310 454656 63316 454708
rect 63368 454696 63374 454708
rect 67634 454696 67640 454708
rect 63368 454668 67640 454696
rect 63368 454656 63374 454668
rect 67634 454656 67640 454668
rect 67692 454656 67698 454708
rect 111794 454656 111800 454708
rect 111852 454696 111858 454708
rect 183554 454696 183560 454708
rect 111852 454668 183560 454696
rect 111852 454656 111858 454668
rect 183554 454656 183560 454668
rect 183612 454696 183618 454708
rect 184290 454696 184296 454708
rect 183612 454668 184296 454696
rect 183612 454656 183618 454668
rect 184290 454656 184296 454668
rect 184348 454656 184354 454708
rect 77294 454112 77300 454164
rect 77352 454152 77358 454164
rect 77352 454124 84194 454152
rect 77352 454112 77358 454124
rect 84166 454084 84194 454124
rect 132586 454084 132592 454096
rect 84166 454056 132592 454084
rect 132586 454044 132592 454056
rect 132644 454044 132650 454096
rect 193950 453500 193956 453552
rect 194008 453540 194014 453552
rect 197354 453540 197360 453552
rect 194008 453512 197360 453540
rect 194008 453500 194014 453512
rect 197354 453500 197360 453512
rect 197412 453500 197418 453552
rect 61746 453364 61752 453416
rect 61804 453404 61810 453416
rect 75914 453404 75920 453416
rect 61804 453376 75920 453404
rect 61804 453364 61810 453376
rect 75914 453364 75920 453376
rect 75972 453364 75978 453416
rect 57698 453296 57704 453348
rect 57756 453336 57762 453348
rect 72418 453336 72424 453348
rect 57756 453308 72424 453336
rect 57756 453296 57762 453308
rect 72418 453296 72424 453308
rect 72476 453296 72482 453348
rect 112438 453296 112444 453348
rect 112496 453336 112502 453348
rect 123018 453336 123024 453348
rect 112496 453308 123024 453336
rect 112496 453296 112502 453308
rect 123018 453296 123024 453308
rect 123076 453296 123082 453348
rect 125502 453296 125508 453348
rect 125560 453336 125566 453348
rect 151078 453336 151084 453348
rect 125560 453308 151084 453336
rect 125560 453296 125566 453308
rect 151078 453296 151084 453308
rect 151136 453296 151142 453348
rect 72694 452616 72700 452668
rect 72752 452656 72758 452668
rect 125502 452656 125508 452668
rect 72752 452628 125508 452656
rect 72752 452616 72758 452628
rect 125502 452616 125508 452628
rect 125560 452616 125566 452668
rect 358722 452616 358728 452668
rect 358780 452656 358786 452668
rect 377398 452656 377404 452668
rect 358780 452628 377404 452656
rect 358780 452616 358786 452628
rect 377398 452616 377404 452628
rect 377456 452616 377462 452668
rect 66162 451936 66168 451988
rect 66220 451976 66226 451988
rect 75178 451976 75184 451988
rect 66220 451948 75184 451976
rect 66220 451936 66226 451948
rect 75178 451936 75184 451948
rect 75236 451936 75242 451988
rect 116670 451936 116676 451988
rect 116728 451976 116734 451988
rect 124306 451976 124312 451988
rect 116728 451948 124312 451976
rect 116728 451936 116734 451948
rect 124306 451936 124312 451948
rect 124364 451936 124370 451988
rect 3418 451868 3424 451920
rect 3476 451908 3482 451920
rect 121454 451908 121460 451920
rect 3476 451880 121460 451908
rect 3476 451868 3482 451880
rect 121454 451868 121460 451880
rect 121512 451868 121518 451920
rect 95878 451188 95884 451240
rect 95936 451228 95942 451240
rect 127618 451228 127624 451240
rect 95936 451200 127624 451228
rect 95936 451188 95942 451200
rect 127618 451188 127624 451200
rect 127676 451188 127682 451240
rect 4798 450508 4804 450560
rect 4856 450548 4862 450560
rect 68094 450548 68100 450560
rect 4856 450520 68100 450548
rect 4856 450508 4862 450520
rect 68094 450508 68100 450520
rect 68152 450508 68158 450560
rect 50798 449964 50804 450016
rect 50856 450004 50862 450016
rect 74534 450004 74540 450016
rect 50856 449976 74540 450004
rect 50856 449964 50862 449976
rect 74534 449964 74540 449976
rect 74592 450004 74598 450016
rect 74810 450004 74816 450016
rect 74592 449976 74816 450004
rect 74592 449964 74598 449976
rect 74810 449964 74816 449976
rect 74868 449964 74874 450016
rect 68094 449896 68100 449948
rect 68152 449936 68158 449948
rect 68554 449936 68560 449948
rect 68152 449908 68560 449936
rect 68152 449896 68158 449908
rect 68554 449896 68560 449908
rect 68612 449936 68618 449948
rect 103514 449936 103520 449948
rect 68612 449908 103520 449936
rect 68612 449896 68618 449908
rect 103514 449896 103520 449908
rect 103572 449936 103578 449948
rect 103698 449936 103704 449948
rect 103572 449908 103704 449936
rect 103572 449896 103578 449908
rect 103698 449896 103704 449908
rect 103756 449896 103762 449948
rect 358722 449896 358728 449948
rect 358780 449936 358786 449948
rect 373994 449936 374000 449948
rect 358780 449908 374000 449936
rect 358780 449896 358786 449908
rect 373994 449896 374000 449908
rect 374052 449896 374058 449948
rect 39942 449828 39948 449880
rect 40000 449868 40006 449880
rect 72694 449868 72700 449880
rect 40000 449840 72700 449868
rect 40000 449828 40006 449840
rect 72694 449828 72700 449840
rect 72752 449828 72758 449880
rect 106918 449828 106924 449880
rect 106976 449868 106982 449880
rect 128998 449868 129004 449880
rect 106976 449840 129004 449868
rect 106976 449828 106982 449840
rect 128998 449828 129004 449840
rect 129056 449828 129062 449880
rect 50890 449148 50896 449200
rect 50948 449188 50954 449200
rect 80882 449188 80888 449200
rect 50948 449160 80888 449188
rect 50948 449148 50954 449160
rect 80882 449148 80888 449160
rect 80940 449148 80946 449200
rect 100662 449148 100668 449200
rect 100720 449188 100726 449200
rect 108298 449188 108304 449200
rect 100720 449160 108304 449188
rect 100720 449148 100726 449160
rect 108298 449148 108304 449160
rect 108356 449148 108362 449200
rect 371510 449148 371516 449200
rect 371568 449188 371574 449200
rect 582650 449188 582656 449200
rect 371568 449160 582656 449188
rect 371568 449148 371574 449160
rect 582650 449148 582656 449160
rect 582708 449148 582714 449200
rect 116578 448604 116584 448656
rect 116636 448644 116642 448656
rect 120718 448644 120724 448656
rect 116636 448616 120724 448644
rect 116636 448604 116642 448616
rect 120718 448604 120724 448616
rect 120776 448604 120782 448656
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 25498 448576 25504 448588
rect 3200 448548 25504 448576
rect 3200 448536 3206 448548
rect 25498 448536 25504 448548
rect 25556 448536 25562 448588
rect 72694 448536 72700 448588
rect 72752 448576 72758 448588
rect 73154 448576 73160 448588
rect 72752 448548 73160 448576
rect 72752 448536 72758 448548
rect 73154 448536 73160 448548
rect 73212 448536 73218 448588
rect 190270 448536 190276 448588
rect 190328 448576 190334 448588
rect 197354 448576 197360 448588
rect 190328 448548 197360 448576
rect 190328 448536 190334 448548
rect 197354 448536 197360 448548
rect 197412 448536 197418 448588
rect 358722 448536 358728 448588
rect 358780 448576 358786 448588
rect 371326 448576 371332 448588
rect 358780 448548 371332 448576
rect 358780 448536 358786 448548
rect 371326 448536 371332 448548
rect 371384 448576 371390 448588
rect 371510 448576 371516 448588
rect 371384 448548 371516 448576
rect 371384 448536 371390 448548
rect 371510 448536 371516 448548
rect 371568 448536 371574 448588
rect 94498 448468 94504 448520
rect 94556 448508 94562 448520
rect 187234 448508 187240 448520
rect 94556 448480 187240 448508
rect 94556 448468 94562 448480
rect 187234 448468 187240 448480
rect 187292 448468 187298 448520
rect 64598 447788 64604 447840
rect 64656 447828 64662 447840
rect 71038 447828 71044 447840
rect 64656 447800 71044 447828
rect 64656 447788 64662 447800
rect 71038 447788 71044 447800
rect 71096 447788 71102 447840
rect 11698 447108 11704 447160
rect 11756 447148 11762 447160
rect 12342 447148 12348 447160
rect 11756 447120 12348 447148
rect 11756 447108 11762 447120
rect 12342 447108 12348 447120
rect 12400 447148 12406 447160
rect 125686 447148 125692 447160
rect 12400 447120 125692 447148
rect 12400 447108 12406 447120
rect 125686 447108 125692 447120
rect 125744 447108 125750 447160
rect 109678 447040 109684 447092
rect 109736 447080 109742 447092
rect 146938 447080 146944 447092
rect 109736 447052 146944 447080
rect 109736 447040 109742 447052
rect 146938 447040 146944 447052
rect 146996 447040 147002 447092
rect 65978 446360 65984 446412
rect 66036 446400 66042 446412
rect 73246 446400 73252 446412
rect 66036 446372 73252 446400
rect 66036 446360 66042 446372
rect 73246 446360 73252 446372
rect 73304 446360 73310 446412
rect 98638 445816 98644 445868
rect 98696 445856 98702 445868
rect 100478 445856 100484 445868
rect 98696 445828 100484 445856
rect 98696 445816 98702 445828
rect 100478 445816 100484 445828
rect 100536 445856 100542 445868
rect 102226 445856 102232 445868
rect 100536 445828 102232 445856
rect 100536 445816 100542 445828
rect 102226 445816 102232 445828
rect 102284 445816 102290 445868
rect 7558 445748 7564 445800
rect 7616 445788 7622 445800
rect 118694 445788 118700 445800
rect 7616 445760 118700 445788
rect 7616 445748 7622 445760
rect 118694 445748 118700 445760
rect 118752 445748 118758 445800
rect 174630 445748 174636 445800
rect 174688 445788 174694 445800
rect 197354 445788 197360 445800
rect 174688 445760 197360 445788
rect 174688 445748 174694 445760
rect 197354 445748 197360 445760
rect 197412 445748 197418 445800
rect 358722 445748 358728 445800
rect 358780 445788 358786 445800
rect 369946 445788 369952 445800
rect 358780 445760 369952 445788
rect 358780 445748 358786 445760
rect 369946 445748 369952 445760
rect 370004 445748 370010 445800
rect 67634 445680 67640 445732
rect 67692 445720 67698 445732
rect 68738 445720 68744 445732
rect 67692 445692 68744 445720
rect 67692 445680 67698 445692
rect 68738 445680 68744 445692
rect 68796 445680 68802 445732
rect 119338 444524 119344 444576
rect 119396 444564 119402 444576
rect 120902 444564 120908 444576
rect 119396 444536 120908 444564
rect 119396 444524 119402 444536
rect 120902 444524 120908 444536
rect 120960 444524 120966 444576
rect 53558 444456 53564 444508
rect 53616 444496 53622 444508
rect 85574 444496 85580 444508
rect 53616 444468 85580 444496
rect 53616 444456 53622 444468
rect 85574 444456 85580 444468
rect 85632 444456 85638 444508
rect 100754 444456 100760 444508
rect 100812 444496 100818 444508
rect 127618 444496 127624 444508
rect 100812 444468 127624 444496
rect 100812 444456 100818 444468
rect 127618 444456 127624 444468
rect 127676 444456 127682 444508
rect 68922 444388 68928 444440
rect 68980 444428 68986 444440
rect 146938 444428 146944 444440
rect 68980 444400 146944 444428
rect 68980 444388 68986 444400
rect 146938 444388 146944 444400
rect 146996 444388 147002 444440
rect 166902 443708 166908 443760
rect 166960 443748 166966 443760
rect 197354 443748 197360 443760
rect 166960 443720 197360 443748
rect 166960 443708 166966 443720
rect 197354 443708 197360 443720
rect 197412 443708 197418 443760
rect 124122 443640 124128 443692
rect 124180 443680 124186 443692
rect 126974 443680 126980 443692
rect 124180 443652 126980 443680
rect 124180 443640 124186 443652
rect 126974 443640 126980 443652
rect 127032 443680 127038 443692
rect 169754 443680 169760 443692
rect 127032 443652 169760 443680
rect 127032 443640 127038 443652
rect 169754 443640 169760 443652
rect 169812 443680 169818 443692
rect 192570 443680 192576 443692
rect 169812 443652 192576 443680
rect 169812 443640 169818 443652
rect 192570 443640 192576 443652
rect 192628 443640 192634 443692
rect 358722 442960 358728 443012
rect 358780 443000 358786 443012
rect 361666 443000 361672 443012
rect 358780 442972 361672 443000
rect 358780 442960 358786 442972
rect 361666 442960 361672 442972
rect 361724 442960 361730 443012
rect 48130 442892 48136 442944
rect 48188 442932 48194 442944
rect 67726 442932 67732 442944
rect 48188 442904 67732 442932
rect 48188 442892 48194 442904
rect 67726 442892 67732 442904
rect 67784 442892 67790 442944
rect 124122 441600 124128 441652
rect 124180 441640 124186 441652
rect 140038 441640 140044 441652
rect 124180 441612 140044 441640
rect 124180 441600 124186 441612
rect 140038 441600 140044 441612
rect 140096 441600 140102 441652
rect 192662 441396 192668 441448
rect 192720 441436 192726 441448
rect 197722 441436 197728 441448
rect 192720 441408 197728 441436
rect 192720 441396 192726 441408
rect 197722 441396 197728 441408
rect 197780 441396 197786 441448
rect 60458 440240 60464 440292
rect 60516 440280 60522 440292
rect 66898 440280 66904 440292
rect 60516 440252 66904 440280
rect 60516 440240 60522 440252
rect 66898 440240 66904 440252
rect 66956 440240 66962 440292
rect 121454 440172 121460 440224
rect 121512 440212 121518 440224
rect 130562 440212 130568 440224
rect 121512 440184 130568 440212
rect 121512 440172 121518 440184
rect 130562 440172 130568 440184
rect 130620 440172 130626 440224
rect 358722 438880 358728 438932
rect 358780 438920 358786 438932
rect 376018 438920 376024 438932
rect 358780 438892 376024 438920
rect 358780 438880 358786 438892
rect 376018 438880 376024 438892
rect 376076 438880 376082 438932
rect 63310 437520 63316 437572
rect 63368 437560 63374 437572
rect 64782 437560 64788 437572
rect 63368 437532 64788 437560
rect 63368 437520 63374 437532
rect 64782 437520 64788 437532
rect 64840 437560 64846 437572
rect 66898 437560 66904 437572
rect 64840 437532 66904 437560
rect 64840 437520 64846 437532
rect 66898 437520 66904 437532
rect 66956 437520 66962 437572
rect 124122 437452 124128 437504
rect 124180 437492 124186 437504
rect 128354 437492 128360 437504
rect 124180 437464 128360 437492
rect 124180 437452 124186 437464
rect 128354 437452 128360 437464
rect 128412 437492 128418 437504
rect 128998 437492 129004 437504
rect 128412 437464 129004 437492
rect 128412 437452 128418 437464
rect 128998 437452 129004 437464
rect 129056 437452 129062 437504
rect 155770 437384 155776 437436
rect 155828 437424 155834 437436
rect 162118 437424 162124 437436
rect 155828 437396 162124 437424
rect 155828 437384 155834 437396
rect 162118 437384 162124 437396
rect 162176 437384 162182 437436
rect 162762 436092 162768 436144
rect 162820 436132 162826 436144
rect 197354 436132 197360 436144
rect 162820 436104 197360 436132
rect 162820 436092 162826 436104
rect 197354 436092 197360 436104
rect 197412 436092 197418 436144
rect 358722 436092 358728 436144
rect 358780 436132 358786 436144
rect 363138 436132 363144 436144
rect 358780 436104 363144 436132
rect 358780 436092 358786 436104
rect 363138 436092 363144 436104
rect 363196 436092 363202 436144
rect 53650 436024 53656 436076
rect 53708 436064 53714 436076
rect 57882 436064 57888 436076
rect 53708 436036 57888 436064
rect 53708 436024 53714 436036
rect 57882 436024 57888 436036
rect 57940 436024 57946 436076
rect 155310 436024 155316 436076
rect 155368 436064 155374 436076
rect 156598 436064 156604 436076
rect 155368 436036 156604 436064
rect 155368 436024 155374 436036
rect 156598 436024 156604 436036
rect 156656 436024 156662 436076
rect 57882 434732 57888 434784
rect 57940 434772 57946 434784
rect 66898 434772 66904 434784
rect 57940 434744 66904 434772
rect 57940 434732 57946 434744
rect 66898 434732 66904 434744
rect 66956 434732 66962 434784
rect 120718 434732 120724 434784
rect 120776 434772 120782 434784
rect 128354 434772 128360 434784
rect 120776 434744 128360 434772
rect 120776 434732 120782 434744
rect 128354 434732 128360 434744
rect 128412 434732 128418 434784
rect 165614 434664 165620 434716
rect 165672 434704 165678 434716
rect 166258 434704 166264 434716
rect 165672 434676 166264 434704
rect 165672 434664 165678 434676
rect 166258 434664 166264 434676
rect 166316 434664 166322 434716
rect 127710 433984 127716 434036
rect 127768 434024 127774 434036
rect 165614 434024 165620 434036
rect 127768 433996 165620 434024
rect 127768 433984 127774 433996
rect 165614 433984 165620 433996
rect 165672 433984 165678 434036
rect 46842 433304 46848 433356
rect 46900 433344 46906 433356
rect 46900 433316 55214 433344
rect 46900 433304 46906 433316
rect 55186 433276 55214 433316
rect 179322 433304 179328 433356
rect 179380 433344 179386 433356
rect 197354 433344 197360 433356
rect 179380 433316 197360 433344
rect 179380 433304 179386 433316
rect 197354 433304 197360 433316
rect 197412 433304 197418 433356
rect 358722 433304 358728 433356
rect 358780 433344 358786 433356
rect 365806 433344 365812 433356
rect 358780 433316 365812 433344
rect 358780 433304 358786 433316
rect 365806 433304 365812 433316
rect 365864 433304 365870 433356
rect 55858 433276 55864 433288
rect 55186 433248 55864 433276
rect 55858 433236 55864 433248
rect 55916 433276 55922 433288
rect 66806 433276 66812 433288
rect 55916 433248 66812 433276
rect 55916 433236 55922 433248
rect 66806 433236 66812 433248
rect 66864 433236 66870 433288
rect 124122 433236 124128 433288
rect 124180 433276 124186 433288
rect 127710 433276 127716 433288
rect 124180 433248 127716 433276
rect 124180 433236 124186 433248
rect 127710 433236 127716 433248
rect 127768 433236 127774 433288
rect 52270 431196 52276 431248
rect 52328 431236 52334 431248
rect 65886 431236 65892 431248
rect 52328 431208 65892 431236
rect 52328 431196 52334 431208
rect 65886 431196 65892 431208
rect 65944 431236 65950 431248
rect 66530 431236 66536 431248
rect 65944 431208 66536 431236
rect 65944 431196 65950 431208
rect 66530 431196 66536 431208
rect 66588 431196 66594 431248
rect 124122 430584 124128 430636
rect 124180 430624 124186 430636
rect 172422 430624 172428 430636
rect 124180 430596 172428 430624
rect 124180 430584 124186 430596
rect 172422 430584 172428 430596
rect 172480 430624 172486 430636
rect 173250 430624 173256 430636
rect 172480 430596 173256 430624
rect 172480 430584 172486 430596
rect 173250 430584 173256 430596
rect 173308 430584 173314 430636
rect 36722 429088 36728 429140
rect 36780 429128 36786 429140
rect 37182 429128 37188 429140
rect 36780 429100 37188 429128
rect 36780 429088 36786 429100
rect 37182 429088 37188 429100
rect 37240 429128 37246 429140
rect 66714 429128 66720 429140
rect 37240 429100 66720 429128
rect 37240 429088 37246 429100
rect 66714 429088 66720 429100
rect 66772 429088 66778 429140
rect 121454 429088 121460 429140
rect 121512 429128 121518 429140
rect 177298 429128 177304 429140
rect 121512 429100 177304 429128
rect 121512 429088 121518 429100
rect 177298 429088 177304 429100
rect 177356 429088 177362 429140
rect 14458 428408 14464 428460
rect 14516 428448 14522 428460
rect 36722 428448 36728 428460
rect 14516 428420 36728 428448
rect 14516 428408 14522 428420
rect 36722 428408 36728 428420
rect 36780 428408 36786 428460
rect 192570 427796 192576 427848
rect 192628 427836 192634 427848
rect 197354 427836 197360 427848
rect 192628 427808 197360 427836
rect 192628 427796 192634 427808
rect 197354 427796 197360 427808
rect 197412 427796 197418 427848
rect 358722 427796 358728 427848
rect 358780 427836 358786 427848
rect 363230 427836 363236 427848
rect 358780 427808 363236 427836
rect 358780 427796 358786 427808
rect 363230 427796 363236 427808
rect 363288 427796 363294 427848
rect 137278 426436 137284 426488
rect 137336 426476 137342 426488
rect 197354 426476 197360 426488
rect 137336 426448 197360 426476
rect 137336 426436 137342 426448
rect 197354 426436 197360 426448
rect 197412 426436 197418 426488
rect 358722 426436 358728 426488
rect 358780 426476 358786 426488
rect 372614 426476 372620 426488
rect 358780 426448 372620 426476
rect 358780 426436 358786 426448
rect 372614 426436 372620 426448
rect 372672 426436 372678 426488
rect 41322 425688 41328 425740
rect 41380 425728 41386 425740
rect 59078 425728 59084 425740
rect 41380 425700 59084 425728
rect 41380 425688 41386 425700
rect 59078 425688 59084 425700
rect 59136 425688 59142 425740
rect 59078 425076 59084 425128
rect 59136 425116 59142 425128
rect 66254 425116 66260 425128
rect 59136 425088 66260 425116
rect 59136 425076 59142 425088
rect 66254 425076 66260 425088
rect 66312 425076 66318 425128
rect 61838 423648 61844 423700
rect 61896 423688 61902 423700
rect 66070 423688 66076 423700
rect 61896 423660 66076 423688
rect 61896 423648 61902 423660
rect 66070 423648 66076 423660
rect 66128 423648 66134 423700
rect 167730 423648 167736 423700
rect 167788 423688 167794 423700
rect 197354 423688 197360 423700
rect 167788 423660 197360 423688
rect 167788 423648 167794 423660
rect 197354 423648 197360 423660
rect 197412 423648 197418 423700
rect 3418 423580 3424 423632
rect 3476 423620 3482 423632
rect 11698 423620 11704 423632
rect 3476 423592 11704 423620
rect 3476 423580 3482 423592
rect 11698 423580 11704 423592
rect 11756 423580 11762 423632
rect 124122 422220 124128 422272
rect 124180 422260 124186 422272
rect 136634 422260 136640 422272
rect 124180 422232 136640 422260
rect 124180 422220 124186 422232
rect 136634 422220 136640 422232
rect 136692 422220 136698 422272
rect 52270 421540 52276 421592
rect 52328 421580 52334 421592
rect 59170 421580 59176 421592
rect 52328 421552 59176 421580
rect 52328 421540 52334 421552
rect 59170 421540 59176 421552
rect 59228 421580 59234 421592
rect 66254 421580 66260 421592
rect 59228 421552 66260 421580
rect 59228 421540 59234 421552
rect 66254 421540 66260 421552
rect 66312 421540 66318 421592
rect 136634 421540 136640 421592
rect 136692 421580 136698 421592
rect 162670 421580 162676 421592
rect 136692 421552 162676 421580
rect 136692 421540 136698 421552
rect 162670 421540 162676 421552
rect 162728 421580 162734 421592
rect 178770 421580 178776 421592
rect 162728 421552 178776 421580
rect 162728 421540 162734 421552
rect 178770 421540 178776 421552
rect 178828 421540 178834 421592
rect 123018 420860 123024 420912
rect 123076 420900 123082 420912
rect 170490 420900 170496 420912
rect 123076 420872 170496 420900
rect 123076 420860 123082 420872
rect 170490 420860 170496 420872
rect 170548 420860 170554 420912
rect 43990 418752 43996 418804
rect 44048 418792 44054 418804
rect 59170 418792 59176 418804
rect 44048 418764 59176 418792
rect 44048 418752 44054 418764
rect 59170 418752 59176 418764
rect 59228 418752 59234 418804
rect 176194 418140 176200 418192
rect 176252 418180 176258 418192
rect 197354 418180 197360 418192
rect 176252 418152 197360 418180
rect 176252 418140 176258 418152
rect 197354 418140 197360 418152
rect 197412 418140 197418 418192
rect 358722 418140 358728 418192
rect 358780 418180 358786 418192
rect 361758 418180 361764 418192
rect 358780 418152 361764 418180
rect 358780 418140 358786 418152
rect 361758 418140 361764 418152
rect 361816 418140 361822 418192
rect 59170 416780 59176 416832
rect 59228 416820 59234 416832
rect 66898 416820 66904 416832
rect 59228 416792 66904 416820
rect 59228 416780 59234 416792
rect 66898 416780 66904 416792
rect 66956 416780 66962 416832
rect 358722 416780 358728 416832
rect 358780 416820 358786 416832
rect 368474 416820 368480 416832
rect 358780 416792 368480 416820
rect 358780 416780 358786 416792
rect 368474 416780 368480 416792
rect 368532 416780 368538 416832
rect 57790 416032 57796 416084
rect 57848 416072 57854 416084
rect 66254 416072 66260 416084
rect 57848 416044 66260 416072
rect 57848 416032 57854 416044
rect 66254 416032 66260 416044
rect 66312 416032 66318 416084
rect 57790 414672 57796 414724
rect 57848 414712 57854 414724
rect 66254 414712 66260 414724
rect 57848 414684 66260 414712
rect 57848 414672 57854 414684
rect 66254 414672 66260 414684
rect 66312 414672 66318 414724
rect 124122 414672 124128 414724
rect 124180 414712 124186 414724
rect 138014 414712 138020 414724
rect 124180 414684 138020 414712
rect 124180 414672 124186 414684
rect 138014 414672 138020 414684
rect 138072 414672 138078 414724
rect 181438 413992 181444 414044
rect 181496 414032 181502 414044
rect 197354 414032 197360 414044
rect 181496 414004 197360 414032
rect 181496 413992 181502 414004
rect 197354 413992 197360 414004
rect 197412 413992 197418 414044
rect 358722 413992 358728 414044
rect 358780 414032 358786 414044
rect 370038 414032 370044 414044
rect 358780 414004 370044 414032
rect 358780 413992 358786 414004
rect 370038 413992 370044 414004
rect 370096 413992 370102 414044
rect 122834 413244 122840 413296
rect 122892 413284 122898 413296
rect 133874 413284 133880 413296
rect 122892 413256 133880 413284
rect 122892 413244 122898 413256
rect 133874 413244 133880 413256
rect 133932 413244 133938 413296
rect 161382 411272 161388 411324
rect 161440 411312 161446 411324
rect 197354 411312 197360 411324
rect 161440 411284 197360 411312
rect 161440 411272 161446 411284
rect 197354 411272 197360 411284
rect 197412 411272 197418 411324
rect 358722 411272 358728 411324
rect 358780 411312 358786 411324
rect 378226 411312 378232 411324
rect 358780 411284 378232 411312
rect 358780 411272 358786 411284
rect 378226 411272 378232 411284
rect 378284 411272 378290 411324
rect 121178 409844 121184 409896
rect 121236 409884 121242 409896
rect 151078 409884 151084 409896
rect 121236 409856 151084 409884
rect 121236 409844 121242 409856
rect 151078 409844 151084 409856
rect 151136 409844 151142 409896
rect 130378 409776 130384 409828
rect 130436 409816 130442 409828
rect 197354 409816 197360 409828
rect 130436 409788 197360 409816
rect 130436 409776 130442 409788
rect 197354 409776 197360 409788
rect 197412 409776 197418 409828
rect 124122 408416 124128 408468
rect 124180 408456 124186 408468
rect 133782 408456 133788 408468
rect 124180 408428 133788 408456
rect 124180 408416 124186 408428
rect 133782 408416 133788 408428
rect 133840 408456 133846 408468
rect 134610 408456 134616 408468
rect 133840 408428 134616 408456
rect 133840 408416 133846 408428
rect 134610 408416 134616 408428
rect 134668 408416 134674 408468
rect 60642 407124 60648 407176
rect 60700 407164 60706 407176
rect 66346 407164 66352 407176
rect 60700 407136 66352 407164
rect 60700 407124 60706 407136
rect 66346 407124 66352 407136
rect 66404 407124 66410 407176
rect 124306 405968 124312 406020
rect 124364 406008 124370 406020
rect 124858 406008 124864 406020
rect 124364 405980 124864 406008
rect 124364 405968 124370 405980
rect 124858 405968 124864 405980
rect 124916 405968 124922 406020
rect 59262 405764 59268 405816
rect 59320 405804 59326 405816
rect 63126 405804 63132 405816
rect 59320 405776 63132 405804
rect 59320 405764 59326 405776
rect 63126 405764 63132 405776
rect 63184 405804 63190 405816
rect 66806 405804 66812 405816
rect 63184 405776 66812 405804
rect 63184 405764 63190 405776
rect 66806 405764 66812 405776
rect 66864 405764 66870 405816
rect 133138 405696 133144 405748
rect 133196 405736 133202 405748
rect 197354 405736 197360 405748
rect 133196 405708 197360 405736
rect 133196 405696 133202 405708
rect 197354 405696 197360 405708
rect 197412 405696 197418 405748
rect 358722 405696 358728 405748
rect 358780 405736 358786 405748
rect 364518 405736 364524 405748
rect 358780 405708 364524 405736
rect 358780 405696 358786 405708
rect 364518 405696 364524 405708
rect 364576 405696 364582 405748
rect 189810 404336 189816 404388
rect 189868 404376 189874 404388
rect 197354 404376 197360 404388
rect 189868 404348 197360 404376
rect 189868 404336 189874 404348
rect 197354 404336 197360 404348
rect 197412 404336 197418 404388
rect 122926 403520 122932 403572
rect 122984 403560 122990 403572
rect 125042 403560 125048 403572
rect 122984 403532 125048 403560
rect 122984 403520 122990 403532
rect 125042 403520 125048 403532
rect 125100 403520 125106 403572
rect 66622 403152 66628 403164
rect 57946 403124 66628 403152
rect 48130 402908 48136 402960
rect 48188 402948 48194 402960
rect 52178 402948 52184 402960
rect 48188 402920 52184 402948
rect 48188 402908 48194 402920
rect 52178 402908 52184 402920
rect 52236 402908 52242 402960
rect 52178 402228 52184 402280
rect 52236 402268 52242 402280
rect 57946 402268 57974 403124
rect 66622 403112 66628 403124
rect 66680 403112 66686 403164
rect 358722 402976 358728 403028
rect 358780 403016 358786 403028
rect 365898 403016 365904 403028
rect 358780 402988 365904 403016
rect 358780 402976 358786 402988
rect 365898 402976 365904 402988
rect 365956 402976 365962 403028
rect 52236 402240 57974 402268
rect 52236 402228 52242 402240
rect 122098 401616 122104 401668
rect 122156 401656 122162 401668
rect 122926 401656 122932 401668
rect 122156 401628 122932 401656
rect 122156 401616 122162 401628
rect 122926 401616 122932 401628
rect 122984 401616 122990 401668
rect 358722 401616 358728 401668
rect 358780 401656 358786 401668
rect 416774 401656 416780 401668
rect 358780 401628 416780 401656
rect 358780 401616 358786 401628
rect 416774 401616 416780 401628
rect 416832 401616 416838 401668
rect 166902 400936 166908 400988
rect 166960 400976 166966 400988
rect 178034 400976 178040 400988
rect 166960 400948 178040 400976
rect 166960 400936 166966 400948
rect 178034 400936 178040 400948
rect 178092 400936 178098 400988
rect 50890 400868 50896 400920
rect 50948 400908 50954 400920
rect 66806 400908 66812 400920
rect 50948 400880 66812 400908
rect 50948 400868 50954 400880
rect 66806 400868 66812 400880
rect 66864 400868 66870 400920
rect 123938 400868 123944 400920
rect 123996 400908 124002 400920
rect 193950 400908 193956 400920
rect 123996 400880 193956 400908
rect 123996 400868 124002 400880
rect 193950 400868 193956 400880
rect 194008 400868 194014 400920
rect 55030 399440 55036 399492
rect 55088 399480 55094 399492
rect 66806 399480 66812 399492
rect 55088 399452 66812 399480
rect 55088 399440 55094 399452
rect 66806 399440 66812 399452
rect 66864 399440 66870 399492
rect 124122 399440 124128 399492
rect 124180 399480 124186 399492
rect 125686 399480 125692 399492
rect 124180 399452 125692 399480
rect 124180 399440 124186 399452
rect 125686 399440 125692 399452
rect 125744 399480 125750 399492
rect 192662 399480 192668 399492
rect 125744 399452 192668 399480
rect 125744 399440 125750 399452
rect 192662 399440 192668 399452
rect 192720 399440 192726 399492
rect 194042 398828 194048 398880
rect 194100 398868 194106 398880
rect 197354 398868 197360 398880
rect 194100 398840 197360 398868
rect 194100 398828 194106 398840
rect 197354 398828 197360 398840
rect 197412 398828 197418 398880
rect 358630 398828 358636 398880
rect 358688 398868 358694 398880
rect 361850 398868 361856 398880
rect 358688 398840 361856 398868
rect 358688 398828 358694 398840
rect 361850 398828 361856 398840
rect 361908 398828 361914 398880
rect 3510 397536 3516 397588
rect 3568 397576 3574 397588
rect 7558 397576 7564 397588
rect 3568 397548 7564 397576
rect 3568 397536 3574 397548
rect 7558 397536 7564 397548
rect 7616 397536 7622 397588
rect 124122 396924 124128 396976
rect 124180 396964 124186 396976
rect 129734 396964 129740 396976
rect 124180 396936 129740 396964
rect 124180 396924 124186 396936
rect 129734 396924 129740 396936
rect 129792 396924 129798 396976
rect 35802 396720 35808 396772
rect 35860 396760 35866 396772
rect 66990 396760 66996 396772
rect 35860 396732 66996 396760
rect 35860 396720 35866 396732
rect 66990 396720 66996 396732
rect 67048 396720 67054 396772
rect 140038 396720 140044 396772
rect 140096 396760 140102 396772
rect 164878 396760 164884 396772
rect 140096 396732 164884 396760
rect 140096 396720 140102 396732
rect 164878 396720 164884 396732
rect 164936 396720 164942 396772
rect 59170 395972 59176 396024
rect 59228 396012 59234 396024
rect 66070 396012 66076 396024
rect 59228 395984 66076 396012
rect 59228 395972 59234 395984
rect 66070 395972 66076 395984
rect 66128 395972 66134 396024
rect 125502 395292 125508 395344
rect 125560 395332 125566 395344
rect 148410 395332 148416 395344
rect 125560 395304 148416 395332
rect 125560 395292 125566 395304
rect 148410 395292 148416 395304
rect 148468 395292 148474 395344
rect 171042 394680 171048 394732
rect 171100 394720 171106 394732
rect 197354 394720 197360 394732
rect 171100 394692 197360 394720
rect 171100 394680 171106 394692
rect 197354 394680 197360 394692
rect 197412 394680 197418 394732
rect 120718 393932 120724 393984
rect 120776 393972 120782 393984
rect 120902 393972 120908 393984
rect 120776 393944 120908 393972
rect 120776 393932 120782 393944
rect 120902 393932 120908 393944
rect 120960 393932 120966 393984
rect 129734 393932 129740 393984
rect 129792 393972 129798 393984
rect 177390 393972 177396 393984
rect 129792 393944 177396 393972
rect 129792 393932 129798 393944
rect 177390 393932 177396 393944
rect 177448 393932 177454 393984
rect 356330 393320 356336 393372
rect 356388 393360 356394 393372
rect 393314 393360 393320 393372
rect 356388 393332 393320 393360
rect 356388 393320 356394 393332
rect 393314 393320 393320 393332
rect 393372 393320 393378 393372
rect 48222 393252 48228 393304
rect 48280 393292 48286 393304
rect 65794 393292 65800 393304
rect 48280 393264 65800 393292
rect 48280 393252 48286 393264
rect 65794 393252 65800 393264
rect 65852 393252 65858 393304
rect 123754 392368 123760 392420
rect 123812 392408 123818 392420
rect 131758 392408 131764 392420
rect 123812 392380 131764 392408
rect 123812 392368 123818 392380
rect 131758 392368 131764 392380
rect 131816 392368 131822 392420
rect 130378 391960 130384 392012
rect 130436 392000 130442 392012
rect 180150 392000 180156 392012
rect 130436 391972 180156 392000
rect 130436 391960 130442 391972
rect 180150 391960 180156 391972
rect 180208 391960 180214 392012
rect 145558 391252 145564 391264
rect 74506 391224 145564 391252
rect 73062 391008 73068 391060
rect 73120 391048 73126 391060
rect 74506 391048 74534 391224
rect 145558 391212 145564 391224
rect 145616 391212 145622 391264
rect 73120 391020 74534 391048
rect 73120 391008 73126 391020
rect 72050 390532 72056 390584
rect 72108 390572 72114 390584
rect 73062 390572 73068 390584
rect 72108 390544 73068 390572
rect 72108 390532 72114 390544
rect 73062 390532 73068 390544
rect 73120 390532 73126 390584
rect 131114 390532 131120 390584
rect 131172 390572 131178 390584
rect 132402 390572 132408 390584
rect 131172 390544 132408 390572
rect 131172 390532 131178 390544
rect 132402 390532 132408 390544
rect 132460 390572 132466 390584
rect 168374 390572 168380 390584
rect 132460 390544 168380 390572
rect 132460 390532 132466 390544
rect 168374 390532 168380 390544
rect 168432 390532 168438 390584
rect 66070 390464 66076 390516
rect 66128 390504 66134 390516
rect 197354 390504 197360 390516
rect 66128 390476 197360 390504
rect 66128 390464 66134 390476
rect 197354 390464 197360 390476
rect 197412 390464 197418 390516
rect 65978 389172 65984 389224
rect 66036 389212 66042 389224
rect 77846 389212 77852 389224
rect 66036 389184 77852 389212
rect 66036 389172 66042 389184
rect 77846 389172 77852 389184
rect 77904 389212 77910 389224
rect 131114 389212 131120 389224
rect 77904 389184 131120 389212
rect 77904 389172 77910 389184
rect 131114 389172 131120 389184
rect 131172 389172 131178 389224
rect 64598 389104 64604 389156
rect 64656 389144 64662 389156
rect 73154 389144 73160 389156
rect 64656 389116 73160 389144
rect 64656 389104 64662 389116
rect 73154 389104 73160 389116
rect 73212 389104 73218 389156
rect 115198 389104 115204 389156
rect 115256 389144 115262 389156
rect 120442 389144 120448 389156
rect 115256 389116 120448 389144
rect 115256 389104 115262 389116
rect 120442 389104 120448 389116
rect 120500 389104 120506 389156
rect 96246 388492 96252 388544
rect 96304 388532 96310 388544
rect 188798 388532 188804 388544
rect 96304 388504 188804 388532
rect 96304 388492 96310 388504
rect 188798 388492 188804 388504
rect 188856 388532 188862 388544
rect 194042 388532 194048 388544
rect 188856 388504 194048 388532
rect 188856 388492 188862 388504
rect 194042 388492 194048 388504
rect 194100 388492 194106 388544
rect 15838 388424 15844 388476
rect 15896 388464 15902 388476
rect 110322 388464 110328 388476
rect 15896 388436 110328 388464
rect 15896 388424 15902 388436
rect 110322 388424 110328 388436
rect 110380 388424 110386 388476
rect 88518 387812 88524 387864
rect 88576 387852 88582 387864
rect 90358 387852 90364 387864
rect 88576 387824 90364 387852
rect 88576 387812 88582 387824
rect 90358 387812 90364 387824
rect 90416 387812 90422 387864
rect 110322 387812 110328 387864
rect 110380 387852 110386 387864
rect 111426 387852 111432 387864
rect 110380 387824 111432 387852
rect 110380 387812 110386 387824
rect 111426 387812 111432 387824
rect 111484 387812 111490 387864
rect 123478 387812 123484 387864
rect 123536 387852 123542 387864
rect 162118 387852 162124 387864
rect 123536 387824 162124 387852
rect 123536 387812 123542 387824
rect 162118 387812 162124 387824
rect 162176 387812 162182 387864
rect 64782 387064 64788 387116
rect 64840 387104 64846 387116
rect 68738 387104 68744 387116
rect 64840 387076 68744 387104
rect 64840 387064 64846 387076
rect 68738 387064 68744 387076
rect 68796 387064 68802 387116
rect 113082 387064 113088 387116
rect 113140 387104 113146 387116
rect 120902 387104 120908 387116
rect 113140 387076 120908 387104
rect 113140 387064 113146 387076
rect 120902 387064 120908 387076
rect 120960 387064 120966 387116
rect 7558 386384 7564 386436
rect 7616 386424 7622 386436
rect 117314 386424 117320 386436
rect 7616 386396 117320 386424
rect 7616 386384 7622 386396
rect 117314 386384 117320 386396
rect 117372 386424 117378 386436
rect 117958 386424 117964 386436
rect 117372 386396 117964 386424
rect 117372 386384 117378 386396
rect 117958 386384 117964 386396
rect 118016 386384 118022 386436
rect 191190 386384 191196 386436
rect 191248 386424 191254 386436
rect 197354 386424 197360 386436
rect 191248 386396 197360 386424
rect 191248 386384 191254 386396
rect 197354 386384 197360 386396
rect 197412 386384 197418 386436
rect 62022 386316 62028 386368
rect 62080 386356 62086 386368
rect 86954 386356 86960 386368
rect 62080 386328 86960 386356
rect 62080 386316 62086 386328
rect 86954 386316 86960 386328
rect 87012 386316 87018 386368
rect 117590 385636 117596 385688
rect 117648 385676 117654 385688
rect 191374 385676 191380 385688
rect 117648 385648 191380 385676
rect 117648 385636 117654 385648
rect 191374 385636 191380 385648
rect 191432 385636 191438 385688
rect 97258 385024 97264 385076
rect 97316 385064 97322 385076
rect 197354 385064 197360 385076
rect 97316 385036 197360 385064
rect 97316 385024 97322 385036
rect 197354 385024 197360 385036
rect 197412 385024 197418 385076
rect 57698 384956 57704 385008
rect 57756 384996 57762 385008
rect 82078 384996 82084 385008
rect 57756 384968 82084 384996
rect 57756 384956 57762 384968
rect 82078 384956 82084 384968
rect 82136 384956 82142 385008
rect 86862 384344 86868 384396
rect 86920 384384 86926 384396
rect 100478 384384 100484 384396
rect 86920 384356 100484 384384
rect 86920 384344 86926 384356
rect 100478 384344 100484 384356
rect 100536 384384 100542 384396
rect 184382 384384 184388 384396
rect 100536 384356 184388 384384
rect 100536 384344 100542 384356
rect 184382 384344 184388 384356
rect 184440 384344 184446 384396
rect 63310 384276 63316 384328
rect 63368 384316 63374 384328
rect 173802 384316 173808 384328
rect 63368 384288 173808 384316
rect 63368 384276 63374 384288
rect 173802 384276 173808 384288
rect 173860 384276 173866 384328
rect 193122 383664 193128 383716
rect 193180 383704 193186 383716
rect 196710 383704 196716 383716
rect 193180 383676 196716 383704
rect 193180 383664 193186 383676
rect 196710 383664 196716 383676
rect 196768 383664 196774 383716
rect 357894 383664 357900 383716
rect 357952 383704 357958 383716
rect 400858 383704 400864 383716
rect 357952 383676 400864 383704
rect 357952 383664 357958 383676
rect 400858 383664 400864 383676
rect 400916 383664 400922 383716
rect 77938 382916 77944 382968
rect 77996 382956 78002 382968
rect 148318 382956 148324 382968
rect 77996 382928 148324 382956
rect 77996 382916 78002 382928
rect 148318 382916 148324 382928
rect 148376 382916 148382 382968
rect 157978 382916 157984 382968
rect 158036 382956 158042 382968
rect 177298 382956 177304 382968
rect 158036 382928 177304 382956
rect 158036 382916 158042 382928
rect 177298 382916 177304 382928
rect 177356 382916 177362 382968
rect 147674 382304 147680 382356
rect 147732 382344 147738 382356
rect 157334 382344 157340 382356
rect 147732 382316 157340 382344
rect 147732 382304 147738 382316
rect 157334 382304 157340 382316
rect 157392 382304 157398 382356
rect 119982 382236 119988 382288
rect 120040 382276 120046 382288
rect 185578 382276 185584 382288
rect 120040 382248 185584 382276
rect 120040 382236 120046 382248
rect 185578 382236 185584 382248
rect 185636 382236 185642 382288
rect 3602 381488 3608 381540
rect 3660 381528 3666 381540
rect 105538 381528 105544 381540
rect 3660 381500 105544 381528
rect 3660 381488 3666 381500
rect 105538 381488 105544 381500
rect 105596 381488 105602 381540
rect 110322 381488 110328 381540
rect 110380 381528 110386 381540
rect 157978 381528 157984 381540
rect 110380 381500 157984 381528
rect 110380 381488 110386 381500
rect 157978 381488 157984 381500
rect 158036 381488 158042 381540
rect 157334 380944 157340 380996
rect 157392 380984 157398 380996
rect 163406 380984 163412 380996
rect 157392 380956 163412 380984
rect 157392 380944 157398 380956
rect 163406 380944 163412 380956
rect 163464 380944 163470 380996
rect 67542 380876 67548 380928
rect 67600 380916 67606 380928
rect 195514 380916 195520 380928
rect 67600 380888 195520 380916
rect 67600 380876 67606 380888
rect 195514 380876 195520 380888
rect 195572 380876 195578 380928
rect 44082 380808 44088 380860
rect 44140 380848 44146 380860
rect 75914 380848 75920 380860
rect 44140 380820 75920 380848
rect 44140 380808 44146 380820
rect 75914 380808 75920 380820
rect 75972 380848 75978 380860
rect 76558 380848 76564 380860
rect 75972 380820 76564 380848
rect 75972 380808 75978 380820
rect 76558 380808 76564 380820
rect 76616 380808 76622 380860
rect 75178 380196 75184 380248
rect 75236 380236 75242 380248
rect 113174 380236 113180 380248
rect 75236 380208 113180 380236
rect 75236 380196 75242 380208
rect 113174 380196 113180 380208
rect 113232 380196 113238 380248
rect 103330 380128 103336 380180
rect 103388 380168 103394 380180
rect 152458 380168 152464 380180
rect 103388 380140 152464 380168
rect 103388 380128 103394 380140
rect 152458 380128 152464 380140
rect 152516 380128 152522 380180
rect 177390 380128 177396 380180
rect 177448 380168 177454 380180
rect 194410 380168 194416 380180
rect 177448 380140 194416 380168
rect 177448 380128 177454 380140
rect 194410 380128 194416 380140
rect 194468 380168 194474 380180
rect 197354 380168 197360 380180
rect 194468 380140 197360 380168
rect 194468 380128 194474 380140
rect 197354 380128 197360 380140
rect 197412 380128 197418 380180
rect 129826 379584 129832 379636
rect 129884 379624 129890 379636
rect 195330 379624 195336 379636
rect 129884 379596 195336 379624
rect 129884 379584 129890 379596
rect 195330 379584 195336 379596
rect 195388 379584 195394 379636
rect 357894 379516 357900 379568
rect 357952 379556 357958 379568
rect 360470 379556 360476 379568
rect 357952 379528 360476 379556
rect 357952 379516 357958 379528
rect 360470 379516 360476 379528
rect 360528 379516 360534 379568
rect 117958 378768 117964 378820
rect 118016 378808 118022 378820
rect 159450 378808 159456 378820
rect 118016 378780 159456 378808
rect 118016 378768 118022 378780
rect 159450 378768 159456 378780
rect 159508 378768 159514 378820
rect 60550 378156 60556 378208
rect 60608 378196 60614 378208
rect 190454 378196 190460 378208
rect 60608 378168 190460 378196
rect 60608 378156 60614 378168
rect 190454 378156 190460 378168
rect 190512 378196 190518 378208
rect 191282 378196 191288 378208
rect 190512 378168 191288 378196
rect 190512 378156 190518 378168
rect 191282 378156 191288 378168
rect 191340 378156 191346 378208
rect 70302 377476 70308 377528
rect 70360 377516 70366 377528
rect 166994 377516 167000 377528
rect 70360 377488 167000 377516
rect 70360 377476 70366 377488
rect 166994 377476 167000 377488
rect 167052 377476 167058 377528
rect 11698 377408 11704 377460
rect 11756 377448 11762 377460
rect 122834 377448 122840 377460
rect 11756 377420 122840 377448
rect 11756 377408 11762 377420
rect 122834 377408 122840 377420
rect 122892 377408 122898 377460
rect 190270 377408 190276 377460
rect 190328 377448 190334 377460
rect 203610 377448 203616 377460
rect 190328 377420 203616 377448
rect 190328 377408 190334 377420
rect 203610 377408 203616 377420
rect 203668 377408 203674 377460
rect 354122 377408 354128 377460
rect 354180 377448 354186 377460
rect 360286 377448 360292 377460
rect 354180 377420 360292 377448
rect 354180 377408 354186 377420
rect 360286 377408 360292 377420
rect 360344 377408 360350 377460
rect 153838 376728 153844 376780
rect 153896 376768 153902 376780
rect 185670 376768 185676 376780
rect 153896 376740 185676 376768
rect 153896 376728 153902 376740
rect 185670 376728 185676 376740
rect 185728 376728 185734 376780
rect 66898 376660 66904 376712
rect 66956 376700 66962 376712
rect 67358 376700 67364 376712
rect 66956 376672 67364 376700
rect 66956 376660 66962 376672
rect 67358 376660 67364 376672
rect 67416 376660 67422 376712
rect 345750 376048 345756 376100
rect 345808 376088 345814 376100
rect 357710 376088 357716 376100
rect 345808 376060 357716 376088
rect 345808 376048 345814 376060
rect 357710 376048 357716 376060
rect 357768 376048 357774 376100
rect 60642 375980 60648 376032
rect 60700 376020 60706 376032
rect 71682 376020 71688 376032
rect 60700 375992 71688 376020
rect 60700 375980 60706 375992
rect 71682 375980 71688 375992
rect 71740 375980 71746 376032
rect 172422 375980 172428 376032
rect 172480 376020 172486 376032
rect 184290 376020 184296 376032
rect 172480 375992 184296 376020
rect 172480 375980 172486 375992
rect 184290 375980 184296 375992
rect 184348 375980 184354 376032
rect 198918 375980 198924 376032
rect 198976 376020 198982 376032
rect 204346 376020 204352 376032
rect 198976 375992 204352 376020
rect 198976 375980 198982 375992
rect 204346 375980 204352 375992
rect 204404 375980 204410 376032
rect 248046 375980 248052 376032
rect 248104 376020 248110 376032
rect 376110 376020 376116 376032
rect 248104 375992 376116 376020
rect 248104 375980 248110 375992
rect 376110 375980 376116 375992
rect 376168 375980 376174 376032
rect 197078 375640 197084 375692
rect 197136 375680 197142 375692
rect 200298 375680 200304 375692
rect 197136 375652 200304 375680
rect 197136 375640 197142 375652
rect 200298 375640 200304 375652
rect 200356 375640 200362 375692
rect 66898 375368 66904 375420
rect 66956 375408 66962 375420
rect 195882 375408 195888 375420
rect 66956 375380 195888 375408
rect 66956 375368 66962 375380
rect 195882 375368 195888 375380
rect 195940 375368 195946 375420
rect 191374 375300 191380 375352
rect 191432 375340 191438 375352
rect 205818 375340 205824 375352
rect 191432 375312 205824 375340
rect 191432 375300 191438 375312
rect 205818 375300 205824 375312
rect 205876 375340 205882 375352
rect 206646 375340 206652 375352
rect 205876 375312 206652 375340
rect 205876 375300 205882 375312
rect 206646 375300 206652 375312
rect 206704 375300 206710 375352
rect 207014 375300 207020 375352
rect 207072 375340 207078 375352
rect 208302 375340 208308 375352
rect 207072 375312 208308 375340
rect 207072 375300 207078 375312
rect 208302 375300 208308 375312
rect 208360 375300 208366 375352
rect 258718 375300 258724 375352
rect 258776 375340 258782 375352
rect 261478 375340 261484 375352
rect 258776 375312 261484 375340
rect 258776 375300 258782 375312
rect 261478 375300 261484 375312
rect 261536 375300 261542 375352
rect 269850 375300 269856 375352
rect 269908 375340 269914 375352
rect 274726 375340 274732 375352
rect 269908 375312 274732 375340
rect 269908 375300 269914 375312
rect 274726 375300 274732 375312
rect 274784 375300 274790 375352
rect 279510 375300 279516 375352
rect 279568 375340 279574 375352
rect 280154 375340 280160 375352
rect 279568 375312 280160 375340
rect 279568 375300 279574 375312
rect 280154 375300 280160 375312
rect 280212 375300 280218 375352
rect 311894 375300 311900 375352
rect 311952 375340 311958 375352
rect 312814 375340 312820 375352
rect 311952 375312 312820 375340
rect 311952 375300 311958 375312
rect 312814 375300 312820 375312
rect 312872 375300 312878 375352
rect 317966 375300 317972 375352
rect 318024 375340 318030 375352
rect 320174 375340 320180 375352
rect 318024 375312 320180 375340
rect 318024 375300 318030 375312
rect 320174 375300 320180 375312
rect 320232 375300 320238 375352
rect 351178 375300 351184 375352
rect 351236 375340 351242 375352
rect 354398 375340 354404 375352
rect 351236 375312 354404 375340
rect 351236 375300 351242 375312
rect 354398 375300 354404 375312
rect 354456 375300 354462 375352
rect 199378 375232 199384 375284
rect 199436 375272 199442 375284
rect 199930 375272 199936 375284
rect 199436 375244 199936 375272
rect 199436 375232 199442 375244
rect 199930 375232 199936 375244
rect 199988 375232 199994 375284
rect 278222 375096 278228 375148
rect 278280 375136 278286 375148
rect 279694 375136 279700 375148
rect 278280 375108 279700 375136
rect 278280 375096 278286 375108
rect 279694 375096 279700 375108
rect 279752 375096 279758 375148
rect 244734 374796 244740 374808
rect 238726 374768 244740 374796
rect 112438 374688 112444 374740
rect 112496 374728 112502 374740
rect 130378 374728 130384 374740
rect 112496 374700 130384 374728
rect 112496 374688 112502 374700
rect 130378 374688 130384 374700
rect 130436 374688 130442 374740
rect 233878 374688 233884 374740
rect 233936 374728 233942 374740
rect 238726 374728 238754 374768
rect 244734 374756 244740 374768
rect 244792 374756 244798 374808
rect 233936 374700 238754 374728
rect 233936 374688 233942 374700
rect 242158 374688 242164 374740
rect 242216 374728 242222 374740
rect 243078 374728 243084 374740
rect 242216 374700 243084 374728
rect 242216 374688 242222 374700
rect 243078 374688 243084 374700
rect 243136 374688 243142 374740
rect 250438 374688 250444 374740
rect 250496 374728 250502 374740
rect 251358 374728 251364 374740
rect 250496 374700 251364 374728
rect 250496 374688 250502 374700
rect 251358 374688 251364 374700
rect 251416 374688 251422 374740
rect 338758 374688 338764 374740
rect 338816 374728 338822 374740
rect 347774 374728 347780 374740
rect 338816 374700 347780 374728
rect 338816 374688 338822 374700
rect 347774 374688 347780 374700
rect 347832 374688 347838 374740
rect 59078 374620 59084 374672
rect 59136 374660 59142 374672
rect 162854 374660 162860 374672
rect 59136 374632 162860 374660
rect 59136 374620 59142 374632
rect 162854 374620 162860 374632
rect 162912 374620 162918 374672
rect 163406 374620 163412 374672
rect 163464 374660 163470 374672
rect 186406 374660 186412 374672
rect 163464 374632 186412 374660
rect 163464 374620 163470 374632
rect 186406 374620 186412 374632
rect 186464 374620 186470 374672
rect 199838 374620 199844 374672
rect 199896 374660 199902 374672
rect 207106 374660 207112 374672
rect 199896 374632 207112 374660
rect 199896 374620 199902 374632
rect 207106 374620 207112 374632
rect 207164 374620 207170 374672
rect 209038 374620 209044 374672
rect 209096 374660 209102 374672
rect 213270 374660 213276 374672
rect 209096 374632 213276 374660
rect 209096 374620 209102 374632
rect 213270 374620 213276 374632
rect 213328 374620 213334 374672
rect 217318 374620 217324 374672
rect 217376 374660 217382 374672
rect 239766 374660 239772 374672
rect 217376 374632 239772 374660
rect 217376 374620 217382 374632
rect 239766 374620 239772 374632
rect 239824 374620 239830 374672
rect 298738 374620 298744 374672
rect 298796 374660 298802 374672
rect 316126 374660 316132 374672
rect 298796 374632 316132 374660
rect 298796 374620 298802 374632
rect 316126 374620 316132 374632
rect 316184 374620 316190 374672
rect 342162 374620 342168 374672
rect 342220 374660 342226 374672
rect 352742 374660 352748 374672
rect 342220 374632 352748 374660
rect 342220 374620 342226 374632
rect 352742 374620 352748 374632
rect 352800 374620 352806 374672
rect 267642 374076 267648 374128
rect 267700 374116 267706 374128
rect 269758 374116 269764 374128
rect 267700 374088 269764 374116
rect 267700 374076 267706 374088
rect 269758 374076 269764 374088
rect 269816 374076 269822 374128
rect 131758 374008 131764 374060
rect 131816 374048 131822 374060
rect 189718 374048 189724 374060
rect 131816 374020 189724 374048
rect 131816 374008 131822 374020
rect 189718 374008 189724 374020
rect 189776 374008 189782 374060
rect 213270 374008 213276 374060
rect 213328 374048 213334 374060
rect 219894 374048 219900 374060
rect 213328 374020 219900 374048
rect 213328 374008 213334 374020
rect 219894 374008 219900 374020
rect 219952 374008 219958 374060
rect 266998 374008 267004 374060
rect 267056 374048 267062 374060
rect 268102 374048 268108 374060
rect 267056 374020 268108 374048
rect 267056 374008 267062 374020
rect 268102 374008 268108 374020
rect 268160 374008 268166 374060
rect 271138 374008 271144 374060
rect 271196 374048 271202 374060
rect 278038 374048 278044 374060
rect 271196 374020 278044 374048
rect 271196 374008 271202 374020
rect 278038 374008 278044 374020
rect 278096 374008 278102 374060
rect 290458 374008 290464 374060
rect 290516 374048 290522 374060
rect 297910 374048 297916 374060
rect 290516 374020 297916 374048
rect 290516 374008 290522 374020
rect 297910 374008 297916 374020
rect 297968 374008 297974 374060
rect 308398 374008 308404 374060
rect 308456 374048 308462 374060
rect 309870 374048 309876 374060
rect 308456 374020 309876 374048
rect 308456 374008 308462 374020
rect 309870 374008 309876 374020
rect 309928 374008 309934 374060
rect 325602 374008 325608 374060
rect 325660 374048 325666 374060
rect 327902 374048 327908 374060
rect 325660 374020 327908 374048
rect 325660 374008 325666 374020
rect 327902 374008 327908 374020
rect 327960 374008 327966 374060
rect 197170 373328 197176 373380
rect 197228 373368 197234 373380
rect 205634 373368 205640 373380
rect 197228 373340 205640 373368
rect 197228 373328 197234 373340
rect 205634 373328 205640 373340
rect 205692 373328 205698 373380
rect 349798 373328 349804 373380
rect 349856 373368 349862 373380
rect 360470 373368 360476 373380
rect 349856 373340 360476 373368
rect 349856 373328 349862 373340
rect 360470 373328 360476 373340
rect 360528 373328 360534 373380
rect 84102 373260 84108 373312
rect 84160 373300 84166 373312
rect 115198 373300 115204 373312
rect 84160 373272 115204 373300
rect 84160 373260 84166 373272
rect 115198 373260 115204 373272
rect 115256 373260 115262 373312
rect 188798 373260 188804 373312
rect 188856 373300 188862 373312
rect 215938 373300 215944 373312
rect 188856 373272 215944 373300
rect 188856 373260 188862 373272
rect 215938 373260 215944 373272
rect 215996 373260 216002 373312
rect 352650 373260 352656 373312
rect 352708 373300 352714 373312
rect 365898 373300 365904 373312
rect 352708 373272 365904 373300
rect 352708 373260 352714 373272
rect 365898 373260 365904 373272
rect 365956 373260 365962 373312
rect 124950 372648 124956 372700
rect 125008 372688 125014 372700
rect 172054 372688 172060 372700
rect 125008 372660 172060 372688
rect 125008 372648 125014 372660
rect 172054 372648 172060 372660
rect 172112 372648 172118 372700
rect 53558 372580 53564 372632
rect 53616 372620 53622 372632
rect 196802 372620 196808 372632
rect 53616 372592 196808 372620
rect 53616 372580 53622 372592
rect 196802 372580 196808 372592
rect 196860 372580 196866 372632
rect 52086 372512 52092 372564
rect 52144 372552 52150 372564
rect 370038 372552 370044 372564
rect 52144 372524 370044 372552
rect 52144 372512 52150 372524
rect 370038 372512 370044 372524
rect 370096 372512 370102 372564
rect 89622 371832 89628 371884
rect 89680 371872 89686 371884
rect 356330 371872 356336 371884
rect 89680 371844 356336 371872
rect 89680 371832 89686 371844
rect 356330 371832 356336 371844
rect 356388 371832 356394 371884
rect 2958 371356 2964 371408
rect 3016 371396 3022 371408
rect 4798 371396 4804 371408
rect 3016 371368 4804 371396
rect 3016 371356 3022 371368
rect 4798 371356 4804 371368
rect 4856 371356 4862 371408
rect 125042 371152 125048 371204
rect 125100 371192 125106 371204
rect 129734 371192 129740 371204
rect 125100 371164 129740 371192
rect 125100 371152 125106 371164
rect 129734 371152 129740 371164
rect 129792 371152 129798 371204
rect 146202 370540 146208 370592
rect 146260 370580 146266 370592
rect 207014 370580 207020 370592
rect 146260 370552 207020 370580
rect 146260 370540 146266 370552
rect 207014 370540 207020 370552
rect 207072 370540 207078 370592
rect 347038 370540 347044 370592
rect 347096 370580 347102 370592
rect 365806 370580 365812 370592
rect 347096 370552 365812 370580
rect 347096 370540 347102 370552
rect 365806 370540 365812 370552
rect 365864 370540 365870 370592
rect 185578 370472 185584 370524
rect 185636 370512 185642 370524
rect 253934 370512 253940 370524
rect 185636 370484 253940 370512
rect 185636 370472 185642 370484
rect 253934 370472 253940 370484
rect 253992 370472 253998 370524
rect 262858 370472 262864 370524
rect 262916 370512 262922 370524
rect 357618 370512 357624 370524
rect 262916 370484 357624 370512
rect 262916 370472 262922 370484
rect 357618 370472 357624 370484
rect 357676 370472 357682 370524
rect 207014 370268 207020 370320
rect 207072 370308 207078 370320
rect 208302 370308 208308 370320
rect 207072 370280 208308 370308
rect 207072 370268 207078 370280
rect 208302 370268 208308 370280
rect 208360 370268 208366 370320
rect 129182 369860 129188 369912
rect 129240 369900 129246 369912
rect 173250 369900 173256 369912
rect 129240 369872 173256 369900
rect 129240 369860 129246 369872
rect 173250 369860 173256 369872
rect 173308 369860 173314 369912
rect 252554 369860 252560 369912
rect 252612 369900 252618 369912
rect 253290 369900 253296 369912
rect 252612 369872 253296 369900
rect 252612 369860 252618 369872
rect 253290 369860 253296 369872
rect 253348 369900 253354 369912
rect 302878 369900 302884 369912
rect 253348 369872 302884 369900
rect 253348 369860 253354 369872
rect 302878 369860 302884 369872
rect 302936 369860 302942 369912
rect 25498 369792 25504 369844
rect 25556 369832 25562 369844
rect 26142 369832 26148 369844
rect 25556 369804 26148 369832
rect 25556 369792 25562 369804
rect 26142 369792 26148 369804
rect 26200 369832 26206 369844
rect 131758 369832 131764 369844
rect 26200 369804 131764 369832
rect 26200 369792 26206 369804
rect 131758 369792 131764 369804
rect 131816 369792 131822 369844
rect 182082 369180 182088 369232
rect 182140 369220 182146 369232
rect 191282 369220 191288 369232
rect 182140 369192 191288 369220
rect 182140 369180 182146 369192
rect 191282 369180 191288 369192
rect 191340 369180 191346 369232
rect 195238 369180 195244 369232
rect 195296 369220 195302 369232
rect 256050 369220 256056 369232
rect 195296 369192 256056 369220
rect 195296 369180 195302 369192
rect 256050 369180 256056 369192
rect 256108 369180 256114 369232
rect 71590 369112 71596 369164
rect 71648 369152 71654 369164
rect 73154 369152 73160 369164
rect 71648 369124 73160 369152
rect 71648 369112 71654 369124
rect 73154 369112 73160 369124
rect 73212 369112 73218 369164
rect 76558 369112 76564 369164
rect 76616 369152 76622 369164
rect 155218 369152 155224 369164
rect 76616 369124 155224 369152
rect 76616 369112 76622 369124
rect 155218 369112 155224 369124
rect 155276 369112 155282 369164
rect 166902 369112 166908 369164
rect 166960 369152 166966 369164
rect 241422 369152 241428 369164
rect 166960 369124 241428 369152
rect 166960 369112 166966 369124
rect 241422 369112 241428 369124
rect 241480 369112 241486 369164
rect 253198 369112 253204 369164
rect 253256 369152 253262 369164
rect 255958 369152 255964 369164
rect 253256 369124 255964 369152
rect 253256 369112 253262 369124
rect 255958 369112 255964 369124
rect 256016 369112 256022 369164
rect 309778 369112 309784 369164
rect 309836 369152 309842 369164
rect 311894 369152 311900 369164
rect 309836 369124 311900 369152
rect 309836 369112 309842 369124
rect 311894 369112 311900 369124
rect 311952 369112 311958 369164
rect 318058 369112 318064 369164
rect 318116 369152 318122 369164
rect 359090 369152 359096 369164
rect 318116 369124 359096 369152
rect 318116 369112 318122 369124
rect 359090 369112 359096 369124
rect 359148 369112 359154 369164
rect 144822 368500 144828 368552
rect 144880 368540 144886 368552
rect 181622 368540 181628 368552
rect 144880 368512 181628 368540
rect 144880 368500 144886 368512
rect 181622 368500 181628 368512
rect 181680 368500 181686 368552
rect 186406 368432 186412 368484
rect 186464 368472 186470 368484
rect 189902 368472 189908 368484
rect 186464 368444 189908 368472
rect 186464 368432 186470 368444
rect 189902 368432 189908 368444
rect 189960 368432 189966 368484
rect 147766 368296 147772 368348
rect 147824 368336 147830 368348
rect 148410 368336 148416 368348
rect 147824 368308 148416 368336
rect 147824 368296 147830 368308
rect 148410 368296 148416 368308
rect 148468 368296 148474 368348
rect 67726 367820 67732 367872
rect 67784 367860 67790 367872
rect 126238 367860 126244 367872
rect 67784 367832 126244 367860
rect 67784 367820 67790 367832
rect 126238 367820 126244 367832
rect 126296 367820 126302 367872
rect 73798 367752 73804 367804
rect 73856 367792 73862 367804
rect 153838 367792 153844 367804
rect 73856 367764 153844 367792
rect 73856 367752 73862 367764
rect 153838 367752 153844 367764
rect 153896 367752 153902 367804
rect 190362 367752 190368 367804
rect 190420 367792 190426 367804
rect 213178 367792 213184 367804
rect 190420 367764 213184 367792
rect 190420 367752 190426 367764
rect 213178 367752 213184 367764
rect 213236 367752 213242 367804
rect 147766 367072 147772 367124
rect 147824 367112 147830 367124
rect 194594 367112 194600 367124
rect 147824 367084 194600 367112
rect 147824 367072 147830 367084
rect 194594 367072 194600 367084
rect 194652 367072 194658 367124
rect 234614 366800 234620 366852
rect 234672 366840 234678 366852
rect 235350 366840 235356 366852
rect 234672 366812 235356 366840
rect 234672 366800 234678 366812
rect 235350 366800 235356 366812
rect 235408 366800 235414 366852
rect 331858 366392 331864 366444
rect 331916 366432 331922 366444
rect 356238 366432 356244 366444
rect 331916 366404 356244 366432
rect 331916 366392 331922 366404
rect 356238 366392 356244 366404
rect 356296 366392 356302 366444
rect 56502 366324 56508 366376
rect 56560 366364 56566 366376
rect 85482 366364 85488 366376
rect 56560 366336 85488 366364
rect 56560 366324 56566 366336
rect 85482 366324 85488 366336
rect 85540 366324 85546 366376
rect 316678 366324 316684 366376
rect 316736 366364 316742 366376
rect 336734 366364 336740 366376
rect 316736 366336 336740 366364
rect 316736 366324 316742 366336
rect 336734 366324 336740 366336
rect 336792 366324 336798 366376
rect 340874 366324 340880 366376
rect 340932 366364 340938 366376
rect 412634 366364 412640 366376
rect 340932 366336 412640 366364
rect 340932 366324 340938 366336
rect 412634 366324 412640 366336
rect 412692 366324 412698 366376
rect 114646 365780 114652 365832
rect 114704 365820 114710 365832
rect 182910 365820 182916 365832
rect 114704 365792 182916 365820
rect 114704 365780 114710 365792
rect 182910 365780 182916 365792
rect 182968 365780 182974 365832
rect 203518 365780 203524 365832
rect 203576 365820 203582 365832
rect 209774 365820 209780 365832
rect 203576 365792 209780 365820
rect 203576 365780 203582 365792
rect 209774 365780 209780 365792
rect 209832 365780 209838 365832
rect 118510 365712 118516 365764
rect 118568 365752 118574 365764
rect 120258 365752 120264 365764
rect 118568 365724 120264 365752
rect 118568 365712 118574 365724
rect 120258 365712 120264 365724
rect 120316 365752 120322 365764
rect 235350 365752 235356 365764
rect 120316 365724 235356 365752
rect 120316 365712 120322 365724
rect 235350 365712 235356 365724
rect 235408 365712 235414 365764
rect 61654 364964 61660 365016
rect 61712 365004 61718 365016
rect 74534 365004 74540 365016
rect 61712 364976 74540 365004
rect 61712 364964 61718 364976
rect 74534 364964 74540 364976
rect 74592 364964 74598 365016
rect 266354 364964 266360 365016
rect 266412 365004 266418 365016
rect 274634 365004 274640 365016
rect 266412 364976 274640 365004
rect 266412 364964 266418 364976
rect 274634 364964 274640 364976
rect 274692 364964 274698 365016
rect 297358 364964 297364 365016
rect 297416 365004 297422 365016
rect 331214 365004 331220 365016
rect 297416 364976 331220 365004
rect 297416 364964 297422 364976
rect 331214 364964 331220 364976
rect 331272 364964 331278 365016
rect 340230 364964 340236 365016
rect 340288 365004 340294 365016
rect 367370 365004 367376 365016
rect 340288 364976 367376 365004
rect 340288 364964 340294 364976
rect 367370 364964 367376 364976
rect 367428 364964 367434 365016
rect 201586 364692 201592 364744
rect 201644 364732 201650 364744
rect 202138 364732 202144 364744
rect 201644 364704 202144 364732
rect 201644 364692 201650 364704
rect 202138 364692 202144 364704
rect 202196 364692 202202 364744
rect 72418 364420 72424 364472
rect 72476 364460 72482 364472
rect 201586 364460 201592 364472
rect 72476 364432 201592 364460
rect 72476 364420 72482 364432
rect 201586 364420 201592 364432
rect 201644 364420 201650 364472
rect 124122 364352 124128 364404
rect 124180 364392 124186 364404
rect 265618 364392 265624 364404
rect 124180 364364 265624 364392
rect 124180 364352 124186 364364
rect 265618 364352 265624 364364
rect 265676 364352 265682 364404
rect 177942 363740 177948 363792
rect 178000 363780 178006 363792
rect 204898 363780 204904 363792
rect 178000 363752 204904 363780
rect 178000 363740 178006 363752
rect 204898 363740 204904 363752
rect 204956 363740 204962 363792
rect 189902 363672 189908 363724
rect 189960 363712 189966 363724
rect 195422 363712 195428 363724
rect 189960 363684 195428 363712
rect 189960 363672 189966 363684
rect 195422 363672 195428 363684
rect 195480 363672 195486 363724
rect 133874 363604 133880 363656
rect 133932 363644 133938 363656
rect 177942 363644 177948 363656
rect 133932 363616 177948 363644
rect 133932 363604 133938 363616
rect 177942 363604 177948 363616
rect 178000 363604 178006 363656
rect 202230 363604 202236 363656
rect 202288 363644 202294 363656
rect 235258 363644 235264 363656
rect 202288 363616 235264 363644
rect 202288 363604 202294 363616
rect 235258 363604 235264 363616
rect 235316 363604 235322 363656
rect 317322 363604 317328 363656
rect 317380 363644 317386 363656
rect 360378 363644 360384 363656
rect 317380 363616 360384 363644
rect 317380 363604 317386 363616
rect 360378 363604 360384 363616
rect 360436 363604 360442 363656
rect 77202 362924 77208 362976
rect 77260 362964 77266 362976
rect 171778 362964 171784 362976
rect 77260 362936 171784 362964
rect 77260 362924 77266 362936
rect 171778 362924 171784 362936
rect 171836 362964 171842 362976
rect 171962 362964 171968 362976
rect 171836 362936 171968 362964
rect 171836 362924 171842 362936
rect 171962 362924 171968 362936
rect 172020 362924 172026 362976
rect 195514 362244 195520 362296
rect 195572 362284 195578 362296
rect 202230 362284 202236 362296
rect 195572 362256 202236 362284
rect 195572 362244 195578 362256
rect 202230 362244 202236 362256
rect 202288 362244 202294 362296
rect 61838 362176 61844 362228
rect 61896 362216 61902 362228
rect 131022 362216 131028 362228
rect 61896 362188 131028 362216
rect 61896 362176 61902 362188
rect 131022 362176 131028 362188
rect 131080 362176 131086 362228
rect 162670 362176 162676 362228
rect 162728 362216 162734 362228
rect 164234 362216 164240 362228
rect 162728 362188 164240 362216
rect 162728 362176 162734 362188
rect 164234 362176 164240 362188
rect 164292 362176 164298 362228
rect 136542 361564 136548 361616
rect 136600 361604 136606 361616
rect 231854 361604 231860 361616
rect 136600 361576 231860 361604
rect 136600 361564 136606 361576
rect 231854 361564 231860 361576
rect 231912 361604 231918 361616
rect 232590 361604 232596 361616
rect 231912 361576 232596 361604
rect 231912 361564 231918 361576
rect 232590 361564 232596 361576
rect 232648 361564 232654 361616
rect 166994 361496 167000 361548
rect 167052 361536 167058 361548
rect 309134 361536 309140 361548
rect 167052 361508 309140 361536
rect 167052 361496 167058 361508
rect 309134 361496 309140 361508
rect 309192 361496 309198 361548
rect 91002 360884 91008 360936
rect 91060 360924 91066 360936
rect 114646 360924 114652 360936
rect 91060 360896 114652 360924
rect 91060 360884 91066 360896
rect 114646 360884 114652 360896
rect 114704 360884 114710 360936
rect 322198 360884 322204 360936
rect 322256 360924 322262 360936
rect 361758 360924 361764 360936
rect 322256 360896 361764 360924
rect 322256 360884 322262 360896
rect 361758 360884 361764 360896
rect 361816 360884 361822 360936
rect 54938 360816 54944 360868
rect 54996 360856 55002 360868
rect 112438 360856 112444 360868
rect 54996 360828 112444 360856
rect 54996 360816 55002 360828
rect 112438 360816 112444 360828
rect 112496 360816 112502 360868
rect 345014 360816 345020 360868
rect 345072 360856 345078 360868
rect 418798 360856 418804 360868
rect 345072 360828 418804 360856
rect 345072 360816 345078 360828
rect 418798 360816 418804 360828
rect 418856 360816 418862 360868
rect 166350 360272 166356 360324
rect 166408 360312 166414 360324
rect 166994 360312 167000 360324
rect 166408 360284 167000 360312
rect 166408 360272 166414 360284
rect 166994 360272 167000 360284
rect 167052 360272 167058 360324
rect 111794 360204 111800 360256
rect 111852 360244 111858 360256
rect 113082 360244 113088 360256
rect 111852 360216 113088 360244
rect 111852 360204 111858 360216
rect 113082 360204 113088 360216
rect 113140 360244 113146 360256
rect 264330 360244 264336 360256
rect 113140 360216 264336 360244
rect 113140 360204 113146 360216
rect 264330 360204 264336 360216
rect 264388 360204 264394 360256
rect 195330 359524 195336 359576
rect 195388 359564 195394 359576
rect 234522 359564 234528 359576
rect 195388 359536 234528 359564
rect 195388 359524 195394 359536
rect 234522 359524 234528 359536
rect 234580 359524 234586 359576
rect 126974 359456 126980 359508
rect 127032 359496 127038 359508
rect 127618 359496 127624 359508
rect 127032 359468 127624 359496
rect 127032 359456 127038 359468
rect 127618 359456 127624 359468
rect 127676 359496 127682 359508
rect 259546 359496 259552 359508
rect 127676 359468 259552 359496
rect 127676 359456 127682 359468
rect 259546 359456 259552 359468
rect 259604 359456 259610 359508
rect 282178 359456 282184 359508
rect 282236 359496 282242 359508
rect 368566 359496 368572 359508
rect 282236 359468 368572 359496
rect 282236 359456 282242 359468
rect 368566 359456 368572 359468
rect 368624 359456 368630 359508
rect 104894 358776 104900 358828
rect 104952 358816 104958 358828
rect 186958 358816 186964 358828
rect 104952 358788 186964 358816
rect 104952 358776 104958 358788
rect 186958 358776 186964 358788
rect 187016 358776 187022 358828
rect 3418 358572 3424 358624
rect 3476 358612 3482 358624
rect 7558 358612 7564 358624
rect 3476 358584 7564 358612
rect 3476 358572 3482 358584
rect 7558 358572 7564 358584
rect 7616 358572 7622 358624
rect 207106 358504 207112 358556
rect 207164 358544 207170 358556
rect 207658 358544 207664 358556
rect 207164 358516 207664 358544
rect 207164 358504 207170 358516
rect 207658 358504 207664 358516
rect 207716 358504 207722 358556
rect 270402 358028 270408 358080
rect 270460 358068 270466 358080
rect 319438 358068 319444 358080
rect 270460 358040 319444 358068
rect 270460 358028 270466 358040
rect 319438 358028 319444 358040
rect 319496 358028 319502 358080
rect 358170 358028 358176 358080
rect 358228 358068 358234 358080
rect 374086 358068 374092 358080
rect 358228 358040 374092 358068
rect 358228 358028 358234 358040
rect 374086 358028 374092 358040
rect 374144 358028 374150 358080
rect 90358 357484 90364 357536
rect 90416 357524 90422 357536
rect 207658 357524 207664 357536
rect 90416 357496 207664 357524
rect 90416 357484 90422 357496
rect 207658 357484 207664 357496
rect 207716 357484 207722 357536
rect 130378 357416 130384 357468
rect 130436 357456 130442 357468
rect 131114 357456 131120 357468
rect 130436 357428 131120 357456
rect 130436 357416 130442 357428
rect 131114 357416 131120 357428
rect 131172 357456 131178 357468
rect 269758 357456 269764 357468
rect 131172 357428 269764 357456
rect 131172 357416 131178 357428
rect 269758 357416 269764 357428
rect 269816 357456 269822 357468
rect 270402 357456 270408 357468
rect 269816 357428 270408 357456
rect 269816 357416 269822 357428
rect 270402 357416 270408 357428
rect 270460 357416 270466 357468
rect 234522 357348 234528 357400
rect 234580 357388 234586 357400
rect 354122 357388 354128 357400
rect 234580 357360 354128 357388
rect 234580 357348 234586 357360
rect 354122 357348 354128 357360
rect 354180 357348 354186 357400
rect 63126 356736 63132 356788
rect 63184 356776 63190 356788
rect 108298 356776 108304 356788
rect 63184 356748 108304 356776
rect 63184 356736 63190 356748
rect 108298 356736 108304 356748
rect 108356 356736 108362 356788
rect 81618 356668 81624 356720
rect 81676 356708 81682 356720
rect 82078 356708 82084 356720
rect 81676 356680 82084 356708
rect 81676 356668 81682 356680
rect 82078 356668 82084 356680
rect 82136 356708 82142 356720
rect 258718 356708 258724 356720
rect 82136 356680 258724 356708
rect 82136 356668 82142 356680
rect 258718 356668 258724 356680
rect 258776 356668 258782 356720
rect 141510 356056 141516 356108
rect 141568 356096 141574 356108
rect 170490 356096 170496 356108
rect 141568 356068 170496 356096
rect 141568 356056 141574 356068
rect 170490 356056 170496 356068
rect 170548 356056 170554 356108
rect 170582 356056 170588 356108
rect 170640 356096 170646 356108
rect 171042 356096 171048 356108
rect 170640 356068 171048 356096
rect 170640 356056 170646 356068
rect 171042 356056 171048 356068
rect 171100 356096 171106 356108
rect 226978 356096 226984 356108
rect 171100 356068 226984 356096
rect 171100 356056 171106 356068
rect 226978 356056 226984 356068
rect 227036 356056 227042 356108
rect 3418 355376 3424 355428
rect 3476 355416 3482 355428
rect 92474 355416 92480 355428
rect 3476 355388 92480 355416
rect 3476 355376 3482 355388
rect 92474 355376 92480 355388
rect 92532 355376 92538 355428
rect 196802 355376 196808 355428
rect 196860 355416 196866 355428
rect 215386 355416 215392 355428
rect 196860 355388 215392 355416
rect 196860 355376 196866 355388
rect 215386 355376 215392 355388
rect 215444 355376 215450 355428
rect 87598 355308 87604 355360
rect 87656 355348 87662 355360
rect 122282 355348 122288 355360
rect 87656 355320 122288 355348
rect 87656 355308 87662 355320
rect 122282 355308 122288 355320
rect 122340 355348 122346 355360
rect 174814 355348 174820 355360
rect 122340 355320 174820 355348
rect 122340 355308 122346 355320
rect 174814 355308 174820 355320
rect 174872 355308 174878 355360
rect 181530 355308 181536 355360
rect 181588 355348 181594 355360
rect 211154 355348 211160 355360
rect 181588 355320 211160 355348
rect 181588 355308 181594 355320
rect 211154 355308 211160 355320
rect 211212 355308 211218 355360
rect 356698 355308 356704 355360
rect 356756 355348 356762 355360
rect 382274 355348 382280 355360
rect 356756 355320 382280 355348
rect 356756 355308 356762 355320
rect 382274 355308 382280 355320
rect 382332 355308 382338 355360
rect 192478 354968 192484 355020
rect 192536 355008 192542 355020
rect 192754 355008 192760 355020
rect 192536 354980 192760 355008
rect 192536 354968 192542 354980
rect 192754 354968 192760 354980
rect 192812 354968 192818 355020
rect 93762 354696 93768 354748
rect 93820 354736 93826 354748
rect 192478 354736 192484 354748
rect 93820 354708 192484 354736
rect 93820 354696 93826 354708
rect 192478 354696 192484 354708
rect 192536 354696 192542 354748
rect 265618 354628 265624 354680
rect 265676 354668 265682 354680
rect 353938 354668 353944 354680
rect 265676 354640 353944 354668
rect 265676 354628 265682 354640
rect 353938 354628 353944 354640
rect 353996 354628 354002 354680
rect 171778 353948 171784 354000
rect 171836 353988 171842 354000
rect 222194 353988 222200 354000
rect 171836 353960 222200 353988
rect 171836 353948 171842 353960
rect 222194 353948 222200 353960
rect 222252 353948 222258 354000
rect 101858 353336 101864 353388
rect 101916 353376 101922 353388
rect 170582 353376 170588 353388
rect 101916 353348 170588 353376
rect 101916 353336 101922 353348
rect 170582 353336 170588 353348
rect 170640 353336 170646 353388
rect 124858 353268 124864 353320
rect 124916 353308 124922 353320
rect 127066 353308 127072 353320
rect 124916 353280 127072 353308
rect 124916 353268 124922 353280
rect 127066 353268 127072 353280
rect 127124 353308 127130 353320
rect 128170 353308 128176 353320
rect 127124 353280 128176 353308
rect 127124 353268 127130 353280
rect 128170 353268 128176 353280
rect 128228 353268 128234 353320
rect 133138 353268 133144 353320
rect 133196 353308 133202 353320
rect 205726 353308 205732 353320
rect 133196 353280 205732 353308
rect 133196 353268 133202 353280
rect 205726 353268 205732 353280
rect 205784 353308 205790 353320
rect 206278 353308 206284 353320
rect 205784 353280 206284 353308
rect 205784 353268 205790 353280
rect 206278 353268 206284 353280
rect 206336 353268 206342 353320
rect 125594 353200 125600 353252
rect 125652 353240 125658 353252
rect 233878 353240 233884 353252
rect 125652 353212 233884 353240
rect 125652 353200 125658 353212
rect 233878 353200 233884 353212
rect 233936 353200 233942 353252
rect 77386 352588 77392 352640
rect 77444 352628 77450 352640
rect 94498 352628 94504 352640
rect 77444 352600 94504 352628
rect 77444 352588 77450 352600
rect 94498 352588 94504 352600
rect 94556 352588 94562 352640
rect 81342 352520 81348 352572
rect 81400 352560 81406 352572
rect 125594 352560 125600 352572
rect 81400 352532 125600 352560
rect 81400 352520 81406 352532
rect 125594 352520 125600 352532
rect 125652 352520 125658 352572
rect 270402 352520 270408 352572
rect 270460 352560 270466 352572
rect 363046 352560 363052 352572
rect 270460 352532 363052 352560
rect 270460 352520 270466 352532
rect 363046 352520 363052 352532
rect 363104 352520 363110 352572
rect 110322 351908 110328 351960
rect 110380 351948 110386 351960
rect 196618 351948 196624 351960
rect 110380 351920 196624 351948
rect 110380 351908 110386 351920
rect 196618 351908 196624 351920
rect 196676 351908 196682 351960
rect 158070 351840 158076 351892
rect 158128 351880 158134 351892
rect 158622 351880 158628 351892
rect 158128 351852 158628 351880
rect 158128 351840 158134 351852
rect 158622 351840 158628 351852
rect 158680 351880 158686 351892
rect 364518 351880 364524 351892
rect 158680 351852 364524 351880
rect 158680 351840 158686 351852
rect 364518 351840 364524 351852
rect 364576 351840 364582 351892
rect 85482 351160 85488 351212
rect 85540 351200 85546 351212
rect 94038 351200 94044 351212
rect 85540 351172 94044 351200
rect 85540 351160 85546 351172
rect 94038 351160 94044 351172
rect 94096 351160 94102 351212
rect 111150 351160 111156 351212
rect 111208 351200 111214 351212
rect 138014 351200 138020 351212
rect 111208 351172 138020 351200
rect 111208 351160 111214 351172
rect 138014 351160 138020 351172
rect 138072 351160 138078 351212
rect 167822 351200 167828 351212
rect 151786 351172 167828 351200
rect 146938 351092 146944 351144
rect 146996 351132 147002 351144
rect 147582 351132 147588 351144
rect 146996 351104 147588 351132
rect 146996 351092 147002 351104
rect 147582 351092 147588 351104
rect 147640 351132 147646 351144
rect 151786 351132 151814 351172
rect 167822 351160 167828 351172
rect 167880 351160 167886 351212
rect 147640 351104 151814 351132
rect 147640 351092 147646 351104
rect 84378 350548 84384 350600
rect 84436 350588 84442 350600
rect 85390 350588 85396 350600
rect 84436 350560 85396 350588
rect 84436 350548 84442 350560
rect 85390 350548 85396 350560
rect 85448 350588 85454 350600
rect 157334 350588 157340 350600
rect 85448 350560 157340 350588
rect 85448 350548 85454 350560
rect 157334 350548 157340 350560
rect 157392 350548 157398 350600
rect 97902 349800 97908 349852
rect 97960 349840 97966 349852
rect 132586 349840 132592 349852
rect 97960 349812 132592 349840
rect 97960 349800 97966 349812
rect 132586 349800 132592 349812
rect 132644 349840 132650 349852
rect 188522 349840 188528 349852
rect 132644 349812 188528 349840
rect 132644 349800 132650 349812
rect 188522 349800 188528 349812
rect 188580 349800 188586 349852
rect 197262 349800 197268 349852
rect 197320 349840 197326 349852
rect 358078 349840 358084 349852
rect 197320 349812 358084 349840
rect 197320 349800 197326 349812
rect 358078 349800 358084 349812
rect 358136 349800 358142 349852
rect 89530 349120 89536 349172
rect 89588 349160 89594 349172
rect 193858 349160 193864 349172
rect 89588 349132 193864 349160
rect 89588 349120 89594 349132
rect 193858 349120 193864 349132
rect 193916 349120 193922 349172
rect 110414 349052 110420 349104
rect 110472 349092 110478 349104
rect 137278 349092 137284 349104
rect 110472 349064 137284 349092
rect 110472 349052 110478 349064
rect 137278 349052 137284 349064
rect 137336 349052 137342 349104
rect 223574 348984 223580 349036
rect 223632 349024 223638 349036
rect 224218 349024 224224 349036
rect 223632 348996 224224 349024
rect 223632 348984 223638 348996
rect 224218 348984 224224 348996
rect 224276 348984 224282 349036
rect 235350 348440 235356 348492
rect 235408 348480 235414 348492
rect 251818 348480 251824 348492
rect 235408 348452 251824 348480
rect 235408 348440 235414 348452
rect 251818 348440 251824 348452
rect 251876 348440 251882 348492
rect 79962 348372 79968 348424
rect 80020 348412 80026 348424
rect 110966 348412 110972 348424
rect 80020 348384 110972 348412
rect 80020 348372 80026 348384
rect 110966 348372 110972 348384
rect 111024 348372 111030 348424
rect 140682 348372 140688 348424
rect 140740 348412 140746 348424
rect 199010 348412 199016 348424
rect 140740 348384 199016 348412
rect 140740 348372 140746 348384
rect 199010 348372 199016 348384
rect 199068 348412 199074 348424
rect 242158 348412 242164 348424
rect 199068 348384 242164 348412
rect 199068 348372 199074 348384
rect 242158 348372 242164 348384
rect 242216 348372 242222 348424
rect 272518 348372 272524 348424
rect 272576 348412 272582 348424
rect 358906 348412 358912 348424
rect 272576 348384 358912 348412
rect 272576 348372 272582 348384
rect 358906 348372 358912 348384
rect 358964 348372 358970 348424
rect 106918 347760 106924 347812
rect 106976 347800 106982 347812
rect 121454 347800 121460 347812
rect 106976 347772 121460 347800
rect 106976 347760 106982 347772
rect 121454 347760 121460 347772
rect 121512 347760 121518 347812
rect 151078 347760 151084 347812
rect 151136 347800 151142 347812
rect 224218 347800 224224 347812
rect 151136 347772 224224 347800
rect 151136 347760 151142 347772
rect 224218 347760 224224 347772
rect 224276 347760 224282 347812
rect 205634 347692 205640 347744
rect 205692 347732 205698 347744
rect 206370 347732 206376 347744
rect 205692 347704 206376 347732
rect 205692 347692 205698 347704
rect 206370 347692 206376 347704
rect 206428 347692 206434 347744
rect 169570 347012 169576 347064
rect 169628 347052 169634 347064
rect 322198 347052 322204 347064
rect 169628 347024 322204 347052
rect 169628 347012 169634 347024
rect 322198 347012 322204 347024
rect 322256 347012 322262 347064
rect 338850 347012 338856 347064
rect 338908 347052 338914 347064
rect 356790 347052 356796 347064
rect 338908 347024 356796 347052
rect 338908 347012 338914 347024
rect 356790 347012 356796 347024
rect 356848 347012 356854 347064
rect 66070 346468 66076 346520
rect 66128 346508 66134 346520
rect 150434 346508 150440 346520
rect 66128 346480 150440 346508
rect 66128 346468 66134 346480
rect 150434 346468 150440 346480
rect 150492 346468 150498 346520
rect 64598 346400 64604 346452
rect 64656 346440 64662 346452
rect 66898 346440 66904 346452
rect 64656 346412 66904 346440
rect 64656 346400 64662 346412
rect 66898 346400 66904 346412
rect 66956 346440 66962 346452
rect 67266 346440 67272 346452
rect 66956 346412 67272 346440
rect 66956 346400 66962 346412
rect 67266 346400 67272 346412
rect 67324 346400 67330 346452
rect 99098 346400 99104 346452
rect 99156 346440 99162 346452
rect 206370 346440 206376 346452
rect 99156 346412 206376 346440
rect 99156 346400 99162 346412
rect 206370 346400 206376 346412
rect 206428 346400 206434 346452
rect 157334 346332 157340 346384
rect 157392 346372 157398 346384
rect 181530 346372 181536 346384
rect 157392 346344 181536 346372
rect 157392 346332 157398 346344
rect 181530 346332 181536 346344
rect 181588 346332 181594 346384
rect 350442 346332 350448 346384
rect 350500 346372 350506 346384
rect 352558 346372 352564 346384
rect 350500 346344 352564 346372
rect 350500 346332 350506 346344
rect 352558 346332 352564 346344
rect 352616 346332 352622 346384
rect 99282 345652 99288 345704
rect 99340 345692 99346 345704
rect 158070 345692 158076 345704
rect 99340 345664 158076 345692
rect 99340 345652 99346 345664
rect 158070 345652 158076 345664
rect 158128 345652 158134 345704
rect 189718 345652 189724 345704
rect 189776 345692 189782 345704
rect 209774 345692 209780 345704
rect 189776 345664 209780 345692
rect 189776 345652 189782 345664
rect 209774 345652 209780 345664
rect 209832 345652 209838 345704
rect 249058 345652 249064 345704
rect 249116 345692 249122 345704
rect 269850 345692 269856 345704
rect 249116 345664 269856 345692
rect 249116 345652 249122 345664
rect 269850 345652 269856 345664
rect 269908 345652 269914 345704
rect 122834 345040 122840 345092
rect 122892 345080 122898 345092
rect 123478 345080 123484 345092
rect 122892 345052 123484 345080
rect 122892 345040 122898 345052
rect 123478 345040 123484 345052
rect 123536 345080 123542 345092
rect 249058 345080 249064 345092
rect 123536 345052 249064 345080
rect 123536 345040 123542 345052
rect 249058 345040 249064 345052
rect 249116 345040 249122 345092
rect 150434 344972 150440 345024
rect 150492 345012 150498 345024
rect 197998 345012 198004 345024
rect 150492 344984 198004 345012
rect 150492 344972 150498 344984
rect 197998 344972 198004 344984
rect 198056 344972 198062 345024
rect 286226 344292 286232 344344
rect 286284 344332 286290 344344
rect 420914 344332 420920 344344
rect 286284 344304 420920 344332
rect 286284 344292 286290 344304
rect 420914 344292 420920 344304
rect 420972 344292 420978 344344
rect 115842 343612 115848 343664
rect 115900 343652 115906 343664
rect 125042 343652 125048 343664
rect 115900 343624 125048 343652
rect 115900 343612 115906 343624
rect 125042 343612 125048 343624
rect 125100 343612 125106 343664
rect 137278 343612 137284 343664
rect 137336 343652 137342 343664
rect 156782 343652 156788 343664
rect 137336 343624 156788 343652
rect 137336 343612 137342 343624
rect 156782 343612 156788 343624
rect 156840 343612 156846 343664
rect 157978 343612 157984 343664
rect 158036 343652 158042 343664
rect 159542 343652 159548 343664
rect 158036 343624 159548 343652
rect 158036 343612 158042 343624
rect 159542 343612 159548 343624
rect 159600 343612 159606 343664
rect 186222 343612 186228 343664
rect 186280 343652 186286 343664
rect 190454 343652 190460 343664
rect 186280 343624 190460 343652
rect 186280 343612 186286 343624
rect 190454 343612 190460 343624
rect 190512 343612 190518 343664
rect 264330 343544 264336 343596
rect 264388 343584 264394 343596
rect 343634 343584 343640 343596
rect 264388 343556 343640 343584
rect 264388 343544 264394 343556
rect 343634 343544 343640 343556
rect 343692 343544 343698 343596
rect 71682 342932 71688 342984
rect 71740 342972 71746 342984
rect 87138 342972 87144 342984
rect 71740 342944 87144 342972
rect 71740 342932 71746 342944
rect 87138 342932 87144 342944
rect 87196 342932 87202 342984
rect 96430 342932 96436 342984
rect 96488 342972 96494 342984
rect 111150 342972 111156 342984
rect 96488 342944 111156 342972
rect 96488 342932 96494 342944
rect 111150 342932 111156 342944
rect 111208 342932 111214 342984
rect 60366 342864 60372 342916
rect 60424 342904 60430 342916
rect 97258 342904 97264 342916
rect 60424 342876 97264 342904
rect 60424 342864 60430 342876
rect 97258 342864 97264 342876
rect 97316 342864 97322 342916
rect 195514 342864 195520 342916
rect 195572 342904 195578 342916
rect 261478 342904 261484 342916
rect 195572 342876 261484 342904
rect 195572 342864 195578 342876
rect 261478 342864 261484 342876
rect 261536 342864 261542 342916
rect 264330 342796 264336 342848
rect 264388 342836 264394 342848
rect 264882 342836 264888 342848
rect 264388 342808 264888 342836
rect 264388 342796 264394 342808
rect 264882 342796 264888 342808
rect 264940 342796 264946 342848
rect 115750 342320 115756 342372
rect 115808 342360 115814 342372
rect 183186 342360 183192 342372
rect 115808 342332 183192 342360
rect 115808 342320 115814 342332
rect 183186 342320 183192 342332
rect 183244 342320 183250 342372
rect 111702 342252 111708 342304
rect 111760 342292 111766 342304
rect 115842 342292 115848 342304
rect 111760 342264 115848 342292
rect 111760 342252 111766 342264
rect 115842 342252 115848 342264
rect 115900 342252 115906 342304
rect 144178 342252 144184 342304
rect 144236 342292 144242 342304
rect 220078 342292 220084 342304
rect 144236 342264 220084 342292
rect 144236 342252 144242 342264
rect 220078 342252 220084 342264
rect 220136 342252 220142 342304
rect 69750 341504 69756 341556
rect 69808 341544 69814 341556
rect 141510 341544 141516 341556
rect 69808 341516 141516 341544
rect 69808 341504 69814 341516
rect 141510 341504 141516 341516
rect 141568 341504 141574 341556
rect 153838 341504 153844 341556
rect 153896 341544 153902 341556
rect 163590 341544 163596 341556
rect 153896 341516 163596 341544
rect 153896 341504 153902 341516
rect 163590 341504 163596 341516
rect 163648 341504 163654 341556
rect 188430 341504 188436 341556
rect 188488 341544 188494 341556
rect 211798 341544 211804 341556
rect 188488 341516 211804 341544
rect 188488 341504 188494 341516
rect 211798 341504 211804 341516
rect 211856 341504 211862 341556
rect 142338 340960 142344 341012
rect 142396 341000 142402 341012
rect 154022 341000 154028 341012
rect 142396 340972 154028 341000
rect 142396 340960 142402 340972
rect 154022 340960 154028 340972
rect 154080 340960 154086 341012
rect 85574 340892 85580 340944
rect 85632 340932 85638 340944
rect 252554 340932 252560 340944
rect 85632 340904 252560 340932
rect 85632 340892 85638 340904
rect 252554 340892 252560 340904
rect 252612 340892 252618 340944
rect 251910 340824 251916 340876
rect 251968 340864 251974 340876
rect 259086 340864 259092 340876
rect 251968 340836 259092 340864
rect 251968 340824 251974 340836
rect 259086 340824 259092 340836
rect 259144 340824 259150 340876
rect 53650 340144 53656 340196
rect 53708 340184 53714 340196
rect 86954 340184 86960 340196
rect 53708 340156 86960 340184
rect 53708 340144 53714 340156
rect 86954 340144 86960 340156
rect 87012 340144 87018 340196
rect 107470 340144 107476 340196
rect 107528 340184 107534 340196
rect 133138 340184 133144 340196
rect 107528 340156 133144 340184
rect 107528 340144 107534 340156
rect 133138 340144 133144 340156
rect 133196 340144 133202 340196
rect 224218 340144 224224 340196
rect 224276 340184 224282 340196
rect 243538 340184 243544 340196
rect 224276 340156 243544 340184
rect 224276 340144 224282 340156
rect 243538 340144 243544 340156
rect 243596 340144 243602 340196
rect 258810 340144 258816 340196
rect 258868 340184 258874 340196
rect 259086 340184 259092 340196
rect 258868 340156 259092 340184
rect 258868 340144 258874 340156
rect 259086 340144 259092 340156
rect 259144 340184 259150 340196
rect 349154 340184 349160 340196
rect 259144 340156 349160 340184
rect 259144 340144 259150 340156
rect 349154 340144 349160 340156
rect 349212 340144 349218 340196
rect 134242 339532 134248 339584
rect 134300 339572 134306 339584
rect 213270 339572 213276 339584
rect 134300 339544 213276 339572
rect 134300 339532 134306 339544
rect 213270 339532 213276 339544
rect 213328 339532 213334 339584
rect 67818 339464 67824 339516
rect 67876 339504 67882 339516
rect 229738 339504 229744 339516
rect 67876 339476 229744 339504
rect 67876 339464 67882 339476
rect 229738 339464 229744 339476
rect 229796 339464 229802 339516
rect 237926 339396 237932 339448
rect 237984 339436 237990 339448
rect 240134 339436 240140 339448
rect 237984 339408 240140 339436
rect 237984 339396 237990 339408
rect 240134 339396 240140 339408
rect 240192 339396 240198 339448
rect 84102 338716 84108 338768
rect 84160 338756 84166 338768
rect 104158 338756 104164 338768
rect 84160 338728 104164 338756
rect 84160 338716 84166 338728
rect 104158 338716 104164 338728
rect 104216 338716 104222 338768
rect 283558 338716 283564 338768
rect 283616 338756 283622 338768
rect 379514 338756 379520 338768
rect 283616 338728 379520 338756
rect 283616 338716 283622 338728
rect 379514 338716 379520 338728
rect 379572 338716 379578 338768
rect 100570 338172 100576 338224
rect 100628 338212 100634 338224
rect 154482 338212 154488 338224
rect 100628 338184 154488 338212
rect 100628 338172 100634 338184
rect 154482 338172 154488 338184
rect 154540 338172 154546 338224
rect 155310 338172 155316 338224
rect 155368 338212 155374 338224
rect 237926 338212 237932 338224
rect 155368 338184 237932 338212
rect 155368 338172 155374 338184
rect 237926 338172 237932 338184
rect 237984 338212 237990 338224
rect 238662 338212 238668 338224
rect 237984 338184 238668 338212
rect 237984 338172 237990 338184
rect 238662 338172 238668 338184
rect 238720 338172 238726 338224
rect 103698 338104 103704 338156
rect 103756 338144 103762 338156
rect 252646 338144 252652 338156
rect 103756 338116 252652 338144
rect 103756 338104 103762 338116
rect 252646 338104 252652 338116
rect 252704 338104 252710 338156
rect 151078 338036 151084 338088
rect 151136 338076 151142 338088
rect 152642 338076 152648 338088
rect 151136 338048 152648 338076
rect 151136 338036 151142 338048
rect 152642 338036 152648 338048
rect 152700 338036 152706 338088
rect 176102 337560 176108 337612
rect 176160 337600 176166 337612
rect 183002 337600 183008 337612
rect 176160 337572 183008 337600
rect 176160 337560 176166 337572
rect 183002 337560 183008 337572
rect 183060 337560 183066 337612
rect 209130 337424 209136 337476
rect 209188 337464 209194 337476
rect 264974 337464 264980 337476
rect 209188 337436 264980 337464
rect 209188 337424 209194 337436
rect 264974 337424 264980 337436
rect 265032 337424 265038 337476
rect 183094 337356 183100 337408
rect 183152 337396 183158 337408
rect 202874 337396 202880 337408
rect 183152 337368 202880 337396
rect 183152 337356 183158 337368
rect 202874 337356 202880 337368
rect 202932 337356 202938 337408
rect 245010 337356 245016 337408
rect 245068 337396 245074 337408
rect 367278 337396 367284 337408
rect 245068 337368 367284 337396
rect 245068 337356 245074 337368
rect 367278 337356 367284 337368
rect 367336 337356 367342 337408
rect 114462 336812 114468 336864
rect 114520 336852 114526 336864
rect 174538 336852 174544 336864
rect 114520 336824 174544 336852
rect 114520 336812 114526 336824
rect 174538 336812 174544 336824
rect 174596 336812 174602 336864
rect 64690 336744 64696 336796
rect 64748 336784 64754 336796
rect 224218 336784 224224 336796
rect 64748 336756 224224 336784
rect 64748 336744 64754 336756
rect 224218 336744 224224 336756
rect 224276 336744 224282 336796
rect 67726 336676 67732 336728
rect 67784 336716 67790 336728
rect 71774 336716 71780 336728
rect 67784 336688 71780 336716
rect 67784 336676 67790 336688
rect 71774 336676 71780 336688
rect 71832 336676 71838 336728
rect 76650 336064 76656 336116
rect 76708 336104 76714 336116
rect 87598 336104 87604 336116
rect 76708 336076 87604 336104
rect 76708 336064 76714 336076
rect 87598 336064 87604 336076
rect 87656 336064 87662 336116
rect 81066 335996 81072 336048
rect 81124 336036 81130 336048
rect 93118 336036 93124 336048
rect 81124 336008 93124 336036
rect 81124 335996 81130 336008
rect 93118 335996 93124 336008
rect 93176 335996 93182 336048
rect 150526 335996 150532 336048
rect 150584 336036 150590 336048
rect 199470 336036 199476 336048
rect 150584 336008 199476 336036
rect 150584 335996 150590 336008
rect 199470 335996 199476 336008
rect 199528 335996 199534 336048
rect 113082 335384 113088 335436
rect 113140 335424 113146 335436
rect 150434 335424 150440 335436
rect 113140 335396 150440 335424
rect 113140 335384 113146 335396
rect 150434 335384 150440 335396
rect 150492 335384 150498 335436
rect 94130 335316 94136 335368
rect 94188 335356 94194 335368
rect 248506 335356 248512 335368
rect 94188 335328 248512 335356
rect 94188 335316 94194 335328
rect 248506 335316 248512 335328
rect 248564 335316 248570 335368
rect 125042 335248 125048 335300
rect 125100 335288 125106 335300
rect 144178 335288 144184 335300
rect 125100 335260 144184 335288
rect 125100 335248 125106 335260
rect 144178 335248 144184 335260
rect 144236 335248 144242 335300
rect 251910 334636 251916 334688
rect 251968 334676 251974 334688
rect 348418 334676 348424 334688
rect 251968 334648 348424 334676
rect 251968 334636 251974 334648
rect 348418 334636 348424 334648
rect 348476 334636 348482 334688
rect 64506 334568 64512 334620
rect 64564 334608 64570 334620
rect 106918 334608 106924 334620
rect 64564 334580 106924 334608
rect 64564 334568 64570 334580
rect 106918 334568 106924 334580
rect 106976 334568 106982 334620
rect 188430 334568 188436 334620
rect 188488 334608 188494 334620
rect 313274 334608 313280 334620
rect 188488 334580 313280 334608
rect 188488 334568 188494 334580
rect 313274 334568 313280 334580
rect 313332 334568 313338 334620
rect 52178 334024 52184 334076
rect 52236 334064 52242 334076
rect 125502 334064 125508 334076
rect 52236 334036 125508 334064
rect 52236 334024 52242 334036
rect 125502 334024 125508 334036
rect 125560 334024 125566 334076
rect 145282 334024 145288 334076
rect 145340 334064 145346 334076
rect 163314 334064 163320 334076
rect 145340 334036 163320 334064
rect 145340 334024 145346 334036
rect 163314 334024 163320 334036
rect 163372 334024 163378 334076
rect 116762 333956 116768 334008
rect 116820 333996 116826 334008
rect 192662 333996 192668 334008
rect 116820 333968 192668 333996
rect 116820 333956 116826 333968
rect 192662 333956 192668 333968
rect 192720 333956 192726 334008
rect 66162 333208 66168 333260
rect 66220 333248 66226 333260
rect 124214 333248 124220 333260
rect 66220 333220 124220 333248
rect 66220 333208 66226 333220
rect 124214 333208 124220 333220
rect 124272 333208 124278 333260
rect 150434 333208 150440 333260
rect 150492 333248 150498 333260
rect 228358 333248 228364 333260
rect 150492 333220 228364 333248
rect 150492 333208 150498 333220
rect 228358 333208 228364 333220
rect 228416 333208 228422 333260
rect 60458 332596 60464 332648
rect 60516 332636 60522 332648
rect 140774 332636 140780 332648
rect 60516 332608 140780 332636
rect 60516 332596 60522 332608
rect 140774 332596 140780 332608
rect 140832 332596 140838 332648
rect 150342 332596 150348 332648
rect 150400 332636 150406 332648
rect 159358 332636 159364 332648
rect 150400 332608 159364 332636
rect 150400 332596 150406 332608
rect 159358 332596 159364 332608
rect 159416 332596 159422 332648
rect 198826 332528 198832 332580
rect 198884 332568 198890 332580
rect 202322 332568 202328 332580
rect 198884 332540 202328 332568
rect 198884 332528 198890 332540
rect 202322 332528 202328 332540
rect 202380 332528 202386 332580
rect 202782 332528 202788 332580
rect 202840 332568 202846 332580
rect 335354 332568 335360 332580
rect 202840 332540 335360 332568
rect 202840 332528 202846 332540
rect 335354 332528 335360 332540
rect 335412 332528 335418 332580
rect 202230 332324 202236 332376
rect 202288 332364 202294 332376
rect 202782 332364 202788 332376
rect 202288 332336 202788 332364
rect 202288 332324 202294 332336
rect 202782 332324 202788 332336
rect 202840 332324 202846 332376
rect 72970 332120 72976 332172
rect 73028 332160 73034 332172
rect 73798 332160 73804 332172
rect 73028 332132 73804 332160
rect 73028 332120 73034 332132
rect 73798 332120 73804 332132
rect 73856 332120 73862 332172
rect 75822 332120 75828 332172
rect 75880 332160 75886 332172
rect 76558 332160 76564 332172
rect 75880 332132 76564 332160
rect 75880 332120 75886 332132
rect 76558 332120 76564 332132
rect 76616 332120 76622 332172
rect 90450 332120 90456 332172
rect 90508 332160 90514 332172
rect 90910 332160 90916 332172
rect 90508 332132 90916 332160
rect 90508 332120 90514 332132
rect 90910 332120 90916 332132
rect 90968 332120 90974 332172
rect 91830 332120 91836 332172
rect 91888 332160 91894 332172
rect 93210 332160 93216 332172
rect 91888 332132 93216 332160
rect 91888 332120 91894 332132
rect 93210 332120 93216 332132
rect 93268 332120 93274 332172
rect 100018 332120 100024 332172
rect 100076 332160 100082 332172
rect 100570 332160 100576 332172
rect 100076 332132 100576 332160
rect 100076 332120 100082 332132
rect 100570 332120 100576 332132
rect 100628 332120 100634 332172
rect 110874 332120 110880 332172
rect 110932 332160 110938 332172
rect 111610 332160 111616 332172
rect 110932 332132 111616 332160
rect 110932 332120 110938 332132
rect 111610 332120 111616 332132
rect 111668 332120 111674 332172
rect 118878 331984 118884 332036
rect 118936 332024 118942 332036
rect 119890 332024 119896 332036
rect 118936 331996 119896 332024
rect 118936 331984 118942 331996
rect 119890 331984 119896 331996
rect 119948 331984 119954 332036
rect 129274 331916 129280 331968
rect 129332 331956 129338 331968
rect 145282 331956 145288 331968
rect 129332 331928 145288 331956
rect 129332 331916 129338 331928
rect 145282 331916 145288 331928
rect 145340 331916 145346 331968
rect 167822 331916 167828 331968
rect 167880 331956 167886 331968
rect 191098 331956 191104 331968
rect 167880 331928 191104 331956
rect 167880 331916 167886 331928
rect 191098 331916 191104 331928
rect 191156 331916 191162 331968
rect 103238 331848 103244 331900
rect 103296 331888 103302 331900
rect 129090 331888 129096 331900
rect 103296 331860 129096 331888
rect 103296 331848 103302 331860
rect 129090 331848 129096 331860
rect 129148 331848 129154 331900
rect 140774 331848 140780 331900
rect 140832 331888 140838 331900
rect 157334 331888 157340 331900
rect 140832 331860 157340 331888
rect 140832 331848 140838 331860
rect 157334 331848 157340 331860
rect 157392 331848 157398 331900
rect 187234 331848 187240 331900
rect 187292 331888 187298 331900
rect 249794 331888 249800 331900
rect 187292 331860 249800 331888
rect 187292 331848 187298 331860
rect 249794 331848 249800 331860
rect 249852 331848 249858 331900
rect 70670 331780 70676 331832
rect 70728 331820 70734 331832
rect 72418 331820 72424 331832
rect 70728 331792 72424 331820
rect 70728 331780 70734 331792
rect 72418 331780 72424 331792
rect 72476 331780 72482 331832
rect 77662 331780 77668 331832
rect 77720 331820 77726 331832
rect 77938 331820 77944 331832
rect 77720 331792 77944 331820
rect 77720 331780 77726 331792
rect 77938 331780 77944 331792
rect 77996 331780 78002 331832
rect 97074 331712 97080 331764
rect 97132 331752 97138 331764
rect 97902 331752 97908 331764
rect 97132 331724 97908 331752
rect 97132 331712 97138 331724
rect 97902 331712 97908 331724
rect 97960 331712 97966 331764
rect 88242 331576 88248 331628
rect 88300 331616 88306 331628
rect 90358 331616 90364 331628
rect 88300 331588 90364 331616
rect 88300 331576 88306 331588
rect 90358 331576 90364 331588
rect 90416 331576 90422 331628
rect 80330 331508 80336 331560
rect 80388 331548 80394 331560
rect 81342 331548 81348 331560
rect 80388 331520 81348 331548
rect 80388 331508 80394 331520
rect 81342 331508 81348 331520
rect 81400 331508 81406 331560
rect 95602 331508 95608 331560
rect 95660 331548 95666 331560
rect 96522 331548 96528 331560
rect 95660 331520 96528 331548
rect 95660 331508 95666 331520
rect 96522 331508 96528 331520
rect 96580 331508 96586 331560
rect 88978 331440 88984 331492
rect 89036 331480 89042 331492
rect 89622 331480 89628 331492
rect 89036 331452 89628 331480
rect 89036 331440 89042 331452
rect 89622 331440 89628 331452
rect 89680 331440 89686 331492
rect 98546 331440 98552 331492
rect 98604 331480 98610 331492
rect 99190 331480 99196 331492
rect 98604 331452 99196 331480
rect 98604 331440 98610 331452
rect 99190 331440 99196 331452
rect 99248 331440 99254 331492
rect 123294 331440 123300 331492
rect 123352 331480 123358 331492
rect 124122 331480 124128 331492
rect 123352 331452 124128 331480
rect 123352 331440 123358 331452
rect 124122 331440 124128 331452
rect 124180 331440 124186 331492
rect 129918 331440 129924 331492
rect 129976 331480 129982 331492
rect 130378 331480 130384 331492
rect 129976 331452 130384 331480
rect 129976 331440 129982 331452
rect 130378 331440 130384 331452
rect 130436 331440 130442 331492
rect 131482 331440 131488 331492
rect 131540 331480 131546 331492
rect 132402 331480 132408 331492
rect 131540 331452 132408 331480
rect 131540 331440 131546 331452
rect 132402 331440 132408 331452
rect 132460 331440 132466 331492
rect 132770 331440 132776 331492
rect 132828 331480 132834 331492
rect 133690 331480 133696 331492
rect 132828 331452 133696 331480
rect 132828 331440 132834 331452
rect 133690 331440 133696 331452
rect 133748 331440 133754 331492
rect 135714 331440 135720 331492
rect 135772 331480 135778 331492
rect 141418 331480 141424 331492
rect 135772 331452 141424 331480
rect 135772 331440 135778 331452
rect 141418 331440 141424 331452
rect 141476 331440 141482 331492
rect 50982 331304 50988 331356
rect 51040 331344 51046 331356
rect 69382 331344 69388 331356
rect 51040 331316 69388 331344
rect 51040 331304 51046 331316
rect 69382 331304 69388 331316
rect 69440 331304 69446 331356
rect 109402 331304 109408 331356
rect 109460 331344 109466 331356
rect 110322 331344 110328 331356
rect 109460 331316 110328 331344
rect 109460 331304 109466 331316
rect 110322 331304 110328 331316
rect 110380 331304 110386 331356
rect 138658 331304 138664 331356
rect 138716 331344 138722 331356
rect 139302 331344 139308 331356
rect 138716 331316 139308 331344
rect 138716 331304 138722 331316
rect 139302 331304 139308 331316
rect 139360 331304 139366 331356
rect 143810 331304 143816 331356
rect 143868 331344 143874 331356
rect 144822 331344 144828 331356
rect 143868 331316 144828 331344
rect 143868 331304 143874 331316
rect 144822 331304 144828 331316
rect 144880 331304 144886 331356
rect 52270 331236 52276 331288
rect 52328 331276 52334 331288
rect 77662 331276 77668 331288
rect 52328 331248 77668 331276
rect 52328 331236 52334 331248
rect 77662 331236 77668 331248
rect 77720 331236 77726 331288
rect 126882 331236 126888 331288
rect 126940 331276 126946 331288
rect 129734 331276 129740 331288
rect 126940 331248 129740 331276
rect 126940 331236 126946 331248
rect 129734 331236 129740 331248
rect 129792 331236 129798 331288
rect 146754 331236 146760 331288
rect 146812 331276 146818 331288
rect 176102 331276 176108 331288
rect 146812 331248 176108 331276
rect 146812 331236 146818 331248
rect 176102 331236 176108 331248
rect 176160 331236 176166 331288
rect 195422 331236 195428 331288
rect 195480 331276 195486 331288
rect 198734 331276 198740 331288
rect 195480 331248 198740 331276
rect 195480 331236 195486 331248
rect 198734 331236 198740 331248
rect 198792 331236 198798 331288
rect 50522 331168 50528 331220
rect 50580 331208 50586 331220
rect 50798 331208 50804 331220
rect 50580 331180 50804 331208
rect 50580 331168 50586 331180
rect 50798 331168 50804 331180
rect 50856 331208 50862 331220
rect 136542 331208 136548 331220
rect 50856 331180 136548 331208
rect 50856 331168 50862 331180
rect 136542 331168 136548 331180
rect 136600 331168 136606 331220
rect 153194 330556 153200 330608
rect 153252 330596 153258 330608
rect 155954 330596 155960 330608
rect 153252 330568 155960 330596
rect 153252 330556 153258 330568
rect 155954 330556 155960 330568
rect 156012 330556 156018 330608
rect 157334 330556 157340 330608
rect 157392 330596 157398 330608
rect 167914 330596 167920 330608
rect 157392 330568 167920 330596
rect 157392 330556 157398 330568
rect 167914 330556 167920 330568
rect 167972 330556 167978 330608
rect 33778 330488 33784 330540
rect 33836 330528 33842 330540
rect 50522 330528 50528 330540
rect 33836 330500 50528 330528
rect 33836 330488 33842 330500
rect 50522 330488 50528 330500
rect 50580 330488 50586 330540
rect 125502 330488 125508 330540
rect 125560 330528 125566 330540
rect 125560 330500 138014 330528
rect 125560 330488 125566 330500
rect 137986 330460 138014 330500
rect 159450 330488 159456 330540
rect 159508 330528 159514 330540
rect 160094 330528 160100 330540
rect 159508 330500 160100 330528
rect 159508 330488 159514 330500
rect 160094 330488 160100 330500
rect 160152 330488 160158 330540
rect 162118 330488 162124 330540
rect 162176 330528 162182 330540
rect 225598 330528 225604 330540
rect 162176 330500 225604 330528
rect 162176 330488 162182 330500
rect 225598 330488 225604 330500
rect 225656 330488 225662 330540
rect 153194 330460 153200 330472
rect 137986 330432 153200 330460
rect 153194 330420 153200 330432
rect 153252 330420 153258 330472
rect 151170 329808 151176 329860
rect 151228 329848 151234 329860
rect 157978 329848 157984 329860
rect 151228 329820 157984 329848
rect 151228 329808 151234 329820
rect 157978 329808 157984 329820
rect 158036 329808 158042 329860
rect 70026 329740 70032 329792
rect 70084 329780 70090 329792
rect 71038 329780 71044 329792
rect 70084 329752 71044 329780
rect 70084 329740 70090 329752
rect 71038 329740 71044 329752
rect 71096 329740 71102 329792
rect 153194 329740 153200 329792
rect 153252 329780 153258 329792
rect 198090 329780 198096 329792
rect 153252 329752 198096 329780
rect 153252 329740 153258 329752
rect 198090 329740 198096 329752
rect 198148 329740 198154 329792
rect 67266 329672 67272 329724
rect 67324 329712 67330 329724
rect 69750 329712 69756 329724
rect 67324 329684 69756 329712
rect 67324 329672 67330 329684
rect 69750 329672 69756 329684
rect 69808 329672 69814 329724
rect 144886 329140 154574 329168
rect 94222 329100 94228 329112
rect 84166 329072 94228 329100
rect 14 328448 20 328500
rect 72 328488 78 328500
rect 84166 328488 84194 329072
rect 94222 329060 94228 329072
rect 94280 329060 94286 329112
rect 115382 329060 115388 329112
rect 115440 329060 115446 329112
rect 132218 329060 132224 329112
rect 132276 329100 132282 329112
rect 132276 329072 132494 329100
rect 132276 329060 132282 329072
rect 72 328460 72924 328488
rect 72 328448 78 328460
rect 72896 328420 72924 328460
rect 73080 328460 84194 328488
rect 73080 328420 73108 328460
rect 115400 328420 115428 329060
rect 132466 328488 132494 329072
rect 144886 328624 144914 329140
rect 145374 329060 145380 329112
rect 145432 329060 145438 329112
rect 152182 329060 152188 329112
rect 152240 329060 152246 329112
rect 137986 328596 144914 328624
rect 137986 328488 138014 328596
rect 132466 328460 138014 328488
rect 145392 328488 145420 329060
rect 152200 328896 152228 329060
rect 152200 328868 152320 328896
rect 152292 328556 152320 328868
rect 154546 328624 154574 329140
rect 155862 329060 155868 329112
rect 155920 329060 155926 329112
rect 156322 329060 156328 329112
rect 156380 329100 156386 329112
rect 157058 329100 157064 329112
rect 156380 329072 157064 329100
rect 156380 329060 156386 329072
rect 157058 329060 157064 329072
rect 157116 329060 157122 329112
rect 164786 329060 164792 329112
rect 164844 329100 164850 329112
rect 182174 329100 182180 329112
rect 164844 329072 182180 329100
rect 164844 329060 164850 329072
rect 182174 329060 182180 329072
rect 182232 329060 182238 329112
rect 186958 329060 186964 329112
rect 187016 329100 187022 329112
rect 220170 329100 220176 329112
rect 187016 329072 220176 329100
rect 187016 329060 187022 329072
rect 220170 329060 220176 329072
rect 220228 329060 220234 329112
rect 226978 329060 226984 329112
rect 227036 329100 227042 329112
rect 322198 329100 322204 329112
rect 227036 329072 322204 329100
rect 227036 329060 227042 329072
rect 322198 329060 322204 329072
rect 322256 329060 322262 329112
rect 155880 328624 155908 329060
rect 156874 328624 156880 328636
rect 154546 328596 156880 328624
rect 156874 328584 156880 328596
rect 156932 328584 156938 328636
rect 152292 328528 152504 328556
rect 145392 328460 146984 328488
rect 72896 328392 73108 328420
rect 103486 328392 115428 328420
rect 146956 328420 146984 328460
rect 146956 328392 147674 328420
rect 40678 327700 40684 327752
rect 40736 327740 40742 327752
rect 103486 327740 103514 328392
rect 147646 328284 147674 328392
rect 152476 328352 152504 328528
rect 156690 328448 156696 328500
rect 156748 328488 156754 328500
rect 159450 328488 159456 328500
rect 156748 328460 159456 328488
rect 156748 328448 156754 328460
rect 159450 328448 159456 328460
rect 159508 328448 159514 328500
rect 159542 328448 159548 328500
rect 159600 328488 159606 328500
rect 164970 328488 164976 328500
rect 159600 328460 164976 328488
rect 159600 328448 159606 328460
rect 164970 328448 164976 328460
rect 165028 328448 165034 328500
rect 156874 328352 156880 328364
rect 152476 328324 156880 328352
rect 156874 328312 156880 328324
rect 156932 328312 156938 328364
rect 156690 328284 156696 328296
rect 147646 328256 156696 328284
rect 156690 328244 156696 328256
rect 156748 328244 156754 328296
rect 215110 327768 215116 327820
rect 215168 327808 215174 327820
rect 292574 327808 292580 327820
rect 215168 327780 292580 327808
rect 215168 327768 215174 327780
rect 292574 327768 292580 327780
rect 292632 327768 292638 327820
rect 40736 327712 103514 327740
rect 40736 327700 40742 327712
rect 163314 327700 163320 327752
rect 163372 327740 163378 327752
rect 186958 327740 186964 327752
rect 163372 327712 186964 327740
rect 163372 327700 163378 327712
rect 186958 327700 186964 327712
rect 187016 327700 187022 327752
rect 272610 327700 272616 327752
rect 272668 327740 272674 327752
rect 362954 327740 362960 327752
rect 272668 327712 362960 327740
rect 272668 327700 272674 327712
rect 362954 327700 362960 327712
rect 363012 327700 363018 327752
rect 156690 327088 156696 327140
rect 156748 327128 156754 327140
rect 236730 327128 236736 327140
rect 156748 327100 236736 327128
rect 156748 327088 156754 327100
rect 236730 327088 236736 327100
rect 236788 327088 236794 327140
rect 240042 327088 240048 327140
rect 240100 327128 240106 327140
rect 272610 327128 272616 327140
rect 240100 327100 272616 327128
rect 240100 327088 240106 327100
rect 272610 327088 272616 327100
rect 272668 327088 272674 327140
rect 180058 326408 180064 326460
rect 180116 326448 180122 326460
rect 206462 326448 206468 326460
rect 180116 326420 206468 326448
rect 180116 326408 180122 326420
rect 206462 326408 206468 326420
rect 206520 326408 206526 326460
rect 157058 326340 157064 326392
rect 157116 326380 157122 326392
rect 195238 326380 195244 326392
rect 157116 326352 195244 326380
rect 157116 326340 157122 326352
rect 195238 326340 195244 326352
rect 195296 326340 195302 326392
rect 214558 326340 214564 326392
rect 214616 326380 214622 326392
rect 344278 326380 344284 326392
rect 214616 326352 344284 326380
rect 214616 326340 214622 326352
rect 344278 326340 344284 326352
rect 344336 326340 344342 326392
rect 48222 325660 48228 325712
rect 48280 325700 48286 325712
rect 66254 325700 66260 325712
rect 48280 325672 66260 325700
rect 48280 325660 48286 325672
rect 66254 325660 66260 325672
rect 66312 325660 66318 325712
rect 158714 325660 158720 325712
rect 158772 325700 158778 325712
rect 171134 325700 171140 325712
rect 158772 325672 171140 325700
rect 158772 325660 158778 325672
rect 171134 325660 171140 325672
rect 171192 325660 171198 325712
rect 204990 325660 204996 325712
rect 205048 325700 205054 325712
rect 269114 325700 269120 325712
rect 205048 325672 269120 325700
rect 205048 325660 205054 325672
rect 269114 325660 269120 325672
rect 269172 325660 269178 325712
rect 188522 325592 188528 325644
rect 188580 325632 188586 325644
rect 214558 325632 214564 325644
rect 188580 325604 214564 325632
rect 188580 325592 188586 325604
rect 214558 325592 214564 325604
rect 214616 325592 214622 325644
rect 214558 325116 214564 325168
rect 214616 325156 214622 325168
rect 215110 325156 215116 325168
rect 214616 325128 215116 325156
rect 214616 325116 214622 325128
rect 215110 325116 215116 325128
rect 215168 325116 215174 325168
rect 170490 324980 170496 325032
rect 170548 325020 170554 325032
rect 186314 325020 186320 325032
rect 170548 324992 186320 325020
rect 170548 324980 170554 324992
rect 186314 324980 186320 324992
rect 186372 324980 186378 325032
rect 162118 324912 162124 324964
rect 162176 324952 162182 324964
rect 234430 324952 234436 324964
rect 162176 324924 234436 324952
rect 162176 324912 162182 324924
rect 234430 324912 234436 324924
rect 234488 324952 234494 324964
rect 251910 324952 251916 324964
rect 234488 324924 251916 324952
rect 234488 324912 234494 324924
rect 251910 324912 251916 324924
rect 251968 324912 251974 324964
rect 219710 324300 219716 324352
rect 219768 324340 219774 324352
rect 220170 324340 220176 324352
rect 219768 324312 220176 324340
rect 219768 324300 219774 324312
rect 220170 324300 220176 324312
rect 220228 324340 220234 324352
rect 276658 324340 276664 324352
rect 220228 324312 276664 324340
rect 220228 324300 220234 324312
rect 276658 324300 276664 324312
rect 276716 324300 276722 324352
rect 158806 324164 158812 324216
rect 158864 324204 158870 324216
rect 160738 324204 160744 324216
rect 158864 324176 160744 324204
rect 158864 324164 158870 324176
rect 160738 324164 160744 324176
rect 160796 324164 160802 324216
rect 158714 323008 158720 323060
rect 158772 323048 158778 323060
rect 214650 323048 214656 323060
rect 158772 323020 214656 323048
rect 158772 323008 158778 323020
rect 214650 323008 214656 323020
rect 214708 323008 214714 323060
rect 203610 322940 203616 322992
rect 203668 322980 203674 322992
rect 280798 322980 280804 322992
rect 203668 322952 280804 322980
rect 203668 322940 203674 322952
rect 280798 322940 280804 322952
rect 280856 322940 280862 322992
rect 64782 322872 64788 322924
rect 64840 322912 64846 322924
rect 65794 322912 65800 322924
rect 64840 322884 65800 322912
rect 64840 322872 64846 322884
rect 65794 322872 65800 322884
rect 65852 322872 65858 322924
rect 158714 322804 158720 322856
rect 158772 322844 158778 322856
rect 161566 322844 161572 322856
rect 158772 322816 161572 322844
rect 158772 322804 158778 322816
rect 161566 322804 161572 322816
rect 161624 322804 161630 322856
rect 65794 322396 65800 322448
rect 65852 322436 65858 322448
rect 66530 322436 66536 322448
rect 65852 322408 66536 322436
rect 65852 322396 65858 322408
rect 66530 322396 66536 322408
rect 66588 322396 66594 322448
rect 159450 322260 159456 322312
rect 159508 322300 159514 322312
rect 220170 322300 220176 322312
rect 159508 322272 220176 322300
rect 159508 322260 159514 322272
rect 220170 322260 220176 322272
rect 220228 322260 220234 322312
rect 238018 322260 238024 322312
rect 238076 322300 238082 322312
rect 259638 322300 259644 322312
rect 238076 322272 259644 322300
rect 238076 322260 238082 322272
rect 259638 322260 259644 322272
rect 259696 322260 259702 322312
rect 162946 322192 162952 322244
rect 163004 322232 163010 322244
rect 246298 322232 246304 322244
rect 163004 322204 246304 322232
rect 163004 322192 163010 322204
rect 246298 322192 246304 322204
rect 246356 322192 246362 322244
rect 273990 322192 273996 322244
rect 274048 322232 274054 322244
rect 317598 322232 317604 322244
rect 274048 322204 317604 322232
rect 274048 322192 274054 322204
rect 317598 322192 317604 322204
rect 317656 322192 317662 322244
rect 326982 322192 326988 322244
rect 327040 322232 327046 322244
rect 340230 322232 340236 322244
rect 327040 322204 340236 322232
rect 327040 322192 327046 322204
rect 340230 322192 340236 322204
rect 340288 322192 340294 322244
rect 254670 321580 254676 321632
rect 254728 321620 254734 321632
rect 325694 321620 325700 321632
rect 254728 321592 325700 321620
rect 254728 321580 254734 321592
rect 325694 321580 325700 321592
rect 325752 321620 325758 321632
rect 326982 321620 326988 321632
rect 325752 321592 326988 321620
rect 325752 321580 325758 321592
rect 326982 321580 326988 321592
rect 327040 321580 327046 321632
rect 4798 321512 4804 321564
rect 4856 321552 4862 321564
rect 66806 321552 66812 321564
rect 4856 321524 66812 321552
rect 4856 321512 4862 321524
rect 66806 321512 66812 321524
rect 66864 321512 66870 321564
rect 174906 320900 174912 320952
rect 174964 320940 174970 320952
rect 240870 320940 240876 320952
rect 174964 320912 240876 320940
rect 174964 320900 174970 320912
rect 240870 320900 240876 320912
rect 240928 320900 240934 320952
rect 158162 320832 158168 320884
rect 158220 320872 158226 320884
rect 228542 320872 228548 320884
rect 158220 320844 228548 320872
rect 158220 320832 158226 320844
rect 228542 320832 228548 320844
rect 228600 320832 228606 320884
rect 166902 320560 166908 320612
rect 166960 320600 166966 320612
rect 170490 320600 170496 320612
rect 166960 320572 170496 320600
rect 166960 320560 166966 320572
rect 170490 320560 170496 320572
rect 170548 320560 170554 320612
rect 158714 320152 158720 320204
rect 158772 320192 158778 320204
rect 163682 320192 163688 320204
rect 158772 320164 163688 320192
rect 158772 320152 158778 320164
rect 163682 320152 163688 320164
rect 163740 320152 163746 320204
rect 240870 320152 240876 320204
rect 240928 320192 240934 320204
rect 356698 320192 356704 320204
rect 240928 320164 356704 320192
rect 240928 320152 240934 320164
rect 356698 320152 356704 320164
rect 356756 320152 356762 320204
rect 158806 320084 158812 320136
rect 158864 320124 158870 320136
rect 166902 320124 166908 320136
rect 158864 320096 166908 320124
rect 158864 320084 158870 320096
rect 166902 320084 166908 320096
rect 166960 320084 166966 320136
rect 167638 319472 167644 319524
rect 167696 319512 167702 319524
rect 200482 319512 200488 319524
rect 167696 319484 200488 319512
rect 167696 319472 167702 319484
rect 200482 319472 200488 319484
rect 200540 319472 200546 319524
rect 4062 319404 4068 319456
rect 4120 319444 4126 319456
rect 11698 319444 11704 319456
rect 4120 319416 11704 319444
rect 4120 319404 4126 319416
rect 11698 319404 11704 319416
rect 11756 319404 11762 319456
rect 53742 319404 53748 319456
rect 53800 319444 53806 319456
rect 66438 319444 66444 319456
rect 53800 319416 66444 319444
rect 53800 319404 53806 319416
rect 66438 319404 66444 319416
rect 66496 319404 66502 319456
rect 171134 319404 171140 319456
rect 171192 319444 171198 319456
rect 210418 319444 210424 319456
rect 171192 319416 210424 319444
rect 171192 319404 171198 319416
rect 210418 319404 210424 319416
rect 210476 319404 210482 319456
rect 213362 319404 213368 319456
rect 213420 319444 213426 319456
rect 283558 319444 283564 319456
rect 213420 319416 283564 319444
rect 213420 319404 213426 319416
rect 283558 319404 283564 319416
rect 283616 319404 283622 319456
rect 327810 319404 327816 319456
rect 327868 319444 327874 319456
rect 371418 319444 371424 319456
rect 327868 319416 371424 319444
rect 327868 319404 327874 319416
rect 371418 319404 371424 319416
rect 371476 319404 371482 319456
rect 202782 318792 202788 318844
rect 202840 318832 202846 318844
rect 308398 318832 308404 318844
rect 202840 318804 308404 318832
rect 202840 318792 202846 318804
rect 308398 318792 308404 318804
rect 308456 318792 308462 318844
rect 64598 318588 64604 318640
rect 64656 318628 64662 318640
rect 66438 318628 66444 318640
rect 64656 318600 66444 318628
rect 64656 318588 64662 318600
rect 66438 318588 66444 318600
rect 66496 318588 66502 318640
rect 160830 318112 160836 318164
rect 160888 318152 160894 318164
rect 166442 318152 166448 318164
rect 160888 318124 166448 318152
rect 160888 318112 160894 318124
rect 166442 318112 166448 318124
rect 166500 318112 166506 318164
rect 167914 318112 167920 318164
rect 167972 318152 167978 318164
rect 193950 318152 193956 318164
rect 167972 318124 193956 318152
rect 167972 318112 167978 318124
rect 193950 318112 193956 318124
rect 194008 318112 194014 318164
rect 194042 318112 194048 318164
rect 194100 318152 194106 318164
rect 216030 318152 216036 318164
rect 194100 318124 216036 318152
rect 194100 318112 194106 318124
rect 216030 318112 216036 318124
rect 216088 318112 216094 318164
rect 54938 318044 54944 318096
rect 54996 318084 55002 318096
rect 64138 318084 64144 318096
rect 54996 318056 64144 318084
rect 54996 318044 55002 318056
rect 64138 318044 64144 318056
rect 64196 318044 64202 318096
rect 156782 318044 156788 318096
rect 156840 318084 156846 318096
rect 167822 318084 167828 318096
rect 156840 318056 167828 318084
rect 156840 318044 156846 318056
rect 167822 318044 167828 318056
rect 167880 318044 167886 318096
rect 170582 318044 170588 318096
rect 170640 318084 170646 318096
rect 199562 318084 199568 318096
rect 170640 318056 199568 318084
rect 170640 318044 170646 318056
rect 199562 318044 199568 318056
rect 199620 318044 199626 318096
rect 213270 318044 213276 318096
rect 213328 318084 213334 318096
rect 251266 318084 251272 318096
rect 213328 318056 251272 318084
rect 213328 318044 213334 318056
rect 251266 318044 251272 318056
rect 251324 318044 251330 318096
rect 340874 317500 340880 317552
rect 340932 317540 340938 317552
rect 342162 317540 342168 317552
rect 340932 317512 342168 317540
rect 340932 317500 340938 317512
rect 342162 317500 342168 317512
rect 342220 317540 342226 317552
rect 396718 317540 396724 317552
rect 342220 317512 396724 317540
rect 342220 317500 342226 317512
rect 396718 317500 396724 317512
rect 396776 317500 396782 317552
rect 228450 317432 228456 317484
rect 228508 317472 228514 317484
rect 347038 317472 347044 317484
rect 228508 317444 347044 317472
rect 228508 317432 228514 317444
rect 347038 317432 347044 317444
rect 347096 317432 347102 317484
rect 186314 317364 186320 317416
rect 186372 317404 186378 317416
rect 204990 317404 204996 317416
rect 186372 317376 204996 317404
rect 186372 317364 186378 317376
rect 204990 317364 204996 317376
rect 205048 317364 205054 317416
rect 262398 317364 262404 317416
rect 262456 317404 262462 317416
rect 262858 317404 262864 317416
rect 262456 317376 262864 317404
rect 262456 317364 262462 317376
rect 262858 317364 262864 317376
rect 262916 317364 262922 317416
rect 4798 316684 4804 316736
rect 4856 316724 4862 316736
rect 64506 316724 64512 316736
rect 4856 316696 64512 316724
rect 4856 316684 4862 316696
rect 64506 316684 64512 316696
rect 64564 316724 64570 316736
rect 66898 316724 66904 316736
rect 64564 316696 66904 316724
rect 64564 316684 64570 316696
rect 66898 316684 66904 316696
rect 66956 316684 66962 316736
rect 160002 316684 160008 316736
rect 160060 316724 160066 316736
rect 161290 316724 161296 316736
rect 160060 316696 161296 316724
rect 160060 316684 160066 316696
rect 161290 316684 161296 316696
rect 161348 316724 161354 316736
rect 166350 316724 166356 316736
rect 161348 316696 166356 316724
rect 161348 316684 161354 316696
rect 166350 316684 166356 316696
rect 166408 316684 166414 316736
rect 165062 316480 165068 316532
rect 165120 316520 165126 316532
rect 165522 316520 165528 316532
rect 165120 316492 165528 316520
rect 165120 316480 165126 316492
rect 165522 316480 165528 316492
rect 165580 316480 165586 316532
rect 208118 316072 208124 316124
rect 208176 316112 208182 316124
rect 209774 316112 209780 316124
rect 208176 316084 209780 316112
rect 208176 316072 208182 316084
rect 209774 316072 209780 316084
rect 209832 316112 209838 316124
rect 210970 316112 210976 316124
rect 209832 316084 210976 316112
rect 209832 316072 209838 316084
rect 210970 316072 210976 316084
rect 211028 316072 211034 316124
rect 240134 316072 240140 316124
rect 240192 316112 240198 316124
rect 262398 316112 262404 316124
rect 240192 316084 262404 316112
rect 240192 316072 240198 316084
rect 262398 316072 262404 316084
rect 262456 316072 262462 316124
rect 165062 316004 165068 316056
rect 165120 316044 165126 316056
rect 246390 316044 246396 316056
rect 165120 316016 246396 316044
rect 165120 316004 165126 316016
rect 246390 316004 246396 316016
rect 246448 316004 246454 316056
rect 158806 315936 158812 315988
rect 158864 315976 158870 315988
rect 168282 315976 168288 315988
rect 158864 315948 168288 315976
rect 158864 315936 158870 315948
rect 168282 315936 168288 315948
rect 168340 315936 168346 315988
rect 168282 315324 168288 315376
rect 168340 315364 168346 315376
rect 182818 315364 182824 315376
rect 168340 315336 182824 315364
rect 168340 315324 168346 315336
rect 182818 315324 182824 315336
rect 182876 315324 182882 315376
rect 204898 315324 204904 315376
rect 204956 315364 204962 315376
rect 232682 315364 232688 315376
rect 204956 315336 232688 315364
rect 204956 315324 204962 315336
rect 232682 315324 232688 315336
rect 232740 315324 232746 315376
rect 177482 315256 177488 315308
rect 177540 315296 177546 315308
rect 223022 315296 223028 315308
rect 177540 315268 223028 315296
rect 177540 315256 177546 315268
rect 223022 315256 223028 315268
rect 223080 315256 223086 315308
rect 232590 315256 232596 315308
rect 232648 315296 232654 315308
rect 244366 315296 244372 315308
rect 232648 315268 244372 315296
rect 232648 315256 232654 315268
rect 244366 315256 244372 315268
rect 244424 315256 244430 315308
rect 52086 314644 52092 314696
rect 52144 314684 52150 314696
rect 56502 314684 56508 314696
rect 52144 314656 56508 314684
rect 52144 314644 52150 314656
rect 56502 314644 56508 314656
rect 56560 314684 56566 314696
rect 66806 314684 66812 314696
rect 56560 314656 66812 314684
rect 56560 314644 56566 314656
rect 66806 314644 66812 314656
rect 66864 314644 66870 314696
rect 195974 314644 195980 314696
rect 196032 314684 196038 314696
rect 198734 314684 198740 314696
rect 196032 314656 198740 314684
rect 196032 314644 196038 314656
rect 198734 314644 198740 314656
rect 198792 314644 198798 314696
rect 222470 314644 222476 314696
rect 222528 314684 222534 314696
rect 223022 314684 223028 314696
rect 222528 314656 223028 314684
rect 222528 314644 222534 314656
rect 223022 314644 223028 314656
rect 223080 314684 223086 314696
rect 255498 314684 255504 314696
rect 223080 314656 255504 314684
rect 223080 314644 223086 314656
rect 255498 314644 255504 314656
rect 255556 314644 255562 314696
rect 60366 314576 60372 314628
rect 60424 314616 60430 314628
rect 66898 314616 66904 314628
rect 60424 314588 66904 314616
rect 60424 314576 60430 314588
rect 66898 314576 66904 314588
rect 66956 314576 66962 314628
rect 223482 313896 223488 313948
rect 223540 313936 223546 313948
rect 240134 313936 240140 313948
rect 223540 313908 240140 313936
rect 223540 313896 223546 313908
rect 240134 313896 240140 313908
rect 240192 313896 240198 313948
rect 302326 313896 302332 313948
rect 302384 313936 302390 313948
rect 358814 313936 358820 313948
rect 302384 313908 358820 313936
rect 302384 313896 302390 313908
rect 358814 313896 358820 313908
rect 358872 313896 358878 313948
rect 238570 313352 238576 313404
rect 238628 313392 238634 313404
rect 271874 313392 271880 313404
rect 238628 313364 271880 313392
rect 238628 313352 238634 313364
rect 271874 313352 271880 313364
rect 271932 313392 271938 313404
rect 272518 313392 272524 313404
rect 271932 313364 272524 313392
rect 271932 313352 271938 313364
rect 272518 313352 272524 313364
rect 272576 313352 272582 313404
rect 158806 313284 158812 313336
rect 158864 313324 158870 313336
rect 192478 313324 192484 313336
rect 158864 313296 192484 313324
rect 158864 313284 158870 313296
rect 192478 313284 192484 313296
rect 192536 313284 192542 313336
rect 241974 313284 241980 313336
rect 242032 313324 242038 313336
rect 242250 313324 242256 313336
rect 242032 313296 242256 313324
rect 242032 313284 242038 313296
rect 242250 313284 242256 313296
rect 242308 313324 242314 313336
rect 302326 313324 302332 313336
rect 242308 313296 302332 313324
rect 242308 313284 242314 313296
rect 302326 313284 302332 313296
rect 302384 313284 302390 313336
rect 161566 312536 161572 312588
rect 161624 312576 161630 312588
rect 235350 312576 235356 312588
rect 161624 312548 235356 312576
rect 161624 312536 161630 312548
rect 235350 312536 235356 312548
rect 235408 312536 235414 312588
rect 293218 312536 293224 312588
rect 293276 312576 293282 312588
rect 338758 312576 338764 312588
rect 293276 312548 338764 312576
rect 293276 312536 293282 312548
rect 338758 312536 338764 312548
rect 338816 312536 338822 312588
rect 202138 311856 202144 311908
rect 202196 311896 202202 311908
rect 209222 311896 209228 311908
rect 202196 311868 209228 311896
rect 202196 311856 202202 311868
rect 209222 311856 209228 311868
rect 209280 311856 209286 311908
rect 227806 311856 227812 311908
rect 227864 311896 227870 311908
rect 228542 311896 228548 311908
rect 227864 311868 228548 311896
rect 227864 311856 227870 311868
rect 228542 311856 228548 311868
rect 228600 311896 228606 311908
rect 282914 311896 282920 311908
rect 228600 311868 282920 311896
rect 228600 311856 228606 311868
rect 282914 311856 282920 311868
rect 282972 311856 282978 311908
rect 238110 311788 238116 311840
rect 238168 311828 238174 311840
rect 239398 311828 239404 311840
rect 238168 311800 239404 311828
rect 238168 311788 238174 311800
rect 239398 311788 239404 311800
rect 239456 311788 239462 311840
rect 187602 311176 187608 311228
rect 187660 311216 187666 311228
rect 194594 311216 194600 311228
rect 187660 311188 194600 311216
rect 187660 311176 187666 311188
rect 194594 311176 194600 311188
rect 194652 311216 194658 311228
rect 238018 311216 238024 311228
rect 194652 311188 238024 311216
rect 194652 311176 194658 311188
rect 238018 311176 238024 311188
rect 238076 311176 238082 311228
rect 239398 311176 239404 311228
rect 239456 311216 239462 311228
rect 239582 311216 239588 311228
rect 239456 311188 239588 311216
rect 239456 311176 239462 311188
rect 239582 311176 239588 311188
rect 239640 311216 239646 311228
rect 254670 311216 254676 311228
rect 239640 311188 254676 311216
rect 239640 311176 239646 311188
rect 254670 311176 254676 311188
rect 254728 311176 254734 311228
rect 11698 311108 11704 311160
rect 11756 311148 11762 311160
rect 67082 311148 67088 311160
rect 11756 311120 67088 311148
rect 11756 311108 11762 311120
rect 67082 311108 67088 311120
rect 67140 311148 67146 311160
rect 67450 311148 67456 311160
rect 67140 311120 67456 311148
rect 67140 311108 67146 311120
rect 67450 311108 67456 311120
rect 67508 311108 67514 311160
rect 197170 311108 197176 311160
rect 197228 311148 197234 311160
rect 287698 311148 287704 311160
rect 197228 311120 287704 311148
rect 197228 311108 197234 311120
rect 287698 311108 287704 311120
rect 287756 311108 287762 311160
rect 158898 310496 158904 310548
rect 158956 310536 158962 310548
rect 194594 310536 194600 310548
rect 158956 310508 194600 310536
rect 158956 310496 158962 310508
rect 194594 310496 194600 310508
rect 194652 310496 194658 310548
rect 158806 310428 158812 310480
rect 158864 310468 158870 310480
rect 164234 310468 164240 310480
rect 158864 310440 164240 310468
rect 158864 310428 158870 310440
rect 164234 310428 164240 310440
rect 164292 310468 164298 310480
rect 165522 310468 165528 310480
rect 164292 310440 165528 310468
rect 164292 310428 164298 310440
rect 165522 310428 165528 310440
rect 165580 310428 165586 310480
rect 238662 310428 238668 310480
rect 238720 310468 238726 310480
rect 240226 310468 240232 310480
rect 238720 310440 240232 310468
rect 238720 310428 238726 310440
rect 240226 310428 240232 310440
rect 240284 310428 240290 310480
rect 165522 309816 165528 309868
rect 165580 309856 165586 309868
rect 177482 309856 177488 309868
rect 165580 309828 177488 309856
rect 165580 309816 165586 309828
rect 177482 309816 177488 309828
rect 177540 309816 177546 309868
rect 35158 309748 35164 309800
rect 35216 309788 35222 309800
rect 62758 309788 62764 309800
rect 35216 309760 62764 309788
rect 35216 309748 35222 309760
rect 62758 309748 62764 309760
rect 62816 309788 62822 309800
rect 66806 309788 66812 309800
rect 62816 309760 66812 309788
rect 62816 309748 62822 309760
rect 66806 309748 66812 309760
rect 66864 309748 66870 309800
rect 171962 309748 171968 309800
rect 172020 309788 172026 309800
rect 223482 309788 223488 309800
rect 172020 309760 223488 309788
rect 172020 309748 172026 309760
rect 223482 309748 223488 309760
rect 223540 309748 223546 309800
rect 262122 309748 262128 309800
rect 262180 309788 262186 309800
rect 313918 309788 313924 309800
rect 262180 309760 313924 309788
rect 262180 309748 262186 309760
rect 313918 309748 313924 309760
rect 313976 309748 313982 309800
rect 208486 309136 208492 309188
rect 208544 309176 208550 309188
rect 209222 309176 209228 309188
rect 208544 309148 209228 309176
rect 208544 309136 208550 309148
rect 209222 309136 209228 309148
rect 209280 309176 209286 309188
rect 279418 309176 279424 309188
rect 209280 309148 279424 309176
rect 209280 309136 209286 309148
rect 279418 309136 279424 309148
rect 279476 309136 279482 309188
rect 158806 308932 158812 308984
rect 158864 308972 158870 308984
rect 162854 308972 162860 308984
rect 158864 308944 162860 308972
rect 158864 308932 158870 308944
rect 162854 308932 162860 308944
rect 162912 308972 162918 308984
rect 166534 308972 166540 308984
rect 162912 308944 166540 308972
rect 162912 308932 162918 308944
rect 166534 308932 166540 308944
rect 166592 308932 166598 308984
rect 282178 307884 282184 307896
rect 200086 307856 282184 307884
rect 200086 307828 200114 307856
rect 282178 307844 282184 307856
rect 282236 307844 282242 307896
rect 199562 307776 199568 307828
rect 199620 307816 199626 307828
rect 200022 307816 200028 307828
rect 199620 307788 200028 307816
rect 199620 307776 199626 307788
rect 200022 307776 200028 307788
rect 200080 307788 200114 307828
rect 200080 307776 200086 307788
rect 239030 307776 239036 307828
rect 239088 307816 239094 307828
rect 381538 307816 381544 307828
rect 239088 307788 381544 307816
rect 239088 307776 239094 307788
rect 381538 307776 381544 307788
rect 381596 307776 381602 307828
rect 61746 307708 61752 307760
rect 61804 307748 61810 307760
rect 66898 307748 66904 307760
rect 61804 307720 66904 307748
rect 61804 307708 61810 307720
rect 66898 307708 66904 307720
rect 66956 307708 66962 307760
rect 197078 307096 197084 307148
rect 197136 307136 197142 307148
rect 204346 307136 204352 307148
rect 197136 307108 204352 307136
rect 197136 307096 197142 307108
rect 204346 307096 204352 307108
rect 204404 307096 204410 307148
rect 190270 307028 190276 307080
rect 190328 307068 190334 307080
rect 204254 307068 204260 307080
rect 190328 307040 204260 307068
rect 190328 307028 190334 307040
rect 204254 307028 204260 307040
rect 204312 307028 204318 307080
rect 207750 306416 207756 306468
rect 207808 306456 207814 306468
rect 243998 306456 244004 306468
rect 207808 306428 244004 306456
rect 207808 306416 207814 306428
rect 243998 306416 244004 306428
rect 244056 306416 244062 306468
rect 158806 306348 158812 306400
rect 158864 306388 158870 306400
rect 170398 306388 170404 306400
rect 158864 306360 170404 306388
rect 158864 306348 158870 306360
rect 170398 306348 170404 306360
rect 170456 306348 170462 306400
rect 209406 306348 209412 306400
rect 209464 306388 209470 306400
rect 267090 306388 267096 306400
rect 209464 306360 267096 306388
rect 209464 306348 209470 306360
rect 267090 306348 267096 306360
rect 267148 306348 267154 306400
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 33778 306320 33784 306332
rect 3384 306292 33784 306320
rect 3384 306280 3390 306292
rect 33778 306280 33784 306292
rect 33836 306280 33842 306332
rect 310422 305600 310428 305652
rect 310480 305640 310486 305652
rect 363230 305640 363236 305652
rect 310480 305612 363236 305640
rect 310480 305600 310486 305612
rect 363230 305600 363236 305612
rect 363288 305600 363294 305652
rect 199470 305056 199476 305108
rect 199528 305096 199534 305108
rect 200114 305096 200120 305108
rect 199528 305068 200120 305096
rect 199528 305056 199534 305068
rect 200114 305056 200120 305068
rect 200172 305096 200178 305108
rect 201402 305096 201408 305108
rect 200172 305068 201408 305096
rect 200172 305056 200178 305068
rect 201402 305056 201408 305068
rect 201460 305056 201466 305108
rect 212718 305056 212724 305108
rect 212776 305096 212782 305108
rect 267826 305096 267832 305108
rect 212776 305068 267832 305096
rect 212776 305056 212782 305068
rect 267826 305056 267832 305068
rect 267884 305056 267890 305108
rect 56410 304988 56416 305040
rect 56468 305028 56474 305040
rect 66806 305028 66812 305040
rect 56468 305000 66812 305028
rect 56468 304988 56474 305000
rect 66806 304988 66812 305000
rect 66864 304988 66870 305040
rect 158806 304988 158812 305040
rect 158864 305028 158870 305040
rect 235994 305028 236000 305040
rect 158864 305000 236000 305028
rect 158864 304988 158870 305000
rect 235994 304988 236000 305000
rect 236052 304988 236058 305040
rect 236086 304988 236092 305040
rect 236144 305028 236150 305040
rect 236730 305028 236736 305040
rect 236144 305000 236736 305028
rect 236144 304988 236150 305000
rect 236730 304988 236736 305000
rect 236788 305028 236794 305040
rect 236788 305000 294000 305028
rect 236788 304988 236794 305000
rect 293972 304960 294000 305000
rect 294598 304960 294604 304972
rect 293972 304932 294604 304960
rect 294598 304920 294604 304932
rect 294656 304960 294662 304972
rect 367094 304960 367100 304972
rect 294656 304932 367100 304960
rect 294656 304920 294662 304932
rect 367094 304920 367100 304932
rect 367152 304920 367158 304972
rect 175182 304308 175188 304360
rect 175240 304348 175246 304360
rect 188430 304348 188436 304360
rect 175240 304320 188436 304348
rect 175240 304308 175246 304320
rect 188430 304308 188436 304320
rect 188488 304308 188494 304360
rect 192754 304308 192760 304360
rect 192812 304348 192818 304360
rect 220170 304348 220176 304360
rect 192812 304320 220176 304348
rect 192812 304308 192818 304320
rect 220170 304308 220176 304320
rect 220228 304308 220234 304360
rect 234522 304308 234528 304360
rect 234580 304348 234586 304360
rect 280982 304348 280988 304360
rect 234580 304320 280988 304348
rect 234580 304308 234586 304320
rect 280982 304308 280988 304320
rect 281040 304308 281046 304360
rect 184290 304240 184296 304292
rect 184348 304280 184354 304292
rect 208946 304280 208952 304292
rect 184348 304252 208952 304280
rect 184348 304240 184354 304252
rect 208946 304240 208952 304252
rect 209004 304240 209010 304292
rect 209038 304240 209044 304292
rect 209096 304280 209102 304292
rect 215202 304280 215208 304292
rect 209096 304252 215208 304280
rect 209096 304240 209102 304252
rect 215202 304240 215208 304252
rect 215260 304280 215266 304292
rect 358078 304280 358084 304292
rect 215260 304252 358084 304280
rect 215260 304240 215266 304252
rect 358078 304240 358084 304252
rect 358136 304240 358142 304292
rect 158806 303968 158812 304020
rect 158864 304008 158870 304020
rect 160830 304008 160836 304020
rect 158864 303980 160836 304008
rect 158864 303968 158870 303980
rect 160830 303968 160836 303980
rect 160888 303968 160894 304020
rect 158806 303628 158812 303680
rect 158864 303668 158870 303680
rect 175182 303668 175188 303680
rect 158864 303640 175188 303668
rect 158864 303628 158870 303640
rect 175182 303628 175188 303640
rect 175240 303628 175246 303680
rect 231670 303628 231676 303680
rect 231728 303668 231734 303680
rect 234522 303668 234528 303680
rect 231728 303640 234528 303668
rect 231728 303628 231734 303640
rect 234522 303628 234528 303640
rect 234580 303628 234586 303680
rect 64690 303560 64696 303612
rect 64748 303600 64754 303612
rect 66898 303600 66904 303612
rect 64748 303572 66904 303600
rect 64748 303560 64754 303572
rect 66898 303560 66904 303572
rect 66956 303560 66962 303612
rect 193398 302880 193404 302932
rect 193456 302920 193462 302932
rect 212718 302920 212724 302932
rect 193456 302892 212724 302920
rect 193456 302880 193462 302892
rect 212718 302880 212724 302892
rect 212776 302880 212782 302932
rect 322198 302880 322204 302932
rect 322256 302920 322262 302932
rect 355318 302920 355324 302932
rect 322256 302892 355324 302920
rect 322256 302880 322262 302892
rect 355318 302880 355324 302892
rect 355376 302880 355382 302932
rect 202230 302268 202236 302320
rect 202288 302308 202294 302320
rect 274082 302308 274088 302320
rect 202288 302280 274088 302308
rect 202288 302268 202294 302280
rect 274082 302268 274088 302280
rect 274140 302268 274146 302320
rect 215294 302200 215300 302252
rect 215352 302240 215358 302252
rect 215846 302240 215852 302252
rect 215352 302212 215852 302240
rect 215352 302200 215358 302212
rect 215846 302200 215852 302212
rect 215904 302240 215910 302252
rect 288434 302240 288440 302252
rect 215904 302212 288440 302240
rect 215904 302200 215910 302212
rect 288434 302200 288440 302212
rect 288492 302200 288498 302252
rect 58986 302132 58992 302184
rect 59044 302172 59050 302184
rect 66898 302172 66904 302184
rect 59044 302144 66904 302172
rect 59044 302132 59050 302144
rect 66898 302132 66904 302144
rect 66956 302132 66962 302184
rect 164970 301520 164976 301572
rect 165028 301560 165034 301572
rect 251358 301560 251364 301572
rect 165028 301532 251364 301560
rect 165028 301520 165034 301532
rect 251358 301520 251364 301532
rect 251416 301520 251422 301572
rect 262950 301520 262956 301572
rect 263008 301560 263014 301572
rect 293954 301560 293960 301572
rect 263008 301532 293960 301560
rect 263008 301520 263014 301532
rect 293954 301520 293960 301532
rect 294012 301520 294018 301572
rect 327718 301520 327724 301572
rect 327776 301560 327782 301572
rect 330478 301560 330484 301572
rect 327776 301532 330484 301560
rect 327776 301520 327782 301532
rect 330478 301520 330484 301532
rect 330536 301520 330542 301572
rect 160002 301452 160008 301504
rect 160060 301492 160066 301504
rect 165614 301492 165620 301504
rect 160060 301464 165620 301492
rect 160060 301452 160066 301464
rect 165614 301452 165620 301464
rect 165672 301492 165678 301504
rect 166074 301492 166080 301504
rect 165672 301464 166080 301492
rect 165672 301452 165678 301464
rect 166074 301452 166080 301464
rect 166132 301452 166138 301504
rect 193858 301452 193864 301504
rect 193916 301492 193922 301504
rect 221550 301492 221556 301504
rect 193916 301464 221556 301492
rect 193916 301452 193922 301464
rect 221550 301452 221556 301464
rect 221608 301452 221614 301504
rect 238018 301452 238024 301504
rect 238076 301492 238082 301504
rect 353938 301492 353944 301504
rect 238076 301464 353944 301492
rect 238076 301452 238082 301464
rect 353938 301452 353944 301464
rect 353996 301452 354002 301504
rect 64690 300840 64696 300892
rect 64748 300880 64754 300892
rect 66806 300880 66812 300892
rect 64748 300852 66812 300880
rect 64748 300840 64754 300852
rect 66806 300840 66812 300852
rect 66864 300840 66870 300892
rect 158990 300296 158996 300348
rect 159048 300336 159054 300348
rect 160094 300336 160100 300348
rect 159048 300308 160100 300336
rect 159048 300296 159054 300308
rect 160094 300296 160100 300308
rect 160152 300336 160158 300348
rect 160922 300336 160928 300348
rect 160152 300308 160928 300336
rect 160152 300296 160158 300308
rect 160922 300296 160928 300308
rect 160980 300296 160986 300348
rect 163682 300160 163688 300212
rect 163740 300200 163746 300212
rect 245746 300200 245752 300212
rect 163740 300172 245752 300200
rect 163740 300160 163746 300172
rect 245746 300160 245752 300172
rect 245804 300160 245810 300212
rect 158806 300092 158812 300144
rect 158864 300132 158870 300144
rect 244458 300132 244464 300144
rect 158864 300104 244464 300132
rect 158864 300092 158870 300104
rect 244458 300092 244464 300104
rect 244516 300092 244522 300144
rect 249150 299480 249156 299532
rect 249208 299520 249214 299532
rect 442994 299520 443000 299532
rect 249208 299492 443000 299520
rect 249208 299480 249214 299492
rect 442994 299480 443000 299492
rect 443052 299480 443058 299532
rect 56318 299412 56324 299464
rect 56376 299452 56382 299464
rect 66622 299452 66628 299464
rect 56376 299424 66628 299452
rect 56376 299412 56382 299424
rect 66622 299412 66628 299424
rect 66680 299412 66686 299464
rect 158806 299412 158812 299464
rect 158864 299452 158870 299464
rect 173250 299452 173256 299464
rect 158864 299424 173256 299452
rect 158864 299412 158870 299424
rect 173250 299412 173256 299424
rect 173308 299412 173314 299464
rect 180242 298800 180248 298852
rect 180300 298840 180306 298852
rect 230382 298840 230388 298852
rect 180300 298812 230388 298840
rect 180300 298800 180306 298812
rect 230382 298800 230388 298812
rect 230440 298800 230446 298852
rect 243446 298800 243452 298852
rect 243504 298840 243510 298852
rect 245654 298840 245660 298852
rect 243504 298812 245660 298840
rect 243504 298800 243510 298812
rect 245654 298800 245660 298812
rect 245712 298840 245718 298852
rect 245712 298812 296714 298840
rect 245712 298800 245718 298812
rect 201310 298732 201316 298784
rect 201368 298772 201374 298784
rect 254670 298772 254676 298784
rect 201368 298744 254676 298772
rect 201368 298732 201374 298744
rect 254670 298732 254676 298744
rect 254728 298732 254734 298784
rect 296686 298772 296714 298812
rect 298094 298772 298100 298784
rect 296686 298744 298100 298772
rect 298094 298732 298100 298744
rect 298152 298772 298158 298784
rect 369854 298772 369860 298784
rect 298152 298744 369860 298772
rect 298152 298732 298158 298744
rect 369854 298732 369860 298744
rect 369912 298732 369918 298784
rect 194318 298120 194324 298172
rect 194376 298160 194382 298172
rect 200298 298160 200304 298172
rect 194376 298132 200304 298160
rect 194376 298120 194382 298132
rect 200298 298120 200304 298132
rect 200356 298160 200362 298172
rect 201310 298160 201316 298172
rect 200356 298132 201316 298160
rect 200356 298120 200362 298132
rect 201310 298120 201316 298132
rect 201368 298120 201374 298172
rect 57882 298052 57888 298104
rect 57940 298092 57946 298104
rect 58986 298092 58992 298104
rect 57940 298064 58992 298092
rect 57940 298052 57946 298064
rect 58986 298052 58992 298064
rect 59044 298052 59050 298104
rect 193950 297508 193956 297560
rect 194008 297548 194014 297560
rect 204254 297548 204260 297560
rect 194008 297520 204260 297548
rect 194008 297508 194014 297520
rect 204254 297508 204260 297520
rect 204312 297508 204318 297560
rect 167822 297440 167828 297492
rect 167880 297480 167886 297492
rect 180242 297480 180248 297492
rect 167880 297452 180248 297480
rect 167880 297440 167886 297452
rect 180242 297440 180248 297452
rect 180300 297440 180306 297492
rect 183370 297440 183376 297492
rect 183428 297480 183434 297492
rect 203518 297480 203524 297492
rect 183428 297452 203524 297480
rect 183428 297440 183434 297452
rect 203518 297440 203524 297452
rect 203576 297440 203582 297492
rect 58986 297372 58992 297424
rect 59044 297412 59050 297424
rect 66806 297412 66812 297424
rect 59044 297384 66812 297412
rect 59044 297372 59050 297384
rect 66806 297372 66812 297384
rect 66864 297372 66870 297424
rect 165154 297372 165160 297424
rect 165212 297412 165218 297424
rect 193398 297412 193404 297424
rect 165212 297384 193404 297412
rect 165212 297372 165218 297384
rect 193398 297372 193404 297384
rect 193456 297372 193462 297424
rect 246390 297372 246396 297424
rect 246448 297412 246454 297424
rect 256694 297412 256700 297424
rect 246448 297384 256700 297412
rect 246448 297372 246454 297384
rect 256694 297372 256700 297384
rect 256752 297372 256758 297424
rect 158806 296692 158812 296744
rect 158864 296732 158870 296744
rect 168282 296732 168288 296744
rect 158864 296704 168288 296732
rect 158864 296692 158870 296704
rect 168282 296692 168288 296704
rect 168340 296692 168346 296744
rect 231118 296692 231124 296744
rect 231176 296732 231182 296744
rect 247126 296732 247132 296744
rect 231176 296704 247132 296732
rect 231176 296692 231182 296704
rect 247126 296692 247132 296704
rect 247184 296692 247190 296744
rect 166810 296012 166816 296064
rect 166868 296052 166874 296064
rect 187050 296052 187056 296064
rect 166868 296024 187056 296052
rect 166868 296012 166874 296024
rect 187050 296012 187056 296024
rect 187108 296012 187114 296064
rect 158806 295944 158812 295996
rect 158864 295984 158870 295996
rect 209038 295984 209044 295996
rect 158864 295956 209044 295984
rect 158864 295944 158870 295956
rect 209038 295944 209044 295956
rect 209096 295944 209102 295996
rect 214558 295400 214564 295452
rect 214616 295440 214622 295452
rect 224310 295440 224316 295452
rect 214616 295412 224316 295440
rect 214616 295400 214622 295412
rect 224310 295400 224316 295412
rect 224368 295400 224374 295452
rect 273162 295400 273168 295452
rect 273220 295440 273226 295452
rect 278222 295440 278228 295452
rect 273220 295412 278228 295440
rect 273220 295400 273226 295412
rect 278222 295400 278228 295412
rect 278280 295400 278286 295452
rect 30282 295332 30288 295384
rect 30340 295372 30346 295384
rect 67174 295372 67180 295384
rect 30340 295344 67180 295372
rect 30340 295332 30346 295344
rect 67174 295332 67180 295344
rect 67232 295332 67238 295384
rect 189902 295332 189908 295384
rect 189960 295372 189966 295384
rect 190362 295372 190368 295384
rect 189960 295344 190368 295372
rect 189960 295332 189966 295344
rect 190362 295332 190368 295344
rect 190420 295372 190426 295384
rect 439406 295372 439412 295384
rect 190420 295344 439412 295372
rect 190420 295332 190426 295344
rect 439406 295332 439412 295344
rect 439464 295332 439470 295384
rect 158806 295264 158812 295316
rect 158864 295304 158870 295316
rect 177390 295304 177396 295316
rect 158864 295276 177396 295304
rect 158864 295264 158870 295276
rect 177390 295264 177396 295276
rect 177448 295264 177454 295316
rect 235258 295264 235264 295316
rect 235316 295304 235322 295316
rect 392670 295304 392676 295316
rect 235316 295276 392676 295304
rect 235316 295264 235322 295276
rect 392670 295264 392676 295276
rect 392728 295264 392734 295316
rect 392670 294584 392676 294636
rect 392728 294624 392734 294636
rect 414658 294624 414664 294636
rect 392728 294596 414664 294624
rect 392728 294584 392734 294596
rect 414658 294584 414664 294596
rect 414716 294584 414722 294636
rect 177298 294040 177304 294092
rect 177356 294080 177362 294092
rect 202230 294080 202236 294092
rect 177356 294052 202236 294080
rect 177356 294040 177362 294052
rect 202230 294040 202236 294052
rect 202288 294040 202294 294092
rect 195330 293972 195336 294024
rect 195388 294012 195394 294024
rect 259730 294012 259736 294024
rect 195388 293984 259736 294012
rect 195388 293972 195394 293984
rect 259730 293972 259736 293984
rect 259788 293972 259794 294024
rect 26142 293904 26148 293956
rect 26200 293944 26206 293956
rect 66806 293944 66812 293956
rect 26200 293916 66812 293944
rect 26200 293904 26206 293916
rect 66806 293904 66812 293916
rect 66864 293904 66870 293956
rect 158806 292612 158812 292664
rect 158864 292652 158870 292664
rect 193858 292652 193864 292664
rect 158864 292624 193864 292652
rect 158864 292612 158870 292624
rect 193858 292612 193864 292624
rect 193916 292612 193922 292664
rect 253198 292652 253204 292664
rect 229066 292624 253204 292652
rect 3602 292544 3608 292596
rect 3660 292584 3666 292596
rect 18598 292584 18604 292596
rect 3660 292556 18604 292584
rect 3660 292544 3666 292556
rect 18598 292544 18604 292556
rect 18656 292544 18662 292596
rect 158898 292544 158904 292596
rect 158956 292584 158962 292596
rect 220170 292584 220176 292596
rect 158956 292556 220176 292584
rect 158956 292544 158962 292556
rect 220170 292544 220176 292556
rect 220228 292544 220234 292596
rect 221550 292544 221556 292596
rect 221608 292584 221614 292596
rect 222102 292584 222108 292596
rect 221608 292556 222108 292584
rect 221608 292544 221614 292556
rect 222102 292544 222108 292556
rect 222160 292584 222166 292596
rect 229066 292584 229094 292624
rect 253198 292612 253204 292624
rect 253256 292612 253262 292664
rect 222160 292556 229094 292584
rect 222160 292544 222166 292556
rect 234430 292544 234436 292596
rect 234488 292584 234494 292596
rect 295426 292584 295432 292596
rect 234488 292556 295432 292584
rect 234488 292544 234494 292556
rect 295426 292544 295432 292556
rect 295484 292544 295490 292596
rect 53558 292476 53564 292528
rect 53616 292516 53622 292528
rect 66806 292516 66812 292528
rect 53616 292488 66812 292516
rect 53616 292476 53622 292488
rect 66806 292476 66812 292488
rect 66864 292476 66870 292528
rect 247126 291796 247132 291848
rect 247184 291836 247190 291848
rect 253934 291836 253940 291848
rect 247184 291808 253940 291836
rect 247184 291796 247190 291808
rect 253934 291796 253940 291808
rect 253992 291796 253998 291848
rect 256050 291796 256056 291848
rect 256108 291836 256114 291848
rect 263778 291836 263784 291848
rect 256108 291808 263784 291836
rect 256108 291796 256114 291808
rect 263778 291796 263784 291808
rect 263836 291796 263842 291848
rect 187510 291320 187516 291372
rect 187568 291360 187574 291372
rect 192570 291360 192576 291372
rect 187568 291332 192576 291360
rect 187568 291320 187574 291332
rect 192570 291320 192576 291332
rect 192628 291320 192634 291372
rect 195146 291252 195152 291304
rect 195204 291292 195210 291304
rect 247310 291292 247316 291304
rect 195204 291264 247316 291292
rect 195204 291252 195210 291264
rect 247310 291252 247316 291264
rect 247368 291252 247374 291304
rect 158806 291184 158812 291236
rect 158864 291224 158870 291236
rect 247126 291224 247132 291236
rect 158864 291196 247132 291224
rect 158864 291184 158870 291196
rect 247126 291184 247132 291196
rect 247184 291184 247190 291236
rect 60458 291116 60464 291168
rect 60516 291156 60522 291168
rect 66346 291156 66352 291168
rect 60516 291128 66352 291156
rect 60516 291116 60522 291128
rect 66346 291116 66352 291128
rect 66404 291116 66410 291168
rect 59170 291048 59176 291100
rect 59228 291088 59234 291100
rect 67082 291088 67088 291100
rect 59228 291060 67088 291088
rect 59228 291048 59234 291060
rect 67082 291048 67088 291060
rect 67140 291048 67146 291100
rect 199562 290776 199568 290828
rect 199620 290816 199626 290828
rect 201494 290816 201500 290828
rect 199620 290788 201500 290816
rect 199620 290776 199626 290788
rect 201494 290776 201500 290788
rect 201552 290776 201558 290828
rect 162210 290436 162216 290488
rect 162268 290476 162274 290488
rect 195146 290476 195152 290488
rect 162268 290448 195152 290476
rect 162268 290436 162274 290448
rect 195146 290436 195152 290448
rect 195204 290436 195210 290488
rect 295886 290436 295892 290488
rect 295944 290476 295950 290488
rect 371234 290476 371240 290488
rect 295944 290448 371240 290476
rect 295944 290436 295950 290448
rect 371234 290436 371240 290448
rect 371292 290436 371298 290488
rect 210418 289892 210424 289944
rect 210476 289932 210482 289944
rect 248414 289932 248420 289944
rect 210476 289904 248420 289932
rect 210476 289892 210482 289904
rect 248414 289892 248420 289904
rect 248472 289892 248478 289944
rect 158806 289824 158812 289876
rect 158864 289864 158870 289876
rect 216674 289864 216680 289876
rect 158864 289836 216680 289864
rect 158864 289824 158870 289836
rect 216674 289824 216680 289836
rect 216732 289824 216738 289876
rect 229738 289824 229744 289876
rect 229796 289864 229802 289876
rect 255314 289864 255320 289876
rect 229796 289836 255320 289864
rect 229796 289824 229802 289836
rect 255314 289824 255320 289836
rect 255372 289824 255378 289876
rect 258902 289824 258908 289876
rect 258960 289864 258966 289876
rect 322290 289864 322296 289876
rect 258960 289836 322296 289864
rect 258960 289824 258966 289836
rect 322290 289824 322296 289836
rect 322348 289824 322354 289876
rect 186958 289756 186964 289808
rect 187016 289796 187022 289808
rect 188430 289796 188436 289808
rect 187016 289768 188436 289796
rect 187016 289756 187022 289768
rect 188430 289756 188436 289768
rect 188488 289756 188494 289808
rect 64138 289212 64144 289264
rect 64196 289252 64202 289264
rect 66806 289252 66812 289264
rect 64196 289224 66812 289252
rect 64196 289212 64202 289224
rect 66806 289212 66812 289224
rect 66864 289212 66870 289264
rect 158806 289212 158812 289264
rect 158864 289252 158870 289264
rect 162762 289252 162768 289264
rect 158864 289224 162768 289252
rect 158864 289212 158870 289224
rect 162762 289212 162768 289224
rect 162820 289212 162826 289264
rect 169018 289076 169024 289128
rect 169076 289116 169082 289128
rect 181438 289116 181444 289128
rect 169076 289088 181444 289116
rect 169076 289076 169082 289088
rect 181438 289076 181444 289088
rect 181496 289076 181502 289128
rect 216674 289076 216680 289128
rect 216732 289116 216738 289128
rect 224862 289116 224868 289128
rect 216732 289088 224868 289116
rect 216732 289076 216738 289088
rect 224862 289076 224868 289088
rect 224920 289076 224926 289128
rect 240502 289076 240508 289128
rect 240560 289116 240566 289128
rect 258902 289116 258908 289128
rect 240560 289088 258908 289116
rect 240560 289076 240566 289088
rect 258902 289076 258908 289088
rect 258960 289076 258966 289128
rect 200022 288464 200028 288516
rect 200080 288504 200086 288516
rect 201678 288504 201684 288516
rect 200080 288476 201684 288504
rect 200080 288464 200086 288476
rect 201678 288464 201684 288476
rect 201736 288464 201742 288516
rect 176102 288396 176108 288448
rect 176160 288436 176166 288448
rect 216674 288436 216680 288448
rect 176160 288408 216680 288436
rect 176160 288396 176166 288408
rect 216674 288396 216680 288408
rect 216732 288396 216738 288448
rect 224862 288396 224868 288448
rect 224920 288436 224926 288448
rect 247494 288436 247500 288448
rect 224920 288408 247500 288436
rect 224920 288396 224926 288408
rect 247494 288396 247500 288408
rect 247552 288396 247558 288448
rect 332594 288396 332600 288448
rect 332652 288436 332658 288448
rect 447134 288436 447140 288448
rect 332652 288408 447140 288436
rect 332652 288396 332658 288408
rect 447134 288396 447140 288408
rect 447192 288396 447198 288448
rect 158898 288328 158904 288380
rect 158956 288368 158962 288380
rect 231118 288368 231124 288380
rect 158956 288340 231124 288368
rect 158956 288328 158962 288340
rect 231118 288328 231124 288340
rect 231176 288328 231182 288380
rect 259546 288192 259552 288244
rect 259604 288232 259610 288244
rect 260098 288232 260104 288244
rect 259604 288204 260104 288232
rect 259604 288192 259610 288204
rect 260098 288192 260104 288204
rect 260156 288192 260162 288244
rect 66162 287784 66168 287836
rect 66220 287824 66226 287836
rect 67358 287824 67364 287836
rect 66220 287796 67364 287824
rect 66220 287784 66226 287796
rect 67358 287784 67364 287796
rect 67416 287784 67422 287836
rect 164970 287648 164976 287700
rect 165028 287688 165034 287700
rect 195146 287688 195152 287700
rect 165028 287660 195152 287688
rect 165028 287648 165034 287660
rect 195146 287648 195152 287660
rect 195204 287648 195210 287700
rect 235350 287648 235356 287700
rect 235408 287688 235414 287700
rect 245838 287688 245844 287700
rect 235408 287660 245844 287688
rect 235408 287648 235414 287660
rect 245838 287648 245844 287660
rect 245896 287648 245902 287700
rect 303614 287648 303620 287700
rect 303672 287688 303678 287700
rect 364334 287688 364340 287700
rect 303672 287660 364340 287688
rect 303672 287648 303678 287660
rect 364334 287648 364340 287660
rect 364392 287648 364398 287700
rect 376110 287648 376116 287700
rect 376168 287688 376174 287700
rect 392578 287688 392584 287700
rect 376168 287660 392584 287688
rect 376168 287648 376174 287660
rect 392578 287648 392584 287660
rect 392636 287648 392642 287700
rect 233142 287104 233148 287156
rect 233200 287144 233206 287156
rect 260098 287144 260104 287156
rect 233200 287116 260104 287144
rect 233200 287104 233206 287116
rect 260098 287104 260104 287116
rect 260156 287104 260162 287156
rect 158806 287036 158812 287088
rect 158864 287076 158870 287088
rect 162118 287076 162124 287088
rect 158864 287048 162124 287076
rect 158864 287036 158870 287048
rect 162118 287036 162124 287048
rect 162176 287036 162182 287088
rect 198734 287036 198740 287088
rect 198792 287076 198798 287088
rect 223574 287076 223580 287088
rect 198792 287048 223580 287076
rect 198792 287036 198798 287048
rect 223574 287036 223580 287048
rect 223632 287036 223638 287088
rect 245838 287036 245844 287088
rect 245896 287076 245902 287088
rect 303614 287076 303620 287088
rect 245896 287048 303620 287076
rect 245896 287036 245902 287048
rect 303614 287036 303620 287048
rect 303672 287036 303678 287088
rect 57606 286968 57612 287020
rect 57664 287008 57670 287020
rect 66806 287008 66812 287020
rect 57664 286980 66812 287008
rect 57664 286968 57670 286980
rect 66806 286968 66812 286980
rect 66864 286968 66870 287020
rect 232682 286968 232688 287020
rect 232740 287008 232746 287020
rect 234246 287008 234252 287020
rect 232740 286980 234252 287008
rect 232740 286968 232746 286980
rect 234246 286968 234252 286980
rect 234304 286968 234310 287020
rect 218606 286628 218612 286680
rect 218664 286668 218670 286680
rect 220078 286668 220084 286680
rect 218664 286640 220084 286668
rect 218664 286628 218670 286640
rect 220078 286628 220084 286640
rect 220136 286628 220142 286680
rect 224218 286356 224224 286408
rect 224276 286396 224282 286408
rect 225046 286396 225052 286408
rect 224276 286368 225052 286396
rect 224276 286356 224282 286368
rect 225046 286356 225052 286368
rect 225104 286356 225110 286408
rect 158806 286288 158812 286340
rect 158864 286328 158870 286340
rect 165062 286328 165068 286340
rect 158864 286300 165068 286328
rect 158864 286288 158870 286300
rect 165062 286288 165068 286300
rect 165120 286288 165126 286340
rect 172054 286288 172060 286340
rect 172112 286328 172118 286340
rect 195330 286328 195336 286340
rect 172112 286300 195336 286328
rect 172112 286288 172118 286300
rect 195330 286288 195336 286300
rect 195388 286288 195394 286340
rect 356698 286084 356704 286136
rect 356756 286124 356762 286136
rect 363598 286124 363604 286136
rect 356756 286096 363604 286124
rect 356756 286084 356762 286096
rect 363598 286084 363604 286096
rect 363656 286084 363662 286136
rect 166442 285948 166448 286000
rect 166500 285988 166506 286000
rect 171870 285988 171876 286000
rect 166500 285960 171876 285988
rect 166500 285948 166506 285960
rect 171870 285948 171876 285960
rect 171928 285948 171934 286000
rect 201402 285812 201408 285864
rect 201460 285852 201466 285864
rect 205542 285852 205548 285864
rect 201460 285824 205548 285852
rect 201460 285812 201466 285824
rect 205542 285812 205548 285824
rect 205600 285812 205606 285864
rect 226536 285824 229094 285852
rect 204990 285744 204996 285796
rect 205048 285784 205054 285796
rect 207014 285784 207020 285796
rect 205048 285756 207020 285784
rect 205048 285744 205054 285756
rect 207014 285744 207020 285756
rect 207072 285744 207078 285796
rect 212902 285744 212908 285796
rect 212960 285784 212966 285796
rect 218054 285784 218060 285796
rect 212960 285756 218060 285784
rect 212960 285744 212966 285756
rect 218054 285744 218060 285756
rect 218112 285744 218118 285796
rect 226536 285728 226564 285824
rect 227622 285744 227628 285796
rect 227680 285784 227686 285796
rect 228910 285784 228916 285796
rect 227680 285756 228916 285784
rect 227680 285744 227686 285756
rect 228910 285744 228916 285756
rect 228968 285744 228974 285796
rect 229066 285784 229094 285824
rect 237374 285784 237380 285796
rect 229066 285756 237380 285784
rect 237374 285744 237380 285756
rect 237432 285744 237438 285796
rect 238478 285744 238484 285796
rect 238536 285784 238542 285796
rect 245010 285784 245016 285796
rect 238536 285756 245016 285784
rect 238536 285744 238542 285756
rect 245010 285744 245016 285756
rect 245068 285744 245074 285796
rect 63402 285676 63408 285728
rect 63460 285716 63466 285728
rect 66254 285716 66260 285728
rect 63460 285688 66260 285716
rect 63460 285676 63466 285688
rect 66254 285676 66260 285688
rect 66312 285676 66318 285728
rect 166350 285676 166356 285728
rect 166408 285716 166414 285728
rect 171962 285716 171968 285728
rect 166408 285688 171968 285716
rect 166408 285676 166414 285688
rect 171962 285676 171968 285688
rect 172020 285676 172026 285728
rect 191098 285676 191104 285728
rect 191156 285716 191162 285728
rect 210878 285716 210884 285728
rect 191156 285688 210884 285716
rect 191156 285676 191162 285688
rect 210878 285676 210884 285688
rect 210936 285676 210942 285728
rect 211798 285676 211804 285728
rect 211856 285716 211862 285728
rect 213822 285716 213828 285728
rect 211856 285688 213828 285716
rect 211856 285676 211862 285688
rect 213822 285676 213828 285688
rect 213880 285676 213886 285728
rect 215202 285676 215208 285728
rect 215260 285716 215266 285728
rect 219158 285716 219164 285728
rect 215260 285688 219164 285716
rect 215260 285676 215266 285688
rect 219158 285676 219164 285688
rect 219216 285676 219222 285728
rect 224310 285676 224316 285728
rect 224368 285716 224374 285728
rect 226518 285716 226524 285728
rect 224368 285688 226524 285716
rect 224368 285676 224374 285688
rect 226518 285676 226524 285688
rect 226576 285676 226582 285728
rect 228358 285676 228364 285728
rect 228416 285716 228422 285728
rect 229278 285716 229284 285728
rect 228416 285688 229284 285716
rect 228416 285676 228422 285688
rect 229278 285676 229284 285688
rect 229336 285676 229342 285728
rect 234430 285676 234436 285728
rect 234488 285716 234494 285728
rect 235166 285716 235172 285728
rect 234488 285688 235172 285716
rect 234488 285676 234494 285688
rect 235166 285676 235172 285688
rect 235224 285676 235230 285728
rect 237558 285676 237564 285728
rect 237616 285716 237622 285728
rect 238570 285716 238576 285728
rect 237616 285688 238576 285716
rect 237616 285676 237622 285688
rect 238570 285676 238576 285688
rect 238628 285676 238634 285728
rect 242342 285676 242348 285728
rect 242400 285716 242406 285728
rect 266998 285716 267004 285728
rect 242400 285688 267004 285716
rect 242400 285676 242406 285688
rect 266998 285676 267004 285688
rect 267056 285676 267062 285728
rect 200114 285268 200120 285320
rect 200172 285308 200178 285320
rect 200942 285308 200948 285320
rect 200172 285280 200948 285308
rect 200172 285268 200178 285280
rect 200942 285268 200948 285280
rect 201000 285268 201006 285320
rect 220814 285268 220820 285320
rect 220872 285308 220878 285320
rect 221274 285308 221280 285320
rect 220872 285280 221280 285308
rect 220872 285268 220878 285280
rect 221274 285268 221280 285280
rect 221332 285268 221338 285320
rect 158162 284928 158168 284980
rect 158220 284968 158226 284980
rect 177574 284968 177580 284980
rect 158220 284940 177580 284968
rect 158220 284928 158226 284940
rect 177574 284928 177580 284940
rect 177632 284928 177638 284980
rect 237466 284928 237472 284980
rect 237524 284968 237530 284980
rect 243906 284968 243912 284980
rect 237524 284940 243912 284968
rect 237524 284928 237530 284940
rect 243906 284928 243912 284940
rect 243964 284928 243970 284980
rect 254670 284928 254676 284980
rect 254728 284968 254734 284980
rect 261570 284968 261576 284980
rect 254728 284940 261576 284968
rect 254728 284928 254734 284940
rect 261570 284928 261576 284940
rect 261628 284928 261634 284980
rect 185670 284384 185676 284436
rect 185728 284424 185734 284436
rect 216766 284424 216772 284436
rect 185728 284396 216772 284424
rect 185728 284384 185734 284396
rect 216766 284384 216772 284396
rect 216824 284384 216830 284436
rect 247034 284384 247040 284436
rect 247092 284424 247098 284436
rect 247678 284424 247684 284436
rect 247092 284396 247684 284424
rect 247092 284384 247098 284396
rect 247678 284384 247684 284396
rect 247736 284424 247742 284436
rect 254578 284424 254584 284436
rect 247736 284396 254584 284424
rect 247736 284384 247742 284396
rect 254578 284384 254584 284396
rect 254636 284384 254642 284436
rect 57882 284316 57888 284368
rect 57940 284356 57946 284368
rect 66806 284356 66812 284368
rect 57940 284328 66812 284356
rect 57940 284316 57946 284328
rect 66806 284316 66812 284328
rect 66864 284316 66870 284368
rect 173250 284316 173256 284368
rect 173308 284356 173314 284368
rect 173308 284328 176700 284356
rect 173308 284316 173314 284328
rect 176672 284288 176700 284328
rect 198734 284316 198740 284368
rect 198792 284356 198798 284368
rect 204622 284356 204628 284368
rect 198792 284328 204628 284356
rect 198792 284316 198798 284328
rect 204622 284316 204628 284328
rect 204680 284316 204686 284368
rect 206646 284316 206652 284368
rect 206704 284356 206710 284368
rect 428458 284356 428464 284368
rect 206704 284328 428464 284356
rect 206704 284316 206710 284328
rect 428458 284316 428464 284328
rect 428516 284316 428522 284368
rect 203334 284288 203340 284300
rect 176672 284260 203340 284288
rect 203334 284248 203340 284260
rect 203392 284248 203398 284300
rect 332594 284248 332600 284300
rect 332652 284288 332658 284300
rect 333882 284288 333888 284300
rect 332652 284260 333888 284288
rect 332652 284248 332658 284260
rect 333882 284248 333888 284260
rect 333940 284288 333946 284300
rect 358170 284288 358176 284300
rect 333940 284260 358176 284288
rect 333940 284248 333946 284260
rect 358170 284248 358176 284260
rect 358228 284248 358234 284300
rect 199470 283908 199476 283960
rect 199528 283948 199534 283960
rect 201402 283948 201408 283960
rect 199528 283920 201408 283948
rect 199528 283908 199534 283920
rect 201402 283908 201408 283920
rect 201460 283908 201466 283960
rect 170582 283568 170588 283620
rect 170640 283608 170646 283620
rect 198826 283608 198832 283620
rect 170640 283580 198832 283608
rect 170640 283568 170646 283580
rect 198826 283568 198832 283580
rect 198884 283568 198890 283620
rect 246298 283568 246304 283620
rect 246356 283608 246362 283620
rect 246850 283608 246856 283620
rect 246356 283580 246856 283608
rect 246356 283568 246362 283580
rect 246850 283568 246856 283580
rect 246908 283608 246914 283620
rect 251174 283608 251180 283620
rect 246908 283580 251180 283608
rect 246908 283568 246914 283580
rect 251174 283568 251180 283580
rect 251232 283568 251238 283620
rect 280982 282956 280988 283008
rect 281040 282996 281046 283008
rect 281718 282996 281724 283008
rect 281040 282968 281724 282996
rect 281040 282956 281046 282968
rect 281718 282956 281724 282968
rect 281776 282956 281782 283008
rect 59170 282888 59176 282940
rect 59228 282928 59234 282940
rect 66806 282928 66812 282940
rect 59228 282900 66812 282928
rect 59228 282888 59234 282900
rect 66806 282888 66812 282900
rect 66864 282888 66870 282940
rect 263594 282888 263600 282940
rect 263652 282928 263658 282940
rect 264882 282928 264888 282940
rect 263652 282900 264888 282928
rect 263652 282888 263658 282900
rect 264882 282888 264888 282900
rect 264940 282928 264946 282940
rect 380158 282928 380164 282940
rect 264940 282900 380164 282928
rect 264940 282888 264946 282900
rect 380158 282888 380164 282900
rect 380216 282888 380222 282940
rect 183278 282820 183284 282872
rect 183336 282860 183342 282872
rect 195146 282860 195152 282872
rect 183336 282832 195152 282860
rect 183336 282820 183342 282832
rect 195146 282820 195152 282832
rect 195204 282820 195210 282872
rect 160094 282140 160100 282192
rect 160152 282180 160158 282192
rect 176654 282180 176660 282192
rect 160152 282152 176660 282180
rect 160152 282140 160158 282152
rect 176654 282140 176660 282152
rect 176712 282140 176718 282192
rect 247494 282140 247500 282192
rect 247552 282180 247558 282192
rect 263594 282180 263600 282192
rect 247552 282152 263600 282180
rect 247552 282140 247558 282152
rect 263594 282140 263600 282152
rect 263652 282140 263658 282192
rect 245930 281664 245936 281716
rect 245988 281704 245994 281716
rect 251082 281704 251088 281716
rect 245988 281676 251088 281704
rect 245988 281664 245994 281676
rect 251082 281664 251088 281676
rect 251140 281664 251146 281716
rect 253198 281664 253204 281716
rect 253256 281704 253262 281716
rect 255498 281704 255504 281716
rect 253256 281676 255504 281704
rect 253256 281664 253262 281676
rect 255498 281664 255504 281676
rect 255556 281664 255562 281716
rect 176654 281528 176660 281580
rect 176712 281568 176718 281580
rect 177942 281568 177948 281580
rect 176712 281540 177948 281568
rect 176712 281528 176718 281540
rect 177942 281528 177948 281540
rect 178000 281568 178006 281580
rect 197354 281568 197360 281580
rect 178000 281540 197360 281568
rect 178000 281528 178006 281540
rect 197354 281528 197360 281540
rect 197412 281528 197418 281580
rect 250622 281460 250628 281512
rect 250680 281500 250686 281512
rect 255498 281500 255504 281512
rect 250680 281472 255504 281500
rect 250680 281460 250686 281472
rect 255498 281460 255504 281472
rect 255556 281460 255562 281512
rect 166534 281392 166540 281444
rect 166592 281432 166598 281444
rect 197354 281432 197360 281444
rect 166592 281404 197360 281432
rect 166592 281392 166598 281404
rect 197354 281392 197360 281404
rect 197412 281392 197418 281444
rect 160830 280780 160836 280832
rect 160888 280820 160894 280832
rect 197170 280820 197176 280832
rect 160888 280792 197176 280820
rect 160888 280780 160894 280792
rect 197170 280780 197176 280792
rect 197228 280820 197234 280832
rect 197446 280820 197452 280832
rect 197228 280792 197452 280820
rect 197228 280780 197234 280792
rect 197446 280780 197452 280792
rect 197504 280780 197510 280832
rect 286410 280780 286416 280832
rect 286468 280820 286474 280832
rect 318058 280820 318064 280832
rect 286468 280792 318064 280820
rect 286468 280780 286474 280792
rect 318058 280780 318064 280792
rect 318116 280780 318122 280832
rect 279050 280576 279056 280628
rect 279108 280616 279114 280628
rect 283558 280616 283564 280628
rect 279108 280588 283564 280616
rect 279108 280576 279114 280588
rect 283558 280576 283564 280588
rect 283616 280576 283622 280628
rect 158806 280236 158812 280288
rect 158864 280276 158870 280288
rect 160922 280276 160928 280288
rect 158864 280248 160928 280276
rect 158864 280236 158870 280248
rect 160922 280236 160928 280248
rect 160980 280236 160986 280288
rect 17862 280168 17868 280220
rect 17920 280208 17926 280220
rect 67542 280208 67548 280220
rect 17920 280180 67548 280208
rect 17920 280168 17926 280180
rect 67542 280168 67548 280180
rect 67600 280168 67606 280220
rect 246114 280168 246120 280220
rect 246172 280208 246178 280220
rect 318794 280208 318800 280220
rect 246172 280180 318800 280208
rect 246172 280168 246178 280180
rect 318794 280168 318800 280180
rect 318852 280168 318858 280220
rect 165522 279760 165528 279812
rect 165580 279800 165586 279812
rect 168558 279800 168564 279812
rect 165580 279772 168564 279800
rect 165580 279760 165586 279772
rect 168558 279760 168564 279772
rect 168616 279760 168622 279812
rect 170398 279488 170404 279540
rect 170456 279528 170462 279540
rect 179414 279528 179420 279540
rect 170456 279500 179420 279528
rect 170456 279488 170462 279500
rect 179414 279488 179420 279500
rect 179472 279488 179478 279540
rect 245930 279488 245936 279540
rect 245988 279528 245994 279540
rect 309778 279528 309784 279540
rect 245988 279500 309784 279528
rect 245988 279488 245994 279500
rect 309778 279488 309784 279500
rect 309836 279488 309842 279540
rect 159358 279420 159364 279472
rect 159416 279460 159422 279472
rect 191834 279460 191840 279472
rect 159416 279432 191840 279460
rect 159416 279420 159422 279432
rect 191834 279420 191840 279432
rect 191892 279420 191898 279472
rect 286318 279420 286324 279472
rect 286376 279460 286382 279472
rect 294598 279460 294604 279472
rect 286376 279432 294604 279460
rect 286376 279420 286382 279432
rect 294598 279420 294604 279432
rect 294656 279420 294662 279472
rect 304258 279420 304264 279472
rect 304316 279460 304322 279472
rect 449894 279460 449900 279472
rect 304316 279432 449900 279460
rect 304316 279420 304322 279432
rect 449894 279420 449900 279432
rect 449952 279420 449958 279472
rect 245930 278944 245936 278996
rect 245988 278984 245994 278996
rect 249150 278984 249156 278996
rect 245988 278956 249156 278984
rect 245988 278944 245994 278956
rect 249150 278944 249156 278956
rect 249208 278944 249214 278996
rect 60274 278740 60280 278792
rect 60332 278780 60338 278792
rect 66622 278780 66628 278792
rect 60332 278752 66628 278780
rect 60332 278740 60338 278752
rect 66622 278740 66628 278752
rect 66680 278740 66686 278792
rect 179414 278740 179420 278792
rect 179472 278780 179478 278792
rect 180702 278780 180708 278792
rect 179472 278752 180708 278780
rect 179472 278740 179478 278752
rect 180702 278740 180708 278752
rect 180760 278780 180766 278792
rect 197354 278780 197360 278792
rect 180760 278752 197360 278780
rect 180760 278740 180766 278752
rect 197354 278740 197360 278752
rect 197412 278740 197418 278792
rect 52178 278672 52184 278724
rect 52236 278712 52242 278724
rect 66806 278712 66812 278724
rect 52236 278684 66812 278712
rect 52236 278672 52242 278684
rect 66806 278672 66812 278684
rect 66864 278672 66870 278724
rect 192662 278672 192668 278724
rect 192720 278712 192726 278724
rect 197170 278712 197176 278724
rect 192720 278684 197176 278712
rect 192720 278672 192726 278684
rect 197170 278672 197176 278684
rect 197228 278712 197234 278724
rect 197446 278712 197452 278724
rect 197228 278684 197452 278712
rect 197228 278672 197234 278684
rect 197446 278672 197452 278684
rect 197504 278672 197510 278724
rect 195882 278604 195888 278656
rect 195940 278644 195946 278656
rect 197354 278644 197360 278656
rect 195940 278616 197360 278644
rect 195940 278604 195946 278616
rect 197354 278604 197360 278616
rect 197412 278604 197418 278656
rect 245930 277992 245936 278044
rect 245988 278032 245994 278044
rect 249886 278032 249892 278044
rect 245988 278004 249892 278032
rect 245988 277992 245994 278004
rect 249886 277992 249892 278004
rect 249944 278032 249950 278044
rect 378226 278032 378232 278044
rect 249944 278004 378232 278032
rect 249944 277992 249950 278004
rect 378226 277992 378232 278004
rect 378284 278032 378290 278044
rect 382918 278032 382924 278044
rect 378284 278004 382924 278032
rect 378284 277992 378290 278004
rect 382918 277992 382924 278004
rect 382976 277992 382982 278044
rect 158622 277380 158628 277432
rect 158680 277420 158686 277432
rect 167638 277420 167644 277432
rect 158680 277392 167644 277420
rect 158680 277380 158686 277392
rect 167638 277380 167644 277392
rect 167696 277380 167702 277432
rect 244366 277380 244372 277432
rect 244424 277420 244430 277432
rect 285030 277420 285036 277432
rect 244424 277392 285036 277420
rect 244424 277380 244430 277392
rect 285030 277380 285036 277392
rect 285088 277380 285094 277432
rect 60550 277312 60556 277364
rect 60608 277352 60614 277364
rect 66254 277352 66260 277364
rect 60608 277324 66260 277352
rect 60608 277312 60614 277324
rect 66254 277312 66260 277324
rect 66312 277312 66318 277364
rect 158806 277312 158812 277364
rect 158864 277352 158870 277364
rect 165154 277352 165160 277364
rect 158864 277324 165160 277352
rect 158864 277312 158870 277324
rect 165154 277312 165160 277324
rect 165212 277312 165218 277364
rect 160922 276632 160928 276684
rect 160980 276672 160986 276684
rect 183278 276672 183284 276684
rect 160980 276644 183284 276672
rect 160980 276632 160986 276644
rect 183278 276632 183284 276644
rect 183336 276632 183342 276684
rect 245746 276632 245752 276684
rect 245804 276672 245810 276684
rect 293954 276672 293960 276684
rect 245804 276644 293960 276672
rect 245804 276632 245810 276644
rect 293954 276632 293960 276644
rect 294012 276672 294018 276684
rect 360194 276672 360200 276684
rect 294012 276644 360200 276672
rect 294012 276632 294018 276644
rect 360194 276632 360200 276644
rect 360252 276632 360258 276684
rect 183278 276088 183284 276140
rect 183336 276128 183342 276140
rect 183336 276100 190454 276128
rect 183336 276088 183342 276100
rect 61838 276020 61844 276072
rect 61896 276060 61902 276072
rect 66806 276060 66812 276072
rect 61896 276032 66812 276060
rect 61896 276020 61902 276032
rect 66806 276020 66812 276032
rect 66864 276020 66870 276072
rect 186222 276020 186228 276072
rect 186280 276060 186286 276072
rect 187234 276060 187240 276072
rect 186280 276032 187240 276060
rect 186280 276020 186286 276032
rect 187234 276020 187240 276032
rect 187292 276020 187298 276072
rect 190426 276060 190454 276100
rect 197446 276060 197452 276072
rect 190426 276032 197452 276060
rect 197446 276020 197452 276032
rect 197504 276020 197510 276072
rect 166902 275952 166908 276004
rect 166960 275992 166966 276004
rect 172514 275992 172520 276004
rect 166960 275964 172520 275992
rect 166960 275952 166966 275964
rect 172514 275952 172520 275964
rect 172572 275992 172578 276004
rect 197262 275992 197268 276004
rect 172572 275964 197268 275992
rect 172572 275952 172578 275964
rect 197262 275952 197268 275964
rect 197320 275992 197326 276004
rect 197538 275992 197544 276004
rect 197320 275964 197544 275992
rect 197320 275952 197326 275964
rect 197538 275952 197544 275964
rect 197596 275952 197602 276004
rect 245930 275952 245936 276004
rect 245988 275992 245994 276004
rect 257338 275992 257344 276004
rect 245988 275964 257344 275992
rect 245988 275952 245994 275964
rect 257338 275952 257344 275964
rect 257396 275952 257402 276004
rect 268378 275952 268384 276004
rect 268436 275992 268442 276004
rect 338850 275992 338856 276004
rect 268436 275964 338856 275992
rect 268436 275952 268442 275964
rect 338850 275952 338856 275964
rect 338908 275952 338914 276004
rect 158806 275884 158812 275936
rect 158864 275924 158870 275936
rect 162210 275924 162216 275936
rect 158864 275896 162216 275924
rect 158864 275884 158870 275896
rect 162210 275884 162216 275896
rect 162268 275884 162274 275936
rect 159818 275272 159824 275324
rect 159876 275312 159882 275324
rect 177390 275312 177396 275324
rect 159876 275284 177396 275312
rect 159876 275272 159882 275284
rect 177390 275272 177396 275284
rect 177448 275272 177454 275324
rect 245930 275272 245936 275324
rect 245988 275312 245994 275324
rect 252830 275312 252836 275324
rect 245988 275284 252836 275312
rect 245988 275272 245994 275284
rect 252830 275272 252836 275284
rect 252888 275272 252894 275324
rect 252830 274660 252836 274712
rect 252888 274700 252894 274712
rect 307110 274700 307116 274712
rect 252888 274672 307116 274700
rect 252888 274660 252894 274672
rect 307110 274660 307116 274672
rect 307168 274660 307174 274712
rect 61930 274592 61936 274644
rect 61988 274632 61994 274644
rect 65886 274632 65892 274644
rect 61988 274604 65892 274632
rect 61988 274592 61994 274604
rect 65886 274592 65892 274604
rect 65944 274592 65950 274644
rect 158806 274592 158812 274644
rect 158864 274632 158870 274644
rect 176102 274632 176108 274644
rect 158864 274604 176108 274632
rect 158864 274592 158870 274604
rect 176102 274592 176108 274604
rect 176160 274592 176166 274644
rect 183462 274524 183468 274576
rect 183520 274564 183526 274576
rect 185026 274564 185032 274576
rect 183520 274536 185032 274564
rect 183520 274524 183526 274536
rect 185026 274524 185032 274536
rect 185084 274524 185090 274576
rect 267182 273980 267188 274032
rect 267240 274020 267246 274032
rect 354122 274020 354128 274032
rect 267240 273992 354128 274020
rect 267240 273980 267246 273992
rect 354122 273980 354128 273992
rect 354180 273980 354186 274032
rect 181714 273912 181720 273964
rect 181772 273952 181778 273964
rect 199470 273952 199476 273964
rect 181772 273924 199476 273952
rect 181772 273912 181778 273924
rect 199470 273912 199476 273924
rect 199528 273912 199534 273964
rect 322198 273912 322204 273964
rect 322256 273952 322262 273964
rect 436738 273952 436744 273964
rect 322256 273924 436744 273952
rect 322256 273912 322262 273924
rect 436738 273912 436744 273924
rect 436796 273912 436802 273964
rect 191834 273436 191840 273488
rect 191892 273476 191898 273488
rect 193030 273476 193036 273488
rect 191892 273448 193036 273476
rect 191892 273436 191898 273448
rect 193030 273436 193036 273448
rect 193088 273476 193094 273488
rect 197446 273476 197452 273488
rect 193088 273448 197452 273476
rect 193088 273436 193094 273448
rect 197446 273436 197452 273448
rect 197504 273436 197510 273488
rect 158806 273232 158812 273284
rect 158864 273272 158870 273284
rect 173342 273272 173348 273284
rect 158864 273244 173348 273272
rect 158864 273232 158870 273244
rect 173342 273232 173348 273244
rect 173400 273232 173406 273284
rect 175090 273164 175096 273216
rect 175148 273204 175154 273216
rect 197446 273204 197452 273216
rect 175148 273176 197452 273204
rect 175148 273164 175154 273176
rect 197446 273164 197452 273176
rect 197504 273164 197510 273216
rect 245838 273164 245844 273216
rect 245896 273204 245902 273216
rect 248598 273204 248604 273216
rect 245896 273176 248604 273204
rect 245896 273164 245902 273176
rect 248598 273164 248604 273176
rect 248656 273204 248662 273216
rect 251266 273204 251272 273216
rect 248656 273176 251272 273204
rect 248656 273164 248662 273176
rect 251266 273164 251272 273176
rect 251324 273164 251330 273216
rect 180242 272484 180248 272536
rect 180300 272524 180306 272536
rect 191374 272524 191380 272536
rect 180300 272496 191380 272524
rect 180300 272484 180306 272496
rect 191374 272484 191380 272496
rect 191432 272484 191438 272536
rect 245930 272484 245936 272536
rect 245988 272524 245994 272536
rect 251266 272524 251272 272536
rect 245988 272496 251272 272524
rect 245988 272484 245994 272496
rect 251266 272484 251272 272496
rect 251324 272524 251330 272536
rect 252462 272524 252468 272536
rect 251324 272496 252468 272524
rect 251324 272484 251330 272496
rect 252462 272484 252468 272496
rect 252520 272484 252526 272536
rect 280890 272484 280896 272536
rect 280948 272524 280954 272536
rect 294598 272524 294604 272536
rect 280948 272496 294604 272524
rect 280948 272484 280954 272496
rect 294598 272484 294604 272496
rect 294656 272484 294662 272536
rect 307662 272484 307668 272536
rect 307720 272524 307726 272536
rect 385034 272524 385040 272536
rect 307720 272496 385040 272524
rect 307720 272484 307726 272496
rect 385034 272484 385040 272496
rect 385092 272484 385098 272536
rect 176102 272280 176108 272332
rect 176160 272320 176166 272332
rect 178678 272320 178684 272332
rect 176160 272292 178684 272320
rect 176160 272280 176166 272292
rect 178678 272280 178684 272292
rect 178736 272280 178742 272332
rect 63126 271872 63132 271924
rect 63184 271912 63190 271924
rect 66254 271912 66260 271924
rect 63184 271884 66260 271912
rect 63184 271872 63190 271884
rect 66254 271872 66260 271884
rect 66312 271872 66318 271924
rect 252462 271872 252468 271924
rect 252520 271912 252526 271924
rect 306374 271912 306380 271924
rect 252520 271884 306380 271912
rect 252520 271872 252526 271884
rect 306374 271872 306380 271884
rect 306432 271912 306438 271924
rect 307662 271912 307668 271924
rect 306432 271884 307668 271912
rect 306432 271872 306438 271884
rect 307662 271872 307668 271884
rect 307720 271872 307726 271924
rect 245930 271192 245936 271244
rect 245988 271232 245994 271244
rect 248598 271232 248604 271244
rect 245988 271204 248604 271232
rect 245988 271192 245994 271204
rect 248598 271192 248604 271204
rect 248656 271192 248662 271244
rect 61930 271124 61936 271176
rect 61988 271164 61994 271176
rect 66898 271164 66904 271176
rect 61988 271136 66904 271164
rect 61988 271124 61994 271136
rect 66898 271124 66904 271136
rect 66956 271124 66962 271176
rect 184750 271124 184756 271176
rect 184808 271164 184814 271176
rect 199562 271164 199568 271176
rect 184808 271136 199568 271164
rect 184808 271124 184814 271136
rect 199562 271124 199568 271136
rect 199620 271124 199626 271176
rect 245838 271124 245844 271176
rect 245896 271164 245902 271176
rect 305178 271164 305184 271176
rect 245896 271136 305184 271164
rect 245896 271124 245902 271136
rect 305178 271124 305184 271136
rect 305236 271164 305242 271176
rect 380894 271164 380900 271176
rect 305236 271136 380900 271164
rect 305236 271124 305242 271136
rect 380894 271124 380900 271136
rect 380952 271124 380958 271176
rect 158806 270784 158812 270836
rect 158864 270824 158870 270836
rect 162210 270824 162216 270836
rect 158864 270796 162216 270824
rect 158864 270784 158870 270796
rect 162210 270784 162216 270796
rect 162268 270784 162274 270836
rect 54938 270512 54944 270564
rect 54996 270552 55002 270564
rect 66898 270552 66904 270564
rect 54996 270524 66904 270552
rect 54996 270512 55002 270524
rect 66898 270512 66904 270524
rect 66956 270512 66962 270564
rect 164142 270512 164148 270564
rect 164200 270552 164206 270564
rect 197446 270552 197452 270564
rect 164200 270524 197452 270552
rect 164200 270512 164206 270524
rect 197446 270512 197452 270524
rect 197504 270512 197510 270564
rect 184382 270444 184388 270496
rect 184440 270484 184446 270496
rect 185762 270484 185768 270496
rect 184440 270456 185768 270484
rect 184440 270444 184446 270456
rect 185762 270444 185768 270456
rect 185820 270444 185826 270496
rect 245930 270172 245936 270224
rect 245988 270212 245994 270224
rect 248506 270212 248512 270224
rect 245988 270184 248512 270212
rect 245988 270172 245994 270184
rect 248506 270172 248512 270184
rect 248564 270172 248570 270224
rect 4062 269764 4068 269816
rect 4120 269804 4126 269816
rect 32398 269804 32404 269816
rect 4120 269776 32404 269804
rect 4120 269764 4126 269776
rect 32398 269764 32404 269776
rect 32456 269764 32462 269816
rect 260098 269764 260104 269816
rect 260156 269804 260162 269816
rect 367738 269804 367744 269816
rect 260156 269776 367744 269804
rect 260156 269764 260162 269776
rect 367738 269764 367744 269776
rect 367796 269764 367802 269816
rect 163682 269084 163688 269136
rect 163740 269124 163746 269136
rect 197446 269124 197452 269136
rect 163740 269096 197452 269124
rect 163740 269084 163746 269096
rect 197446 269084 197452 269096
rect 197504 269084 197510 269136
rect 12434 269016 12440 269068
rect 12492 269056 12498 269068
rect 14458 269056 14464 269068
rect 12492 269028 14464 269056
rect 12492 269016 12498 269028
rect 14458 269016 14464 269028
rect 14516 269016 14522 269068
rect 63310 269016 63316 269068
rect 63368 269056 63374 269068
rect 64782 269056 64788 269068
rect 63368 269028 64788 269056
rect 63368 269016 63374 269028
rect 64782 269016 64788 269028
rect 64840 269016 64846 269068
rect 158806 269016 158812 269068
rect 158864 269056 158870 269068
rect 170582 269056 170588 269068
rect 158864 269028 170588 269056
rect 158864 269016 158870 269028
rect 170582 269016 170588 269028
rect 170640 269016 170646 269068
rect 172422 269016 172428 269068
rect 172480 269056 172486 269068
rect 178678 269056 178684 269068
rect 172480 269028 178684 269056
rect 172480 269016 172486 269028
rect 178678 269016 178684 269028
rect 178736 269016 178742 269068
rect 181530 269016 181536 269068
rect 181588 269056 181594 269068
rect 184290 269056 184296 269068
rect 181588 269028 184296 269056
rect 181588 269016 181594 269028
rect 184290 269016 184296 269028
rect 184348 269016 184354 269068
rect 194410 269016 194416 269068
rect 194468 269056 194474 269068
rect 194686 269056 194692 269068
rect 194468 269028 194692 269056
rect 194468 269016 194474 269028
rect 194686 269016 194692 269028
rect 194744 269016 194750 269068
rect 291838 268948 291844 269000
rect 291896 268988 291902 269000
rect 293218 268988 293224 269000
rect 291896 268960 293224 268988
rect 291896 268948 291902 268960
rect 293218 268948 293224 268960
rect 293276 268948 293282 269000
rect 161290 268336 161296 268388
rect 161348 268376 161354 268388
rect 187326 268376 187332 268388
rect 161348 268348 187332 268376
rect 161348 268336 161354 268348
rect 187326 268336 187332 268348
rect 187384 268336 187390 268388
rect 311986 268336 311992 268388
rect 312044 268376 312050 268388
rect 367186 268376 367192 268388
rect 312044 268348 367192 268376
rect 312044 268336 312050 268348
rect 367186 268336 367192 268348
rect 367244 268336 367250 268388
rect 194686 267996 194692 268048
rect 194744 268036 194750 268048
rect 198274 268036 198280 268048
rect 194744 268008 198280 268036
rect 194744 267996 194750 268008
rect 198274 267996 198280 268008
rect 198332 267996 198338 268048
rect 64782 267860 64788 267912
rect 64840 267900 64846 267912
rect 66806 267900 66812 267912
rect 64840 267872 66812 267900
rect 64840 267860 64846 267872
rect 66806 267860 66812 267872
rect 66864 267860 66870 267912
rect 187326 267724 187332 267776
rect 187384 267764 187390 267776
rect 197538 267764 197544 267776
rect 187384 267736 197544 267764
rect 187384 267724 187390 267736
rect 197538 267724 197544 267736
rect 197596 267724 197602 267776
rect 244458 267724 244464 267776
rect 244516 267764 244522 267776
rect 311986 267764 311992 267776
rect 244516 267736 311992 267764
rect 244516 267724 244522 267736
rect 311986 267724 311992 267736
rect 312044 267724 312050 267776
rect 187602 267656 187608 267708
rect 187660 267696 187666 267708
rect 197446 267696 197452 267708
rect 187660 267668 197452 267696
rect 187660 267656 187666 267668
rect 197446 267656 197452 267668
rect 197504 267656 197510 267708
rect 245746 267656 245752 267708
rect 245804 267696 245810 267708
rect 259638 267696 259644 267708
rect 245804 267668 259644 267696
rect 245804 267656 245810 267668
rect 259638 267656 259644 267668
rect 259696 267656 259702 267708
rect 194318 267112 194324 267164
rect 194376 267152 194382 267164
rect 197538 267152 197544 267164
rect 194376 267124 197544 267152
rect 194376 267112 194382 267124
rect 197538 267112 197544 267124
rect 197596 267112 197602 267164
rect 3142 266976 3148 267028
rect 3200 267016 3206 267028
rect 12434 267016 12440 267028
rect 3200 266988 12440 267016
rect 3200 266976 3206 266988
rect 12434 266976 12440 266988
rect 12492 266976 12498 267028
rect 259638 266976 259644 267028
rect 259696 267016 259702 267028
rect 336090 267016 336096 267028
rect 259696 266988 336096 267016
rect 259696 266976 259702 266988
rect 336090 266976 336096 266988
rect 336148 266976 336154 267028
rect 191282 266908 191288 266960
rect 191340 266948 191346 266960
rect 193214 266948 193220 266960
rect 191340 266920 193220 266948
rect 191340 266908 191346 266920
rect 193214 266908 193220 266920
rect 193272 266908 193278 266960
rect 12434 266364 12440 266416
rect 12492 266404 12498 266416
rect 13078 266404 13084 266416
rect 12492 266376 13084 266404
rect 12492 266364 12498 266376
rect 13078 266364 13084 266376
rect 13136 266364 13142 266416
rect 256786 266364 256792 266416
rect 256844 266364 256850 266416
rect 158806 266296 158812 266348
rect 158864 266336 158870 266348
rect 172054 266336 172060 266348
rect 158864 266308 172060 266336
rect 158864 266296 158870 266308
rect 172054 266296 172060 266308
rect 172112 266296 172118 266348
rect 246022 266296 246028 266348
rect 246080 266336 246086 266348
rect 256804 266336 256832 266364
rect 358170 266336 358176 266348
rect 246080 266308 358176 266336
rect 246080 266296 246086 266308
rect 358170 266296 358176 266308
rect 358228 266336 358234 266348
rect 583294 266336 583300 266348
rect 358228 266308 583300 266336
rect 358228 266296 358234 266308
rect 583294 266296 583300 266308
rect 583352 266296 583358 266348
rect 180610 265684 180616 265736
rect 180668 265724 180674 265736
rect 181438 265724 181444 265736
rect 180668 265696 181444 265724
rect 180668 265684 180674 265696
rect 181438 265684 181444 265696
rect 181496 265684 181502 265736
rect 189810 265684 189816 265736
rect 189868 265724 189874 265736
rect 196618 265724 196624 265736
rect 189868 265696 196624 265724
rect 189868 265684 189874 265696
rect 196618 265684 196624 265696
rect 196676 265684 196682 265736
rect 167730 265616 167736 265668
rect 167788 265656 167794 265668
rect 194318 265656 194324 265668
rect 167788 265628 194324 265656
rect 167788 265616 167794 265628
rect 194318 265616 194324 265628
rect 194376 265616 194382 265668
rect 245838 265616 245844 265668
rect 245896 265656 245902 265668
rect 252554 265656 252560 265668
rect 245896 265628 252560 265656
rect 245896 265616 245902 265628
rect 252554 265616 252560 265628
rect 252612 265616 252618 265668
rect 276750 265616 276756 265668
rect 276808 265656 276814 265668
rect 292574 265656 292580 265668
rect 276808 265628 292580 265656
rect 276808 265616 276814 265628
rect 292574 265616 292580 265628
rect 292632 265616 292638 265668
rect 54846 264936 54852 264988
rect 54904 264976 54910 264988
rect 66806 264976 66812 264988
rect 54904 264948 66812 264976
rect 54904 264936 54910 264948
rect 66806 264936 66812 264948
rect 66864 264936 66870 264988
rect 158806 264868 158812 264920
rect 158864 264908 158870 264920
rect 188522 264908 188528 264920
rect 158864 264880 188528 264908
rect 158864 264868 158870 264880
rect 188522 264868 188528 264880
rect 188580 264868 188586 264920
rect 190362 264868 190368 264920
rect 190420 264908 190426 264920
rect 197446 264908 197452 264920
rect 190420 264880 197452 264908
rect 190420 264868 190426 264880
rect 197446 264868 197452 264880
rect 197504 264868 197510 264920
rect 257430 264256 257436 264308
rect 257488 264296 257494 264308
rect 291194 264296 291200 264308
rect 257488 264268 291200 264296
rect 257488 264256 257494 264268
rect 291194 264256 291200 264268
rect 291252 264256 291258 264308
rect 55122 264188 55128 264240
rect 55180 264228 55186 264240
rect 62114 264228 62120 264240
rect 55180 264200 62120 264228
rect 55180 264188 55186 264200
rect 62114 264188 62120 264200
rect 62172 264188 62178 264240
rect 170582 264188 170588 264240
rect 170640 264228 170646 264240
rect 177298 264228 177304 264240
rect 170640 264200 177304 264228
rect 170640 264188 170646 264200
rect 177298 264188 177304 264200
rect 177356 264188 177362 264240
rect 259362 264188 259368 264240
rect 259420 264228 259426 264240
rect 377490 264228 377496 264240
rect 259420 264200 377496 264228
rect 259420 264188 259426 264200
rect 377490 264188 377496 264200
rect 377548 264188 377554 264240
rect 62114 263576 62120 263628
rect 62172 263616 62178 263628
rect 63218 263616 63224 263628
rect 62172 263588 63224 263616
rect 62172 263576 62178 263588
rect 63218 263576 63224 263588
rect 63276 263616 63282 263628
rect 66898 263616 66904 263628
rect 63276 263588 66904 263616
rect 63276 263576 63282 263588
rect 66898 263576 66904 263588
rect 66956 263576 66962 263628
rect 182082 263576 182088 263628
rect 182140 263616 182146 263628
rect 197446 263616 197452 263628
rect 182140 263588 197452 263616
rect 182140 263576 182146 263588
rect 197446 263576 197452 263588
rect 197504 263576 197510 263628
rect 158806 263508 158812 263560
rect 158864 263548 158870 263560
rect 166258 263548 166264 263560
rect 158864 263520 166264 263548
rect 158864 263508 158870 263520
rect 166258 263508 166264 263520
rect 166316 263508 166322 263560
rect 245010 262964 245016 263016
rect 245068 263004 245074 263016
rect 246390 263004 246396 263016
rect 245068 262976 246396 263004
rect 245068 262964 245074 262976
rect 246390 262964 246396 262976
rect 246448 262964 246454 263016
rect 43990 262828 43996 262880
rect 44048 262868 44054 262880
rect 52454 262868 52460 262880
rect 44048 262840 52460 262868
rect 44048 262828 44054 262840
rect 52454 262828 52460 262840
rect 52512 262828 52518 262880
rect 172422 262828 172428 262880
rect 172480 262868 172486 262880
rect 194686 262868 194692 262880
rect 172480 262840 194692 262868
rect 172480 262828 172486 262840
rect 194686 262828 194692 262840
rect 194744 262828 194750 262880
rect 52454 262216 52460 262268
rect 52512 262256 52518 262268
rect 53558 262256 53564 262268
rect 52512 262228 53564 262256
rect 52512 262216 52518 262228
rect 53558 262216 53564 262228
rect 53616 262256 53622 262268
rect 66806 262256 66812 262268
rect 53616 262228 66812 262256
rect 53616 262216 53622 262228
rect 66806 262216 66812 262228
rect 66864 262216 66870 262268
rect 159450 262216 159456 262268
rect 159508 262256 159514 262268
rect 181438 262256 181444 262268
rect 159508 262228 181444 262256
rect 159508 262216 159514 262228
rect 181438 262216 181444 262228
rect 181496 262256 181502 262268
rect 182082 262256 182088 262268
rect 181496 262228 182088 262256
rect 181496 262216 181502 262228
rect 182082 262216 182088 262228
rect 182140 262216 182146 262268
rect 193122 262216 193128 262268
rect 193180 262256 193186 262268
rect 194778 262256 194784 262268
rect 193180 262228 194784 262256
rect 193180 262216 193186 262228
rect 194778 262216 194784 262228
rect 194836 262256 194842 262268
rect 194836 262228 197308 262256
rect 194836 262216 194842 262228
rect 156782 262148 156788 262200
rect 156840 262188 156846 262200
rect 159542 262188 159548 262200
rect 156840 262160 159548 262188
rect 156840 262148 156846 262160
rect 159542 262148 159548 262160
rect 159600 262148 159606 262200
rect 178770 262188 178776 262200
rect 161446 262160 178776 262188
rect 158622 262080 158628 262132
rect 158680 262120 158686 262132
rect 161446 262120 161474 262160
rect 178770 262148 178776 262160
rect 178828 262148 178834 262200
rect 197280 262188 197308 262228
rect 245838 262216 245844 262268
rect 245896 262256 245902 262268
rect 248506 262256 248512 262268
rect 245896 262228 248512 262256
rect 245896 262216 245902 262228
rect 248506 262216 248512 262228
rect 248564 262216 248570 262268
rect 258902 262216 258908 262268
rect 258960 262256 258966 262268
rect 356790 262256 356796 262268
rect 258960 262228 356796 262256
rect 258960 262216 258966 262228
rect 356790 262216 356796 262228
rect 356848 262216 356854 262268
rect 198090 262188 198096 262200
rect 197280 262160 198096 262188
rect 198090 262148 198096 262160
rect 198148 262148 198154 262200
rect 158680 262092 161474 262120
rect 158680 262080 158686 262092
rect 254578 261536 254584 261588
rect 254636 261576 254642 261588
rect 300118 261576 300124 261588
rect 254636 261548 300124 261576
rect 254636 261536 254642 261548
rect 300118 261536 300124 261548
rect 300176 261536 300182 261588
rect 32398 261468 32404 261520
rect 32456 261508 32462 261520
rect 51074 261508 51080 261520
rect 32456 261480 51080 261508
rect 32456 261468 32462 261480
rect 51074 261468 51080 261480
rect 51132 261468 51138 261520
rect 188430 261468 188436 261520
rect 188488 261508 188494 261520
rect 196802 261508 196808 261520
rect 188488 261480 196808 261508
rect 188488 261468 188494 261480
rect 196802 261468 196808 261480
rect 196860 261468 196866 261520
rect 57606 260924 57612 260976
rect 57664 260964 57670 260976
rect 66806 260964 66812 260976
rect 57664 260936 66812 260964
rect 57664 260924 57670 260936
rect 66806 260924 66812 260936
rect 66864 260924 66870 260976
rect 51074 260856 51080 260908
rect 51132 260896 51138 260908
rect 52178 260896 52184 260908
rect 51132 260868 52184 260896
rect 51132 260856 51138 260868
rect 52178 260856 52184 260868
rect 52236 260896 52242 260908
rect 66254 260896 66260 260908
rect 52236 260868 66260 260896
rect 52236 260856 52242 260868
rect 66254 260856 66260 260868
rect 66312 260856 66318 260908
rect 167086 260856 167092 260908
rect 167144 260896 167150 260908
rect 197446 260896 197452 260908
rect 167144 260868 197452 260896
rect 167144 260856 167150 260868
rect 197446 260856 197452 260868
rect 197504 260856 197510 260908
rect 246022 260788 246028 260840
rect 246080 260828 246086 260840
rect 255498 260828 255504 260840
rect 246080 260800 255504 260828
rect 246080 260788 246086 260800
rect 255498 260788 255504 260800
rect 255556 260828 255562 260840
rect 317322 260828 317328 260840
rect 255556 260800 317328 260828
rect 255556 260788 255562 260800
rect 317322 260788 317328 260800
rect 317380 260828 317386 260840
rect 318058 260828 318064 260840
rect 317380 260800 318064 260828
rect 317380 260788 317386 260800
rect 318058 260788 318064 260800
rect 318116 260788 318122 260840
rect 157978 260108 157984 260160
rect 158036 260148 158042 260160
rect 191282 260148 191288 260160
rect 158036 260120 191288 260148
rect 158036 260108 158042 260120
rect 191282 260108 191288 260120
rect 191340 260108 191346 260160
rect 303706 260108 303712 260160
rect 303764 260148 303770 260160
rect 373994 260148 374000 260160
rect 303764 260120 374000 260148
rect 303764 260108 303770 260120
rect 373994 260108 374000 260120
rect 374052 260108 374058 260160
rect 158898 259428 158904 259480
rect 158956 259468 158962 259480
rect 166258 259468 166264 259480
rect 158956 259440 166264 259468
rect 158956 259428 158962 259440
rect 166258 259428 166264 259440
rect 166316 259428 166322 259480
rect 188430 259428 188436 259480
rect 188488 259468 188494 259480
rect 197446 259468 197452 259480
rect 188488 259440 197452 259468
rect 188488 259428 188494 259440
rect 197446 259428 197452 259440
rect 197504 259428 197510 259480
rect 245654 259428 245660 259480
rect 245712 259468 245718 259480
rect 303706 259468 303712 259480
rect 245712 259440 303712 259468
rect 245712 259428 245718 259440
rect 303706 259428 303712 259440
rect 303764 259428 303770 259480
rect 182082 259360 182088 259412
rect 182140 259400 182146 259412
rect 185670 259400 185676 259412
rect 182140 259372 185676 259400
rect 182140 259360 182146 259372
rect 185670 259360 185676 259372
rect 185728 259360 185734 259412
rect 245838 259360 245844 259412
rect 245896 259400 245902 259412
rect 260926 259400 260932 259412
rect 245896 259372 260932 259400
rect 245896 259360 245902 259372
rect 260926 259360 260932 259372
rect 260984 259400 260990 259412
rect 262122 259400 262128 259412
rect 260984 259372 262128 259400
rect 260984 259360 260990 259372
rect 262122 259360 262128 259372
rect 262180 259360 262186 259412
rect 262122 258748 262128 258800
rect 262180 258788 262186 258800
rect 292758 258788 292764 258800
rect 262180 258760 292764 258788
rect 262180 258748 262186 258760
rect 292758 258748 292764 258760
rect 292816 258788 292822 258800
rect 361666 258788 361672 258800
rect 292816 258760 361672 258788
rect 292816 258748 292822 258760
rect 361666 258748 361672 258760
rect 361724 258748 361730 258800
rect 165062 258680 165068 258732
rect 165120 258720 165126 258732
rect 174722 258720 174728 258732
rect 165120 258692 174728 258720
rect 165120 258680 165126 258692
rect 174722 258680 174728 258692
rect 174780 258680 174786 258732
rect 288526 258680 288532 258732
rect 288584 258720 288590 258732
rect 369946 258720 369952 258732
rect 288584 258692 369952 258720
rect 288584 258680 288590 258692
rect 369946 258680 369952 258692
rect 370004 258680 370010 258732
rect 175090 258544 175096 258596
rect 175148 258584 175154 258596
rect 176102 258584 176108 258596
rect 175148 258556 176108 258584
rect 175148 258544 175154 258556
rect 176102 258544 176108 258556
rect 176160 258544 176166 258596
rect 191834 258476 191840 258528
rect 191892 258516 191898 258528
rect 197446 258516 197452 258528
rect 191892 258488 197452 258516
rect 191892 258476 191898 258488
rect 197446 258476 197452 258488
rect 197504 258476 197510 258528
rect 182082 258176 182088 258188
rect 161446 258148 182088 258176
rect 66254 258108 66260 258120
rect 62040 258080 66260 258108
rect 34422 258000 34428 258052
rect 34480 258040 34486 258052
rect 61378 258040 61384 258052
rect 34480 258012 61384 258040
rect 34480 258000 34486 258012
rect 61378 258000 61384 258012
rect 61436 258040 61442 258052
rect 62040 258040 62068 258080
rect 66254 258068 66260 258080
rect 66312 258068 66318 258120
rect 158806 258068 158812 258120
rect 158864 258108 158870 258120
rect 161446 258108 161474 258148
rect 182082 258136 182088 258148
rect 182140 258136 182146 258188
rect 189718 258136 189724 258188
rect 189776 258176 189782 258188
rect 191834 258176 191840 258188
rect 189776 258148 191840 258176
rect 189776 258136 189782 258148
rect 191834 258136 191840 258148
rect 191892 258136 191898 258188
rect 158864 258080 161474 258108
rect 158864 258068 158870 258080
rect 185578 258068 185584 258120
rect 185636 258108 185642 258120
rect 191098 258108 191104 258120
rect 185636 258080 191104 258108
rect 185636 258068 185642 258080
rect 191098 258068 191104 258080
rect 191156 258068 191162 258120
rect 245654 258068 245660 258120
rect 245712 258108 245718 258120
rect 288526 258108 288532 258120
rect 245712 258080 288532 258108
rect 245712 258068 245718 258080
rect 288526 258068 288532 258080
rect 288584 258068 288590 258120
rect 61436 258012 62068 258040
rect 61436 258000 61442 258012
rect 245838 258000 245844 258052
rect 245896 258040 245902 258052
rect 256694 258040 256700 258052
rect 245896 258012 256700 258040
rect 245896 258000 245902 258012
rect 256694 258000 256700 258012
rect 256752 258000 256758 258052
rect 273898 257388 273904 257440
rect 273956 257428 273962 257440
rect 348418 257428 348424 257440
rect 273956 257400 348424 257428
rect 273956 257388 273962 257400
rect 348418 257388 348424 257400
rect 348476 257388 348482 257440
rect 162210 257320 162216 257372
rect 162268 257360 162274 257372
rect 184198 257360 184204 257372
rect 162268 257332 184204 257360
rect 162268 257320 162274 257332
rect 184198 257320 184204 257332
rect 184256 257320 184262 257372
rect 250530 257320 250536 257372
rect 250588 257360 250594 257372
rect 441614 257360 441620 257372
rect 250588 257332 441620 257360
rect 250588 257320 250594 257332
rect 441614 257320 441620 257332
rect 441672 257320 441678 257372
rect 159266 257048 159272 257100
rect 159324 257088 159330 257100
rect 160830 257088 160836 257100
rect 159324 257060 160836 257088
rect 159324 257048 159330 257060
rect 160830 257048 160836 257060
rect 160888 257048 160894 257100
rect 189718 256776 189724 256828
rect 189776 256816 189782 256828
rect 197446 256816 197452 256828
rect 189776 256788 197452 256816
rect 189776 256776 189782 256788
rect 197446 256776 197452 256788
rect 197504 256776 197510 256828
rect 64506 256708 64512 256760
rect 64564 256748 64570 256760
rect 66898 256748 66904 256760
rect 64564 256720 66904 256748
rect 64564 256708 64570 256720
rect 66898 256708 66904 256720
rect 66956 256708 66962 256760
rect 184198 256708 184204 256760
rect 184256 256748 184262 256760
rect 184658 256748 184664 256760
rect 184256 256720 184664 256748
rect 184256 256708 184262 256720
rect 184658 256708 184664 256720
rect 184716 256748 184722 256760
rect 197538 256748 197544 256760
rect 184716 256720 197544 256748
rect 184716 256708 184722 256720
rect 197538 256708 197544 256720
rect 197596 256708 197602 256760
rect 256694 256708 256700 256760
rect 256752 256748 256758 256760
rect 260098 256748 260104 256760
rect 256752 256720 260104 256748
rect 256752 256708 256758 256720
rect 260098 256708 260104 256720
rect 260156 256708 260162 256760
rect 178034 256640 178040 256692
rect 178092 256680 178098 256692
rect 179322 256680 179328 256692
rect 178092 256652 179328 256680
rect 178092 256640 178098 256652
rect 179322 256640 179328 256652
rect 179380 256680 179386 256692
rect 197446 256680 197452 256692
rect 179380 256652 197452 256680
rect 179380 256640 179386 256652
rect 197446 256640 197452 256652
rect 197504 256640 197510 256692
rect 245838 256640 245844 256692
rect 245896 256680 245902 256692
rect 254118 256680 254124 256692
rect 245896 256652 254124 256680
rect 245896 256640 245902 256652
rect 254118 256640 254124 256652
rect 254176 256640 254182 256692
rect 245838 256028 245844 256080
rect 245896 256068 245902 256080
rect 258166 256068 258172 256080
rect 245896 256040 258172 256068
rect 245896 256028 245902 256040
rect 258166 256028 258172 256040
rect 258224 256028 258230 256080
rect 162210 255960 162216 256012
rect 162268 256000 162274 256012
rect 178034 256000 178040 256012
rect 162268 255972 178040 256000
rect 162268 255960 162274 255972
rect 178034 255960 178040 255972
rect 178092 255960 178098 256012
rect 254118 255960 254124 256012
rect 254176 256000 254182 256012
rect 309226 256000 309232 256012
rect 254176 255972 309232 256000
rect 254176 255960 254182 255972
rect 309226 255960 309232 255972
rect 309284 256000 309290 256012
rect 363138 256000 363144 256012
rect 309284 255972 363144 256000
rect 309284 255960 309290 255972
rect 363138 255960 363144 255972
rect 363196 255960 363202 256012
rect 60458 255280 60464 255332
rect 60516 255320 60522 255332
rect 66806 255320 66812 255332
rect 60516 255292 66812 255320
rect 60516 255280 60522 255292
rect 66806 255280 66812 255292
rect 66864 255280 66870 255332
rect 158806 255280 158812 255332
rect 158864 255320 158870 255332
rect 173802 255320 173808 255332
rect 158864 255292 173808 255320
rect 158864 255280 158870 255292
rect 173802 255280 173808 255292
rect 173860 255280 173866 255332
rect 257522 255280 257528 255332
rect 257580 255320 257586 255332
rect 300854 255320 300860 255332
rect 257580 255292 300860 255320
rect 257580 255280 257586 255292
rect 300854 255280 300860 255292
rect 300912 255280 300918 255332
rect 194410 255212 194416 255264
rect 194468 255252 194474 255264
rect 197446 255252 197452 255264
rect 194468 255224 197452 255252
rect 194468 255212 194474 255224
rect 197446 255212 197452 255224
rect 197504 255212 197510 255264
rect 246022 255212 246028 255264
rect 246080 255252 246086 255264
rect 251358 255252 251364 255264
rect 246080 255224 251364 255252
rect 246080 255212 246086 255224
rect 251358 255212 251364 255224
rect 251416 255252 251422 255264
rect 252462 255252 252468 255264
rect 251416 255224 252468 255252
rect 251416 255212 251422 255224
rect 252462 255212 252468 255224
rect 252520 255212 252526 255264
rect 245838 255144 245844 255196
rect 245896 255184 245902 255196
rect 247310 255184 247316 255196
rect 245896 255156 247316 255184
rect 245896 255144 245902 255156
rect 247310 255144 247316 255156
rect 247368 255144 247374 255196
rect 252462 254600 252468 254652
rect 252520 254640 252526 254652
rect 322198 254640 322204 254652
rect 252520 254612 322204 254640
rect 252520 254600 252526 254612
rect 322198 254600 322204 254612
rect 322256 254600 322262 254652
rect 158806 254532 158812 254584
rect 158864 254572 158870 254584
rect 189718 254572 189724 254584
rect 158864 254544 189724 254572
rect 158864 254532 158870 254544
rect 189718 254532 189724 254544
rect 189776 254532 189782 254584
rect 258166 254532 258172 254584
rect 258224 254572 258230 254584
rect 384298 254572 384304 254584
rect 258224 254544 384304 254572
rect 258224 254532 258230 254544
rect 384298 254532 384304 254544
rect 384356 254532 384362 254584
rect 3142 253920 3148 253972
rect 3200 253960 3206 253972
rect 10962 253960 10968 253972
rect 3200 253932 10968 253960
rect 3200 253920 3206 253932
rect 10962 253920 10968 253932
rect 11020 253960 11026 253972
rect 11698 253960 11704 253972
rect 11020 253932 11704 253960
rect 11020 253920 11026 253932
rect 11698 253920 11704 253932
rect 11756 253920 11762 253972
rect 63310 253920 63316 253972
rect 63368 253960 63374 253972
rect 66806 253960 66812 253972
rect 63368 253932 66812 253960
rect 63368 253920 63374 253932
rect 66806 253920 66812 253932
rect 66864 253920 66870 253972
rect 158898 253920 158904 253972
rect 158956 253960 158962 253972
rect 162762 253960 162768 253972
rect 158956 253932 162768 253960
rect 158956 253920 158962 253932
rect 162762 253920 162768 253932
rect 162820 253920 162826 253972
rect 247034 253920 247040 253972
rect 247092 253960 247098 253972
rect 247310 253960 247316 253972
rect 247092 253932 247316 253960
rect 247092 253920 247098 253932
rect 247310 253920 247316 253932
rect 247368 253920 247374 253972
rect 246022 253852 246028 253904
rect 246080 253892 246086 253904
rect 267826 253892 267832 253904
rect 246080 253864 267832 253892
rect 246080 253852 246086 253864
rect 267826 253852 267832 253864
rect 267884 253892 267890 253904
rect 269022 253892 269028 253904
rect 267884 253864 269028 253892
rect 267884 253852 267890 253864
rect 269022 253852 269028 253864
rect 269080 253852 269086 253904
rect 314654 253240 314660 253292
rect 314712 253280 314718 253292
rect 358998 253280 359004 253292
rect 314712 253252 359004 253280
rect 314712 253240 314718 253252
rect 358998 253240 359004 253252
rect 359056 253240 359062 253292
rect 39942 253172 39948 253224
rect 40000 253212 40006 253224
rect 60090 253212 60096 253224
rect 40000 253184 60096 253212
rect 40000 253172 40006 253184
rect 60090 253172 60096 253184
rect 60148 253172 60154 253224
rect 185762 253172 185768 253224
rect 185820 253212 185826 253224
rect 197906 253212 197912 253224
rect 185820 253184 197912 253212
rect 185820 253172 185826 253184
rect 197906 253172 197912 253184
rect 197964 253212 197970 253224
rect 198366 253212 198372 253224
rect 197964 253184 198372 253212
rect 197964 253172 197970 253184
rect 198366 253172 198372 253184
rect 198424 253172 198430 253224
rect 269022 253172 269028 253224
rect 269080 253212 269086 253224
rect 300946 253212 300952 253224
rect 269080 253184 300952 253212
rect 269080 253172 269086 253184
rect 300946 253172 300952 253184
rect 301004 253212 301010 253224
rect 372614 253212 372620 253224
rect 301004 253184 372620 253212
rect 301004 253172 301010 253184
rect 372614 253172 372620 253184
rect 372672 253172 372678 253224
rect 158806 252628 158812 252680
rect 158864 252668 158870 252680
rect 176102 252668 176108 252680
rect 158864 252640 176108 252668
rect 158864 252628 158870 252640
rect 176102 252628 176108 252640
rect 176160 252628 176166 252680
rect 60090 252560 60096 252612
rect 60148 252600 60154 252612
rect 60366 252600 60372 252612
rect 60148 252572 60372 252600
rect 60148 252560 60154 252572
rect 60366 252560 60372 252572
rect 60424 252600 60430 252612
rect 66806 252600 66812 252612
rect 60424 252572 66812 252600
rect 60424 252560 60430 252572
rect 66806 252560 66812 252572
rect 66864 252560 66870 252612
rect 159634 252560 159640 252612
rect 159692 252600 159698 252612
rect 195882 252600 195888 252612
rect 159692 252572 195888 252600
rect 159692 252560 159698 252572
rect 195882 252560 195888 252572
rect 195940 252600 195946 252612
rect 197446 252600 197452 252612
rect 195940 252572 197452 252600
rect 195940 252560 195946 252572
rect 197446 252560 197452 252572
rect 197504 252560 197510 252612
rect 245654 252560 245660 252612
rect 245712 252600 245718 252612
rect 314654 252600 314660 252612
rect 245712 252572 314660 252600
rect 245712 252560 245718 252572
rect 314654 252560 314660 252572
rect 314712 252560 314718 252612
rect 246022 252492 246028 252544
rect 246080 252532 246086 252544
rect 263686 252532 263692 252544
rect 246080 252504 263692 252532
rect 246080 252492 246086 252504
rect 263686 252492 263692 252504
rect 263744 252492 263750 252544
rect 245838 252220 245844 252272
rect 245896 252260 245902 252272
rect 249794 252260 249800 252272
rect 245896 252232 249800 252260
rect 245896 252220 245902 252232
rect 249794 252220 249800 252232
rect 249852 252260 249858 252272
rect 251082 252260 251088 252272
rect 249852 252232 251088 252260
rect 249852 252220 249858 252232
rect 251082 252220 251088 252232
rect 251140 252220 251146 252272
rect 173434 251988 173440 252000
rect 161446 251960 173440 251988
rect 159358 251880 159364 251932
rect 159416 251920 159422 251932
rect 161446 251920 161474 251960
rect 173434 251948 173440 251960
rect 173492 251948 173498 252000
rect 159416 251892 161474 251920
rect 159416 251880 159422 251892
rect 173802 251880 173808 251932
rect 173860 251920 173866 251932
rect 194318 251920 194324 251932
rect 173860 251892 194324 251920
rect 173860 251880 173866 251892
rect 194318 251880 194324 251892
rect 194376 251880 194382 251932
rect 291102 251880 291108 251932
rect 291160 251920 291166 251932
rect 302234 251920 302240 251932
rect 291160 251892 302240 251920
rect 291160 251880 291166 251892
rect 302234 251880 302240 251892
rect 302292 251880 302298 251932
rect 309870 251880 309876 251932
rect 309928 251920 309934 251932
rect 345658 251920 345664 251932
rect 309928 251892 345664 251920
rect 309928 251880 309934 251892
rect 345658 251880 345664 251892
rect 345716 251880 345722 251932
rect 162762 251812 162768 251864
rect 162820 251852 162826 251864
rect 183278 251852 183284 251864
rect 162820 251824 183284 251852
rect 162820 251812 162826 251824
rect 183278 251812 183284 251824
rect 183336 251852 183342 251864
rect 183554 251852 183560 251864
rect 183336 251824 183560 251852
rect 183336 251812 183342 251824
rect 183554 251812 183560 251824
rect 183612 251812 183618 251864
rect 263686 251812 263692 251864
rect 263744 251852 263750 251864
rect 460934 251852 460940 251864
rect 263744 251824 460940 251852
rect 263744 251812 263750 251824
rect 460934 251812 460940 251824
rect 460992 251812 460998 251864
rect 65886 251744 65892 251796
rect 65944 251784 65950 251796
rect 66990 251784 66996 251796
rect 65944 251756 66996 251784
rect 65944 251744 65950 251756
rect 66990 251744 66996 251756
rect 67048 251744 67054 251796
rect 194318 251608 194324 251660
rect 194376 251648 194382 251660
rect 197078 251648 197084 251660
rect 194376 251620 197084 251648
rect 194376 251608 194382 251620
rect 197078 251608 197084 251620
rect 197136 251608 197142 251660
rect 191374 251200 191380 251252
rect 191432 251240 191438 251252
rect 193122 251240 193128 251252
rect 191432 251212 193128 251240
rect 191432 251200 191438 251212
rect 193122 251200 193128 251212
rect 193180 251200 193186 251252
rect 158806 251132 158812 251184
rect 158864 251172 158870 251184
rect 166350 251172 166356 251184
rect 158864 251144 166356 251172
rect 158864 251132 158870 251144
rect 166350 251132 166356 251144
rect 166408 251132 166414 251184
rect 307754 250520 307760 250572
rect 307812 250560 307818 250572
rect 356054 250560 356060 250572
rect 307812 250532 356060 250560
rect 307812 250520 307818 250532
rect 356054 250520 356060 250532
rect 356112 250520 356118 250572
rect 160922 250452 160928 250504
rect 160980 250492 160986 250504
rect 167730 250492 167736 250504
rect 160980 250464 167736 250492
rect 160980 250452 160986 250464
rect 167730 250452 167736 250464
rect 167788 250452 167794 250504
rect 173342 250452 173348 250504
rect 173400 250492 173406 250504
rect 191742 250492 191748 250504
rect 173400 250464 191748 250492
rect 173400 250452 173406 250464
rect 191742 250452 191748 250464
rect 191800 250452 191806 250504
rect 317322 250452 317328 250504
rect 317380 250492 317386 250504
rect 368474 250492 368480 250504
rect 317380 250464 368480 250492
rect 317380 250452 317386 250464
rect 368474 250452 368480 250464
rect 368532 250452 368538 250504
rect 252462 249840 252468 249892
rect 252520 249880 252526 249892
rect 285122 249880 285128 249892
rect 252520 249852 285128 249880
rect 252520 249840 252526 249852
rect 285122 249840 285128 249852
rect 285180 249840 285186 249892
rect 191098 249772 191104 249824
rect 191156 249812 191162 249824
rect 197446 249812 197452 249824
rect 191156 249784 197452 249812
rect 191156 249772 191162 249784
rect 197446 249772 197452 249784
rect 197504 249772 197510 249824
rect 247310 249772 247316 249824
rect 247368 249812 247374 249824
rect 316034 249812 316040 249824
rect 247368 249784 316040 249812
rect 247368 249772 247374 249784
rect 316034 249772 316040 249784
rect 316092 249812 316098 249824
rect 317322 249812 317328 249824
rect 316092 249784 317328 249812
rect 316092 249772 316098 249784
rect 317322 249772 317328 249784
rect 317380 249772 317386 249824
rect 246022 249704 246028 249756
rect 246080 249744 246086 249756
rect 251818 249744 251824 249756
rect 246080 249716 251824 249744
rect 246080 249704 246086 249716
rect 251818 249704 251824 249716
rect 251876 249744 251882 249756
rect 252462 249744 252468 249756
rect 251876 249716 252468 249744
rect 251876 249704 251882 249716
rect 252462 249704 252468 249716
rect 252520 249704 252526 249756
rect 191742 249500 191748 249552
rect 191800 249540 191806 249552
rect 197446 249540 197452 249552
rect 191800 249512 197452 249540
rect 191800 249500 191806 249512
rect 197446 249500 197452 249512
rect 197504 249500 197510 249552
rect 181530 249364 181536 249416
rect 181588 249404 181594 249416
rect 189810 249404 189816 249416
rect 181588 249376 189816 249404
rect 181588 249364 181594 249376
rect 189810 249364 189816 249376
rect 189868 249364 189874 249416
rect 284938 249092 284944 249144
rect 284996 249132 285002 249144
rect 307846 249132 307852 249144
rect 284996 249104 307852 249132
rect 284996 249092 285002 249104
rect 307846 249092 307852 249104
rect 307904 249092 307910 249144
rect 265710 249024 265716 249076
rect 265768 249064 265774 249076
rect 429838 249064 429844 249076
rect 265768 249036 429844 249064
rect 265768 249024 265774 249036
rect 429838 249024 429844 249036
rect 429896 249024 429902 249076
rect 193122 248684 193128 248736
rect 193180 248724 193186 248736
rect 197446 248724 197452 248736
rect 193180 248696 197452 248724
rect 193180 248684 193186 248696
rect 197446 248684 197452 248696
rect 197504 248684 197510 248736
rect 175918 248480 175924 248532
rect 175976 248520 175982 248532
rect 181714 248520 181720 248532
rect 175976 248492 181720 248520
rect 175976 248480 175982 248492
rect 181714 248480 181720 248492
rect 181772 248480 181778 248532
rect 67542 248412 67548 248464
rect 67600 248452 67606 248464
rect 67910 248452 67916 248464
rect 67600 248424 67916 248452
rect 67600 248412 67606 248424
rect 67910 248412 67916 248424
rect 67968 248412 67974 248464
rect 158806 248412 158812 248464
rect 158864 248452 158870 248464
rect 187142 248452 187148 248464
rect 158864 248424 187148 248452
rect 158864 248412 158870 248424
rect 187142 248412 187148 248424
rect 187200 248412 187206 248464
rect 67542 248276 67548 248328
rect 67600 248316 67606 248328
rect 67910 248316 67916 248328
rect 67600 248288 67916 248316
rect 67600 248276 67606 248288
rect 67910 248276 67916 248288
rect 67968 248276 67974 248328
rect 196710 247160 196716 247172
rect 180766 247132 196716 247160
rect 159542 247052 159548 247104
rect 159600 247092 159606 247104
rect 180766 247092 180794 247132
rect 196710 247120 196716 247132
rect 196768 247160 196774 247172
rect 197262 247160 197268 247172
rect 196768 247132 197268 247160
rect 196768 247120 196774 247132
rect 197262 247120 197268 247132
rect 197320 247120 197326 247172
rect 159600 247064 180794 247092
rect 159600 247052 159606 247064
rect 195330 247052 195336 247104
rect 195388 247092 195394 247104
rect 197722 247092 197728 247104
rect 195388 247064 197728 247092
rect 195388 247052 195394 247064
rect 197722 247052 197728 247064
rect 197780 247052 197786 247104
rect 245010 247052 245016 247104
rect 245068 247092 245074 247104
rect 245654 247092 245660 247104
rect 245068 247064 245660 247092
rect 245068 247052 245074 247064
rect 245654 247052 245660 247064
rect 245712 247052 245718 247104
rect 245838 247052 245844 247104
rect 245896 247092 245902 247104
rect 267826 247092 267832 247104
rect 245896 247064 267832 247092
rect 245896 247052 245902 247064
rect 267826 247052 267832 247064
rect 267884 247052 267890 247104
rect 60642 246984 60648 247036
rect 60700 247024 60706 247036
rect 66806 247024 66812 247036
rect 60700 246996 66812 247024
rect 60700 246984 60706 246996
rect 66806 246984 66812 246996
rect 66864 246984 66870 247036
rect 158806 246372 158812 246424
rect 158864 246412 158870 246424
rect 176194 246412 176200 246424
rect 158864 246384 176200 246412
rect 158864 246372 158870 246384
rect 176194 246372 176200 246384
rect 176252 246412 176258 246424
rect 184198 246412 184204 246424
rect 176252 246384 184204 246412
rect 176252 246372 176258 246384
rect 184198 246372 184204 246384
rect 184256 246372 184262 246424
rect 245654 246372 245660 246424
rect 245712 246412 245718 246424
rect 253106 246412 253112 246424
rect 245712 246384 253112 246412
rect 245712 246372 245718 246384
rect 253106 246372 253112 246384
rect 253164 246372 253170 246424
rect 257338 246372 257344 246424
rect 257396 246412 257402 246424
rect 269114 246412 269120 246424
rect 257396 246384 269120 246412
rect 257396 246372 257402 246384
rect 269114 246372 269120 246384
rect 269172 246372 269178 246424
rect 274082 246372 274088 246424
rect 274140 246412 274146 246424
rect 291194 246412 291200 246424
rect 274140 246384 291200 246412
rect 274140 246372 274146 246384
rect 291194 246372 291200 246384
rect 291252 246372 291258 246424
rect 162118 246304 162124 246356
rect 162176 246344 162182 246356
rect 199470 246344 199476 246356
rect 162176 246316 199476 246344
rect 162176 246304 162182 246316
rect 199470 246304 199476 246316
rect 199528 246304 199534 246356
rect 246298 246304 246304 246356
rect 246356 246344 246362 246356
rect 283558 246344 283564 246356
rect 246356 246316 283564 246344
rect 246356 246304 246362 246316
rect 283558 246304 283564 246316
rect 283616 246304 283622 246356
rect 64598 245624 64604 245676
rect 64656 245664 64662 245676
rect 66806 245664 66812 245676
rect 64656 245636 66812 245664
rect 64656 245624 64662 245636
rect 66806 245624 66812 245636
rect 66864 245624 66870 245676
rect 194226 245624 194232 245676
rect 194284 245664 194290 245676
rect 194594 245664 194600 245676
rect 194284 245636 194600 245664
rect 194284 245624 194290 245636
rect 194594 245624 194600 245636
rect 194652 245624 194658 245676
rect 48130 245556 48136 245608
rect 48188 245596 48194 245608
rect 66898 245596 66904 245608
rect 48188 245568 66904 245596
rect 48188 245556 48194 245568
rect 66898 245556 66904 245568
rect 66956 245556 66962 245608
rect 180518 245556 180524 245608
rect 180576 245596 180582 245608
rect 181622 245596 181628 245608
rect 180576 245568 181628 245596
rect 180576 245556 180582 245568
rect 181622 245556 181628 245568
rect 181680 245556 181686 245608
rect 260742 244944 260748 244996
rect 260800 244984 260806 244996
rect 313274 244984 313280 244996
rect 260800 244956 313280 244984
rect 260800 244944 260806 244956
rect 313274 244944 313280 244956
rect 313332 244984 313338 244996
rect 352650 244984 352656 244996
rect 313332 244956 352656 244984
rect 313332 244944 313338 244956
rect 352650 244944 352656 244956
rect 352708 244944 352714 244996
rect 158806 244876 158812 244928
rect 158864 244916 158870 244928
rect 171778 244916 171784 244928
rect 158864 244888 171784 244916
rect 158864 244876 158870 244888
rect 171778 244876 171784 244888
rect 171836 244876 171842 244928
rect 180150 244876 180156 244928
rect 180208 244916 180214 244928
rect 189074 244916 189080 244928
rect 180208 244888 189080 244916
rect 180208 244876 180214 244888
rect 189074 244876 189080 244888
rect 189132 244876 189138 244928
rect 190362 244876 190368 244928
rect 190420 244916 190426 244928
rect 197354 244916 197360 244928
rect 190420 244888 197360 244916
rect 190420 244876 190426 244888
rect 197354 244876 197360 244888
rect 197412 244876 197418 244928
rect 270402 244876 270408 244928
rect 270460 244916 270466 244928
rect 583018 244916 583024 244928
rect 270460 244888 583024 244916
rect 270460 244876 270466 244888
rect 583018 244876 583024 244888
rect 583076 244876 583082 244928
rect 67082 244400 67088 244452
rect 67140 244440 67146 244452
rect 67358 244440 67364 244452
rect 67140 244412 67364 244440
rect 67140 244400 67146 244412
rect 67358 244400 67364 244412
rect 67416 244400 67422 244452
rect 158806 244264 158812 244316
rect 158864 244304 158870 244316
rect 177298 244304 177304 244316
rect 158864 244276 177304 244304
rect 158864 244264 158870 244276
rect 177298 244264 177304 244276
rect 177356 244264 177362 244316
rect 269942 244264 269948 244316
rect 270000 244304 270006 244316
rect 270402 244304 270408 244316
rect 270000 244276 270408 244304
rect 270000 244264 270006 244276
rect 270402 244264 270408 244276
rect 270460 244264 270466 244316
rect 59262 244196 59268 244248
rect 59320 244236 59326 244248
rect 67450 244236 67456 244248
rect 59320 244208 67456 244236
rect 59320 244196 59326 244208
rect 67450 244196 67456 244208
rect 67508 244196 67514 244248
rect 246390 244196 246396 244248
rect 246448 244236 246454 244248
rect 249978 244236 249984 244248
rect 246448 244208 249984 244236
rect 246448 244196 246454 244208
rect 249978 244196 249984 244208
rect 250036 244196 250042 244248
rect 262122 243380 262128 243432
rect 262180 243420 262186 243432
rect 262398 243420 262404 243432
rect 262180 243392 262404 243420
rect 262180 243380 262186 243392
rect 262398 243380 262404 243392
rect 262456 243380 262462 243432
rect 158806 242972 158812 243024
rect 158864 243012 158870 243024
rect 181714 243012 181720 243024
rect 158864 242984 181720 243012
rect 158864 242972 158870 242984
rect 181714 242972 181720 242984
rect 181772 242972 181778 243024
rect 190178 242972 190184 243024
rect 190236 243012 190242 243024
rect 197354 243012 197360 243024
rect 190236 242984 197360 243012
rect 190236 242972 190242 242984
rect 197354 242972 197360 242984
rect 197412 242972 197418 243024
rect 245746 242972 245752 243024
rect 245804 243012 245810 243024
rect 262122 243012 262128 243024
rect 245804 242984 262128 243012
rect 245804 242972 245810 242984
rect 262122 242972 262128 242984
rect 262180 242972 262186 243024
rect 156966 242904 156972 242956
rect 157024 242944 157030 242956
rect 191190 242944 191196 242956
rect 157024 242916 191196 242944
rect 157024 242904 157030 242916
rect 191190 242904 191196 242916
rect 191248 242904 191254 242956
rect 262766 242904 262772 242956
rect 262824 242944 262830 242956
rect 409874 242944 409880 242956
rect 262824 242916 409880 242944
rect 262824 242904 262830 242916
rect 409874 242904 409880 242916
rect 409932 242904 409938 242956
rect 161014 242224 161020 242276
rect 161072 242264 161078 242276
rect 164142 242264 164148 242276
rect 161072 242236 164148 242264
rect 161072 242224 161078 242236
rect 164142 242224 164148 242236
rect 164200 242264 164206 242276
rect 177482 242264 177488 242276
rect 164200 242236 177488 242264
rect 164200 242224 164206 242236
rect 177482 242224 177488 242236
rect 177540 242224 177546 242276
rect 156874 242156 156880 242208
rect 156932 242196 156938 242208
rect 187510 242196 187516 242208
rect 156932 242168 187516 242196
rect 156932 242156 156938 242168
rect 187510 242156 187516 242168
rect 187568 242196 187574 242208
rect 199562 242196 199568 242208
rect 187568 242168 199568 242196
rect 187568 242156 187574 242168
rect 199562 242156 199568 242168
rect 199620 242156 199626 242208
rect 310606 242156 310612 242208
rect 310664 242196 310670 242208
rect 345750 242196 345756 242208
rect 310664 242168 345756 242196
rect 310664 242156 310670 242168
rect 345750 242156 345756 242168
rect 345808 242156 345814 242208
rect 153102 241476 153108 241528
rect 153160 241516 153166 241528
rect 156690 241516 156696 241528
rect 153160 241488 156696 241516
rect 153160 241476 153166 241488
rect 156690 241476 156696 241488
rect 156748 241476 156754 241528
rect 246114 241476 246120 241528
rect 246172 241516 246178 241528
rect 310606 241516 310612 241528
rect 246172 241488 310612 241516
rect 246172 241476 246178 241488
rect 310606 241476 310612 241488
rect 310664 241476 310670 241528
rect 57790 241408 57796 241460
rect 57848 241448 57854 241460
rect 83320 241448 83326 241460
rect 57848 241420 83326 241448
rect 57848 241408 57854 241420
rect 83320 241408 83326 241420
rect 83378 241408 83384 241460
rect 111104 241408 111110 241460
rect 111162 241448 111168 241460
rect 159634 241448 159640 241460
rect 111162 241420 159640 241448
rect 111162 241408 111168 241420
rect 159634 241408 159640 241420
rect 159692 241408 159698 241460
rect 67082 241340 67088 241392
rect 67140 241380 67146 241392
rect 73798 241380 73804 241392
rect 67140 241352 73804 241380
rect 67140 241340 67146 241352
rect 73798 241340 73804 241352
rect 73856 241340 73862 241392
rect 3326 241068 3332 241120
rect 3384 241108 3390 241120
rect 7558 241108 7564 241120
rect 3384 241080 7564 241108
rect 3384 241068 3390 241080
rect 7558 241068 7564 241080
rect 7616 241068 7622 241120
rect 159450 240796 159456 240848
rect 159508 240836 159514 240848
rect 170582 240836 170588 240848
rect 159508 240808 170588 240836
rect 159508 240796 159514 240808
rect 170582 240796 170588 240808
rect 170640 240796 170646 240848
rect 171870 240796 171876 240848
rect 171928 240836 171934 240848
rect 187050 240836 187056 240848
rect 171928 240808 187056 240836
rect 171928 240796 171934 240808
rect 187050 240796 187056 240808
rect 187108 240796 187114 240848
rect 195790 240796 195796 240848
rect 195848 240836 195854 240848
rect 197906 240836 197912 240848
rect 195848 240808 197912 240836
rect 195848 240796 195854 240808
rect 197906 240796 197912 240808
rect 197964 240796 197970 240848
rect 288342 240796 288348 240848
rect 288400 240836 288406 240848
rect 298738 240836 298744 240848
rect 288400 240808 298744 240836
rect 288400 240796 288406 240808
rect 298738 240796 298744 240808
rect 298796 240796 298802 240848
rect 98362 240728 98368 240780
rect 98420 240768 98426 240780
rect 160922 240768 160928 240780
rect 98420 240740 160928 240768
rect 98420 240728 98426 240740
rect 160922 240728 160928 240740
rect 160980 240728 160986 240780
rect 165154 240728 165160 240780
rect 165212 240768 165218 240780
rect 179414 240768 179420 240780
rect 165212 240740 179420 240768
rect 165212 240728 165218 240740
rect 179414 240728 179420 240740
rect 179472 240728 179478 240780
rect 245654 240728 245660 240780
rect 245712 240768 245718 240780
rect 452654 240768 452660 240780
rect 245712 240740 452660 240768
rect 245712 240728 245718 240740
rect 452654 240728 452660 240740
rect 452712 240728 452718 240780
rect 238726 240264 248414 240292
rect 200114 240184 200120 240236
rect 200172 240224 200178 240236
rect 200172 240196 209774 240224
rect 200172 240184 200178 240196
rect 77294 240116 77300 240168
rect 77352 240156 77358 240168
rect 77846 240156 77852 240168
rect 77352 240128 77852 240156
rect 77352 240116 77358 240128
rect 77846 240116 77852 240128
rect 77904 240116 77910 240168
rect 89714 240116 89720 240168
rect 89772 240156 89778 240168
rect 90358 240156 90364 240168
rect 89772 240128 90364 240156
rect 89772 240116 89778 240128
rect 90358 240116 90364 240128
rect 90416 240116 90422 240168
rect 91094 240116 91100 240168
rect 91152 240156 91158 240168
rect 91830 240156 91836 240168
rect 91152 240128 91836 240156
rect 91152 240116 91158 240128
rect 91830 240116 91836 240128
rect 91888 240116 91894 240168
rect 139394 240116 139400 240168
rect 139452 240156 139458 240168
rect 140038 240156 140044 240168
rect 139452 240128 140044 240156
rect 139452 240116 139458 240128
rect 140038 240116 140044 240128
rect 140096 240116 140102 240168
rect 186314 240116 186320 240168
rect 186372 240156 186378 240168
rect 202874 240156 202880 240168
rect 186372 240128 202880 240156
rect 186372 240116 186378 240128
rect 202874 240116 202880 240128
rect 202932 240156 202938 240168
rect 203426 240156 203432 240168
rect 202932 240128 203432 240156
rect 202932 240116 202938 240128
rect 203426 240116 203432 240128
rect 203484 240116 203490 240168
rect 209746 240156 209774 240196
rect 220722 240156 220728 240168
rect 209746 240128 220728 240156
rect 220722 240116 220728 240128
rect 220780 240116 220786 240168
rect 220906 240116 220912 240168
rect 220964 240156 220970 240168
rect 223298 240156 223304 240168
rect 220964 240128 223304 240156
rect 220964 240116 220970 240128
rect 223298 240116 223304 240128
rect 223356 240116 223362 240168
rect 232130 240116 232136 240168
rect 232188 240156 232194 240168
rect 238726 240156 238754 240264
rect 245654 240224 245660 240236
rect 232188 240128 238754 240156
rect 242636 240196 245660 240224
rect 232188 240116 232194 240128
rect 242636 240100 242664 240196
rect 245654 240184 245660 240196
rect 245712 240184 245718 240236
rect 248386 240156 248414 240264
rect 287238 240156 287244 240168
rect 248386 240128 287244 240156
rect 287238 240116 287244 240128
rect 287296 240156 287302 240168
rect 288342 240156 288348 240168
rect 287296 240128 288348 240156
rect 287296 240116 287302 240128
rect 288342 240116 288348 240128
rect 288400 240116 288406 240168
rect 69474 240048 69480 240100
rect 69532 240088 69538 240100
rect 72510 240088 72516 240100
rect 69532 240060 72516 240088
rect 69532 240048 69538 240060
rect 72510 240048 72516 240060
rect 72568 240048 72574 240100
rect 72602 240048 72608 240100
rect 72660 240088 72666 240100
rect 73062 240088 73068 240100
rect 72660 240060 73068 240088
rect 72660 240048 72666 240060
rect 73062 240048 73068 240060
rect 73120 240048 73126 240100
rect 81894 240048 81900 240100
rect 81952 240088 81958 240100
rect 82722 240088 82728 240100
rect 81952 240060 82728 240088
rect 81952 240048 81958 240060
rect 82722 240048 82728 240060
rect 82780 240048 82786 240100
rect 85574 240048 85580 240100
rect 85632 240088 85638 240100
rect 86862 240088 86868 240100
rect 85632 240060 86868 240088
rect 85632 240048 85638 240060
rect 86862 240048 86868 240060
rect 86920 240048 86926 240100
rect 93026 240048 93032 240100
rect 93084 240088 93090 240100
rect 93762 240088 93768 240100
rect 93084 240060 93768 240088
rect 93084 240048 93090 240060
rect 93762 240048 93768 240060
rect 93820 240048 93826 240100
rect 103790 240048 103796 240100
rect 103848 240088 103854 240100
rect 104802 240088 104808 240100
rect 103848 240060 104808 240088
rect 103848 240048 103854 240060
rect 104802 240048 104808 240060
rect 104860 240048 104866 240100
rect 114646 240048 114652 240100
rect 114704 240088 114710 240100
rect 115198 240088 115204 240100
rect 114704 240060 115204 240088
rect 114704 240048 114710 240060
rect 115198 240048 115204 240060
rect 115256 240048 115262 240100
rect 119338 240048 119344 240100
rect 119396 240088 119402 240100
rect 119982 240088 119988 240100
rect 119396 240060 119988 240088
rect 119396 240048 119402 240060
rect 119982 240048 119988 240060
rect 120040 240048 120046 240100
rect 127158 240048 127164 240100
rect 127216 240088 127222 240100
rect 128262 240088 128268 240100
rect 127216 240060 128268 240088
rect 127216 240048 127222 240060
rect 128262 240048 128268 240060
rect 128320 240048 128326 240100
rect 131850 240048 131856 240100
rect 131908 240088 131914 240100
rect 132310 240088 132316 240100
rect 131908 240060 132316 240088
rect 131908 240048 131914 240060
rect 132310 240048 132316 240060
rect 132368 240048 132374 240100
rect 142890 240048 142896 240100
rect 142948 240088 142954 240100
rect 143442 240088 143448 240100
rect 142948 240060 143448 240088
rect 142948 240048 142954 240060
rect 143442 240048 143448 240060
rect 143500 240048 143506 240100
rect 143626 240048 143632 240100
rect 143684 240088 143690 240100
rect 144270 240088 144276 240100
rect 143684 240060 144276 240088
rect 143684 240048 143690 240060
rect 144270 240048 144276 240060
rect 144328 240048 144334 240100
rect 153286 240048 153292 240100
rect 153344 240088 153350 240100
rect 153838 240088 153844 240100
rect 153344 240060 153844 240088
rect 153344 240048 153350 240060
rect 153838 240048 153844 240060
rect 153896 240048 153902 240100
rect 195238 240048 195244 240100
rect 195296 240088 195302 240100
rect 201126 240088 201132 240100
rect 195296 240060 201132 240088
rect 195296 240048 195302 240060
rect 201126 240048 201132 240060
rect 201184 240048 201190 240100
rect 228726 240048 228732 240100
rect 228784 240088 228790 240100
rect 228784 240060 238754 240088
rect 228784 240048 228790 240060
rect 67358 239980 67364 240032
rect 67416 240020 67422 240032
rect 69658 240020 69664 240032
rect 67416 239992 69664 240020
rect 67416 239980 67422 239992
rect 69658 239980 69664 239992
rect 69716 239980 69722 240032
rect 199838 239980 199844 240032
rect 199896 240020 199902 240032
rect 201034 240020 201040 240032
rect 199896 239992 201040 240020
rect 199896 239980 199902 239992
rect 201034 239980 201040 239992
rect 201092 239980 201098 240032
rect 232590 239980 232596 240032
rect 232648 240020 232654 240032
rect 237466 240020 237472 240032
rect 232648 239992 237472 240020
rect 232648 239980 232654 239992
rect 237466 239980 237472 239992
rect 237524 239980 237530 240032
rect 80698 239912 80704 239964
rect 80756 239952 80762 239964
rect 81250 239952 81256 239964
rect 80756 239924 81256 239952
rect 80756 239912 80762 239924
rect 81250 239912 81256 239924
rect 81308 239912 81314 239964
rect 88794 239912 88800 239964
rect 88852 239952 88858 239964
rect 89530 239952 89536 239964
rect 88852 239924 89536 239952
rect 88852 239912 88858 239924
rect 89530 239912 89536 239924
rect 89588 239912 89594 239964
rect 110690 239912 110696 239964
rect 110748 239952 110754 239964
rect 111702 239952 111708 239964
rect 110748 239924 111708 239952
rect 110748 239912 110754 239924
rect 111702 239912 111708 239924
rect 111760 239912 111766 239964
rect 153746 239912 153752 239964
rect 153804 239952 153810 239964
rect 154482 239952 154488 239964
rect 153804 239924 154488 239952
rect 153804 239912 153810 239924
rect 154482 239912 154488 239924
rect 154540 239912 154546 239964
rect 238726 239952 238754 240060
rect 242618 240048 242624 240100
rect 242676 240048 242682 240100
rect 257522 239952 257528 239964
rect 238726 239924 257528 239952
rect 257522 239912 257528 239924
rect 257580 239912 257586 239964
rect 99650 239776 99656 239828
rect 99708 239816 99714 239828
rect 100570 239816 100576 239828
rect 99708 239788 100576 239816
rect 99708 239776 99714 239788
rect 100570 239776 100576 239788
rect 100628 239776 100634 239828
rect 133322 239708 133328 239760
rect 133380 239748 133386 239760
rect 133782 239748 133788 239760
rect 133380 239720 133788 239748
rect 133380 239708 133386 239720
rect 133782 239708 133788 239720
rect 133840 239708 133846 239760
rect 84102 239436 84108 239488
rect 84160 239476 84166 239488
rect 97350 239476 97356 239488
rect 84160 239448 97356 239476
rect 84160 239436 84166 239448
rect 97350 239436 97356 239448
rect 97408 239436 97414 239488
rect 108942 239436 108948 239488
rect 109000 239476 109006 239488
rect 206002 239476 206008 239488
rect 109000 239448 206008 239476
rect 109000 239436 109006 239448
rect 206002 239436 206008 239448
rect 206060 239436 206066 239488
rect 305086 239436 305092 239488
rect 305144 239476 305150 239488
rect 322934 239476 322940 239488
rect 305144 239448 322940 239476
rect 305144 239436 305150 239448
rect 322934 239436 322940 239448
rect 322992 239436 322998 239488
rect 68922 239368 68928 239420
rect 68980 239408 68986 239420
rect 191834 239408 191840 239420
rect 68980 239380 191840 239408
rect 68980 239368 68986 239380
rect 191834 239368 191840 239380
rect 191892 239368 191898 239420
rect 224402 239368 224408 239420
rect 224460 239408 224466 239420
rect 232038 239408 232044 239420
rect 224460 239380 232044 239408
rect 224460 239368 224466 239380
rect 232038 239368 232044 239380
rect 232096 239368 232102 239420
rect 317506 239368 317512 239420
rect 317564 239408 317570 239420
rect 342254 239408 342260 239420
rect 317564 239380 342260 239408
rect 317564 239368 317570 239380
rect 342254 239368 342260 239380
rect 342312 239368 342318 239420
rect 92566 239232 92572 239284
rect 92624 239272 92630 239284
rect 93118 239272 93124 239284
rect 92624 239244 93124 239272
rect 92624 239232 92630 239244
rect 93118 239232 93124 239244
rect 93176 239232 93182 239284
rect 105538 239232 105544 239284
rect 105596 239272 105602 239284
rect 106182 239272 106188 239284
rect 105596 239244 106188 239272
rect 105596 239232 105602 239244
rect 106182 239232 106188 239244
rect 106240 239232 106246 239284
rect 120810 239232 120816 239284
rect 120868 239272 120874 239284
rect 121362 239272 121368 239284
rect 120868 239244 121368 239272
rect 120868 239232 120874 239244
rect 121362 239232 121368 239244
rect 121420 239232 121426 239284
rect 128906 239232 128912 239284
rect 128964 239272 128970 239284
rect 129550 239272 129556 239284
rect 128964 239244 129556 239272
rect 128964 239232 128970 239244
rect 129550 239232 129556 239244
rect 129608 239232 129614 239284
rect 141418 239232 141424 239284
rect 141476 239272 141482 239284
rect 141970 239272 141976 239284
rect 141476 239244 141976 239272
rect 141476 239232 141482 239244
rect 141970 239232 141976 239244
rect 142028 239232 142034 239284
rect 144178 239232 144184 239284
rect 144236 239272 144242 239284
rect 144822 239272 144828 239284
rect 144236 239244 144828 239272
rect 144236 239232 144242 239244
rect 144822 239232 144828 239244
rect 144880 239232 144886 239284
rect 147122 239232 147128 239284
rect 147180 239272 147186 239284
rect 147582 239272 147588 239284
rect 147180 239244 147588 239272
rect 147180 239232 147186 239244
rect 147582 239232 147588 239244
rect 147640 239232 147646 239284
rect 117314 239164 117320 239216
rect 117372 239204 117378 239216
rect 117958 239204 117964 239216
rect 117372 239176 117964 239204
rect 117372 239164 117378 239176
rect 117958 239164 117964 239176
rect 118016 239164 118022 239216
rect 115106 239096 115112 239148
rect 115164 239136 115170 239148
rect 115842 239136 115848 239148
rect 115164 239108 115848 239136
rect 115164 239096 115170 239108
rect 115842 239096 115848 239108
rect 115900 239096 115906 239148
rect 273162 238824 273168 238876
rect 273220 238864 273226 238876
rect 283190 238864 283196 238876
rect 273220 238836 283196 238864
rect 273220 238824 273226 238836
rect 283190 238824 283196 238836
rect 283248 238824 283254 238876
rect 240318 238756 240324 238808
rect 240376 238796 240382 238808
rect 240870 238796 240876 238808
rect 240376 238768 240876 238796
rect 240376 238756 240382 238768
rect 240870 238756 240876 238768
rect 240928 238796 240934 238808
rect 317506 238796 317512 238808
rect 240928 238768 317512 238796
rect 240928 238756 240934 238768
rect 317506 238756 317512 238768
rect 317564 238756 317570 238808
rect 13078 238688 13084 238740
rect 13136 238728 13142 238740
rect 92566 238728 92572 238740
rect 13136 238700 92572 238728
rect 13136 238688 13142 238700
rect 92566 238688 92572 238700
rect 92624 238688 92630 238740
rect 222286 238688 222292 238740
rect 222344 238728 222350 238740
rect 273162 238728 273168 238740
rect 222344 238700 273168 238728
rect 222344 238688 222350 238700
rect 273162 238688 273168 238700
rect 273220 238688 273226 238740
rect 50890 238620 50896 238672
rect 50948 238660 50954 238672
rect 75914 238660 75920 238672
rect 50948 238632 75920 238660
rect 50948 238620 50954 238632
rect 75914 238620 75920 238632
rect 75972 238620 75978 238672
rect 121638 238620 121644 238672
rect 121696 238660 121702 238672
rect 183370 238660 183376 238672
rect 121696 238632 183376 238660
rect 121696 238620 121702 238632
rect 183370 238620 183376 238632
rect 183428 238620 183434 238672
rect 206002 238620 206008 238672
rect 206060 238660 206066 238672
rect 219894 238660 219900 238672
rect 206060 238632 219900 238660
rect 206060 238620 206066 238632
rect 219894 238620 219900 238632
rect 219952 238620 219958 238672
rect 113174 238552 113180 238604
rect 113232 238592 113238 238604
rect 222304 238592 222332 238688
rect 241790 238620 241796 238672
rect 241848 238660 241854 238672
rect 252646 238660 252652 238672
rect 241848 238632 252652 238660
rect 241848 238620 241854 238632
rect 252646 238620 252652 238632
rect 252704 238620 252710 238672
rect 113232 238564 222332 238592
rect 113232 238552 113238 238564
rect 239214 238144 239220 238196
rect 239272 238184 239278 238196
rect 242710 238184 242716 238196
rect 239272 238156 242716 238184
rect 239272 238144 239278 238156
rect 242710 238144 242716 238156
rect 242768 238144 242774 238196
rect 259362 238076 259368 238128
rect 259420 238116 259426 238128
rect 262950 238116 262956 238128
rect 259420 238088 262956 238116
rect 259420 238076 259426 238088
rect 262950 238076 262956 238088
rect 263008 238076 263014 238128
rect 199378 238008 199384 238060
rect 199436 238048 199442 238060
rect 200206 238048 200212 238060
rect 199436 238020 200212 238048
rect 199436 238008 199442 238020
rect 200206 238008 200212 238020
rect 200264 238008 200270 238060
rect 224770 238008 224776 238060
rect 224828 238048 224834 238060
rect 232958 238048 232964 238060
rect 224828 238020 232964 238048
rect 224828 238008 224834 238020
rect 232958 238008 232964 238020
rect 233016 238008 233022 238060
rect 285122 238008 285128 238060
rect 285180 238048 285186 238060
rect 385678 238048 385684 238060
rect 285180 238020 385684 238048
rect 285180 238008 285186 238020
rect 385678 238008 385684 238020
rect 385736 238008 385742 238060
rect 191834 237668 191840 237720
rect 191892 237708 191898 237720
rect 194410 237708 194416 237720
rect 191892 237680 194416 237708
rect 191892 237668 191898 237680
rect 194410 237668 194416 237680
rect 194468 237708 194474 237720
rect 199378 237708 199384 237720
rect 194468 237680 199384 237708
rect 194468 237668 194474 237680
rect 199378 237668 199384 237680
rect 199436 237668 199442 237720
rect 237466 237532 237472 237584
rect 237524 237572 237530 237584
rect 239398 237572 239404 237584
rect 237524 237544 239404 237572
rect 237524 237532 237530 237544
rect 239398 237532 239404 237544
rect 239456 237532 239462 237584
rect 236822 237464 236828 237516
rect 236880 237504 236886 237516
rect 238018 237504 238024 237516
rect 236880 237476 238024 237504
rect 236880 237464 236886 237476
rect 238018 237464 238024 237476
rect 238076 237464 238082 237516
rect 75914 237396 75920 237448
rect 75972 237436 75978 237448
rect 76558 237436 76564 237448
rect 75972 237408 76564 237436
rect 75972 237396 75978 237408
rect 76558 237396 76564 237408
rect 76616 237396 76622 237448
rect 92566 237396 92572 237448
rect 92624 237436 92630 237448
rect 93118 237436 93124 237448
rect 92624 237408 93124 237436
rect 92624 237396 92630 237408
rect 93118 237396 93124 237408
rect 93176 237396 93182 237448
rect 207106 237396 207112 237448
rect 207164 237436 207170 237448
rect 207934 237436 207940 237448
rect 207164 237408 207940 237436
rect 207164 237396 207170 237408
rect 207934 237396 207940 237408
rect 207992 237396 207998 237448
rect 214190 237396 214196 237448
rect 214248 237436 214254 237448
rect 214650 237436 214656 237448
rect 214248 237408 214656 237436
rect 214248 237396 214254 237408
rect 214650 237396 214656 237408
rect 214708 237396 214714 237448
rect 215662 237396 215668 237448
rect 215720 237436 215726 237448
rect 216490 237436 216496 237448
rect 215720 237408 216496 237436
rect 215720 237396 215726 237408
rect 216490 237396 216496 237408
rect 216548 237396 216554 237448
rect 55030 237328 55036 237380
rect 55088 237368 55094 237380
rect 77386 237368 77392 237380
rect 55088 237340 77392 237368
rect 55088 237328 55094 237340
rect 77386 237328 77392 237340
rect 77444 237328 77450 237380
rect 199562 237328 199568 237380
rect 199620 237368 199626 237380
rect 202966 237368 202972 237380
rect 199620 237340 202972 237368
rect 199620 237328 199626 237340
rect 202966 237328 202972 237340
rect 203024 237328 203030 237380
rect 155954 237260 155960 237312
rect 156012 237300 156018 237312
rect 160738 237300 160744 237312
rect 156012 237272 160744 237300
rect 156012 237260 156018 237272
rect 160738 237260 160744 237272
rect 160796 237260 160802 237312
rect 149054 236784 149060 236836
rect 149112 236824 149118 236836
rect 149238 236824 149244 236836
rect 149112 236796 149244 236824
rect 149112 236784 149118 236796
rect 149238 236784 149244 236796
rect 149296 236784 149302 236836
rect 128998 236716 129004 236768
rect 129056 236756 129062 236768
rect 136818 236756 136824 236768
rect 129056 236728 136824 236756
rect 129056 236716 129062 236728
rect 136818 236716 136824 236728
rect 136876 236716 136882 236768
rect 139486 236716 139492 236768
rect 139544 236756 139550 236768
rect 156966 236756 156972 236768
rect 139544 236728 156972 236756
rect 139544 236716 139550 236728
rect 156966 236716 156972 236728
rect 157024 236716 157030 236768
rect 177298 236716 177304 236768
rect 177356 236756 177362 236768
rect 192938 236756 192944 236768
rect 177356 236728 192944 236756
rect 177356 236716 177362 236728
rect 192938 236716 192944 236728
rect 192996 236716 193002 236768
rect 67726 236648 67732 236700
rect 67784 236688 67790 236700
rect 236638 236688 236644 236700
rect 67784 236660 236644 236688
rect 67784 236648 67790 236660
rect 236638 236648 236644 236660
rect 236696 236688 236702 236700
rect 248598 236688 248604 236700
rect 236696 236660 248604 236688
rect 236696 236648 236702 236660
rect 248598 236648 248604 236660
rect 248656 236648 248662 236700
rect 313366 236648 313372 236700
rect 313424 236688 313430 236700
rect 333974 236688 333980 236700
rect 313424 236660 333980 236688
rect 313424 236648 313430 236660
rect 333974 236648 333980 236660
rect 334032 236648 334038 236700
rect 342898 236648 342904 236700
rect 342956 236688 342962 236700
rect 363690 236688 363696 236700
rect 342956 236660 363696 236688
rect 342956 236648 342962 236660
rect 363690 236648 363696 236660
rect 363748 236648 363754 236700
rect 284938 236036 284944 236088
rect 284996 236076 285002 236088
rect 286410 236076 286416 236088
rect 284996 236048 286416 236076
rect 284996 236036 285002 236048
rect 286410 236036 286416 236048
rect 286468 236036 286474 236088
rect 202966 235968 202972 236020
rect 203024 236008 203030 236020
rect 203518 236008 203524 236020
rect 203024 235980 203524 236008
rect 203024 235968 203030 235980
rect 203518 235968 203524 235980
rect 203576 235968 203582 236020
rect 204070 235968 204076 236020
rect 204128 236008 204134 236020
rect 226978 236008 226984 236020
rect 204128 235980 226984 236008
rect 204128 235968 204134 235980
rect 226978 235968 226984 235980
rect 227036 235968 227042 236020
rect 239398 235968 239404 236020
rect 239456 236008 239462 236020
rect 313366 236008 313372 236020
rect 239456 235980 313372 236008
rect 239456 235968 239462 235980
rect 313366 235968 313372 235980
rect 313424 235968 313430 236020
rect 46842 235900 46848 235952
rect 46900 235940 46906 235952
rect 143626 235940 143632 235952
rect 46900 235912 143632 235940
rect 46900 235900 46906 235912
rect 143626 235900 143632 235912
rect 143684 235940 143690 235952
rect 144178 235940 144184 235952
rect 143684 235912 144184 235940
rect 143684 235900 143690 235912
rect 144178 235900 144184 235912
rect 144236 235900 144242 235952
rect 149054 235900 149060 235952
rect 149112 235940 149118 235952
rect 167638 235940 167644 235952
rect 149112 235912 167644 235940
rect 149112 235900 149118 235912
rect 167638 235900 167644 235912
rect 167696 235900 167702 235952
rect 57698 235832 57704 235884
rect 57756 235872 57762 235884
rect 103514 235872 103520 235884
rect 57756 235844 103520 235872
rect 57756 235832 57762 235844
rect 103514 235832 103520 235844
rect 103572 235872 103578 235884
rect 104710 235872 104716 235884
rect 103572 235844 104716 235872
rect 103572 235832 103578 235844
rect 104710 235832 104716 235844
rect 104768 235832 104774 235884
rect 125594 235832 125600 235884
rect 125652 235872 125658 235884
rect 139486 235872 139492 235884
rect 125652 235844 139492 235872
rect 125652 235832 125658 235844
rect 139486 235832 139492 235844
rect 139544 235832 139550 235884
rect 199470 235832 199476 235884
rect 199528 235872 199534 235884
rect 223758 235872 223764 235884
rect 199528 235844 223764 235872
rect 199528 235832 199534 235844
rect 223758 235832 223764 235844
rect 223816 235832 223822 235884
rect 201126 235560 201132 235612
rect 201184 235600 201190 235612
rect 206370 235600 206376 235612
rect 201184 235572 206376 235600
rect 201184 235560 201190 235572
rect 206370 235560 206376 235572
rect 206428 235560 206434 235612
rect 139578 235220 139584 235272
rect 139636 235260 139642 235272
rect 150434 235260 150440 235272
rect 139636 235232 150440 235260
rect 139636 235220 139642 235232
rect 150434 235220 150440 235232
rect 150492 235220 150498 235272
rect 182082 235220 182088 235272
rect 182140 235260 182146 235272
rect 196618 235260 196624 235272
rect 182140 235232 196624 235260
rect 182140 235220 182146 235232
rect 196618 235220 196624 235232
rect 196676 235220 196682 235272
rect 270402 235220 270408 235272
rect 270460 235260 270466 235272
rect 294690 235260 294696 235272
rect 270460 235232 294696 235260
rect 270460 235220 270466 235232
rect 294690 235220 294696 235232
rect 294748 235220 294754 235272
rect 174630 235084 174636 235136
rect 174688 235124 174694 235136
rect 177298 235124 177304 235136
rect 174688 235096 177304 235124
rect 174688 235084 174694 235096
rect 177298 235084 177304 235096
rect 177356 235084 177362 235136
rect 195974 234880 195980 234932
rect 196032 234920 196038 234932
rect 199378 234920 199384 234932
rect 196032 234892 199384 234920
rect 196032 234880 196038 234892
rect 199378 234880 199384 234892
rect 199436 234880 199442 234932
rect 214742 234676 214748 234728
rect 214800 234716 214806 234728
rect 215110 234716 215116 234728
rect 214800 234688 215116 234716
rect 214800 234676 214806 234688
rect 215110 234676 215116 234688
rect 215168 234716 215174 234728
rect 233326 234716 233332 234728
rect 215168 234688 233332 234716
rect 215168 234676 215174 234688
rect 233326 234676 233332 234688
rect 233384 234676 233390 234728
rect 240778 234676 240784 234728
rect 240836 234716 240842 234728
rect 246022 234716 246028 234728
rect 240836 234688 246028 234716
rect 240836 234676 240842 234688
rect 246022 234676 246028 234688
rect 246080 234676 246086 234728
rect 155218 234608 155224 234660
rect 155276 234648 155282 234660
rect 184750 234648 184756 234660
rect 155276 234620 184756 234648
rect 155276 234608 155282 234620
rect 184750 234608 184756 234620
rect 184808 234648 184814 234660
rect 185026 234648 185032 234660
rect 184808 234620 185032 234648
rect 184808 234608 184814 234620
rect 185026 234608 185032 234620
rect 185084 234608 185090 234660
rect 223758 234608 223764 234660
rect 223816 234648 223822 234660
rect 224218 234648 224224 234660
rect 223816 234620 224224 234648
rect 223816 234608 223822 234620
rect 224218 234608 224224 234620
rect 224276 234608 224282 234660
rect 230198 234608 230204 234660
rect 230256 234648 230262 234660
rect 231946 234648 231952 234660
rect 230256 234620 231952 234648
rect 230256 234608 230262 234620
rect 231946 234608 231952 234620
rect 232004 234648 232010 234660
rect 434806 234648 434812 234660
rect 232004 234620 434812 234648
rect 232004 234608 232010 234620
rect 434806 234608 434812 234620
rect 434864 234608 434870 234660
rect 149238 234540 149244 234592
rect 149296 234580 149302 234592
rect 231854 234580 231860 234592
rect 149296 234552 231860 234580
rect 149296 234540 149302 234552
rect 231854 234540 231860 234552
rect 231912 234540 231918 234592
rect 267642 234540 267648 234592
rect 267700 234580 267706 234592
rect 269758 234580 269764 234592
rect 267700 234552 269764 234580
rect 267700 234540 267734 234552
rect 269758 234540 269764 234552
rect 269816 234540 269822 234592
rect 324314 234540 324320 234592
rect 324372 234580 324378 234592
rect 325602 234580 325608 234592
rect 324372 234552 325608 234580
rect 324372 234540 324378 234552
rect 325602 234540 325608 234552
rect 325660 234580 325666 234592
rect 327718 234580 327724 234592
rect 325660 234552 327724 234580
rect 325660 234540 325666 234552
rect 327718 234540 327724 234552
rect 327776 234540 327782 234592
rect 158070 234472 158076 234524
rect 158128 234512 158134 234524
rect 162302 234512 162308 234524
rect 158128 234484 162308 234512
rect 158128 234472 158134 234484
rect 162302 234472 162308 234484
rect 162360 234472 162366 234524
rect 201310 234472 201316 234524
rect 201368 234512 201374 234524
rect 218146 234512 218152 234524
rect 201368 234484 218152 234512
rect 201368 234472 201374 234484
rect 218146 234472 218152 234484
rect 218204 234472 218210 234524
rect 219894 234472 219900 234524
rect 219952 234512 219958 234524
rect 267706 234512 267734 234540
rect 219952 234484 267734 234512
rect 219952 234472 219958 234484
rect 138014 233928 138020 233980
rect 138072 233968 138078 233980
rect 148318 233968 148324 233980
rect 138072 233940 148324 233968
rect 138072 233928 138078 233940
rect 148318 233928 148324 233940
rect 148376 233928 148382 233980
rect 60274 233860 60280 233912
rect 60332 233900 60338 233912
rect 147674 233900 147680 233912
rect 60332 233872 147680 233900
rect 60332 233860 60338 233872
rect 147674 233860 147680 233872
rect 147732 233860 147738 233912
rect 176102 233860 176108 233912
rect 176160 233900 176166 233912
rect 191190 233900 191196 233912
rect 176160 233872 191196 233900
rect 176160 233860 176166 233872
rect 191190 233860 191196 233872
rect 191248 233860 191254 233912
rect 104894 233180 104900 233232
rect 104952 233220 104958 233232
rect 188430 233220 188436 233232
rect 104952 233192 188436 233220
rect 104952 233180 104958 233192
rect 188430 233180 188436 233192
rect 188488 233180 188494 233232
rect 191282 233180 191288 233232
rect 191340 233220 191346 233232
rect 222838 233220 222844 233232
rect 191340 233192 222844 233220
rect 191340 233180 191346 233192
rect 222838 233180 222844 233192
rect 222896 233220 222902 233232
rect 223390 233220 223396 233232
rect 222896 233192 223396 233220
rect 222896 233180 222902 233192
rect 223390 233180 223396 233192
rect 223448 233180 223454 233232
rect 192478 233112 192484 233164
rect 192536 233152 192542 233164
rect 206830 233152 206836 233164
rect 192536 233124 206836 233152
rect 192536 233112 192542 233124
rect 206830 233112 206836 233124
rect 206888 233112 206894 233164
rect 232958 232568 232964 232620
rect 233016 232608 233022 232620
rect 242158 232608 242164 232620
rect 233016 232580 242164 232608
rect 233016 232568 233022 232580
rect 242158 232568 242164 232580
rect 242216 232568 242222 232620
rect 61930 232500 61936 232552
rect 61988 232540 61994 232552
rect 123478 232540 123484 232552
rect 61988 232512 123484 232540
rect 61988 232500 61994 232512
rect 123478 232500 123484 232512
rect 123536 232500 123542 232552
rect 150434 232500 150440 232552
rect 150492 232540 150498 232552
rect 191650 232540 191656 232552
rect 150492 232512 191656 232540
rect 150492 232500 150498 232512
rect 191650 232500 191656 232512
rect 191708 232500 191714 232552
rect 226150 232500 226156 232552
rect 226208 232540 226214 232552
rect 284386 232540 284392 232552
rect 226208 232512 284392 232540
rect 226208 232500 226214 232512
rect 284386 232500 284392 232512
rect 284444 232500 284450 232552
rect 285030 232500 285036 232552
rect 285088 232540 285094 232552
rect 378778 232540 378784 232552
rect 285088 232512 378784 232540
rect 285088 232500 285094 232512
rect 378778 232500 378784 232512
rect 378836 232500 378842 232552
rect 139486 231860 139492 231872
rect 128372 231832 139492 231860
rect 114278 231752 114284 231804
rect 114336 231792 114342 231804
rect 128372 231792 128400 231832
rect 139486 231820 139492 231832
rect 139544 231820 139550 231872
rect 114336 231764 128400 231792
rect 114336 231752 114342 231764
rect 147674 231752 147680 231804
rect 147732 231792 147738 231804
rect 173250 231792 173256 231804
rect 147732 231764 173256 231792
rect 147732 231752 147738 231764
rect 173250 231752 173256 231764
rect 173308 231752 173314 231804
rect 191650 231752 191656 231804
rect 191708 231792 191714 231804
rect 224402 231792 224408 231804
rect 191708 231764 224408 231792
rect 191708 231752 191714 231764
rect 224402 231752 224408 231764
rect 224460 231752 224466 231804
rect 240042 231752 240048 231804
rect 240100 231792 240106 231804
rect 291286 231792 291292 231804
rect 240100 231764 291292 231792
rect 240100 231752 240106 231764
rect 291286 231752 291292 231764
rect 291344 231792 291350 231804
rect 291838 231792 291844 231804
rect 291344 231764 291844 231792
rect 291344 231752 291350 231764
rect 291838 231752 291844 231764
rect 291896 231752 291902 231804
rect 156598 231684 156604 231736
rect 156656 231724 156662 231736
rect 157978 231724 157984 231736
rect 156656 231696 157984 231724
rect 156656 231684 156662 231696
rect 157978 231684 157984 231696
rect 158036 231684 158042 231736
rect 129550 231208 129556 231260
rect 129608 231248 129614 231260
rect 143350 231248 143356 231260
rect 129608 231220 143356 231248
rect 129608 231208 129614 231220
rect 143350 231208 143356 231220
rect 143408 231208 143414 231260
rect 100570 231140 100576 231192
rect 100628 231180 100634 231192
rect 108298 231180 108304 231192
rect 100628 231152 108304 231180
rect 100628 231140 100634 231152
rect 108298 231140 108304 231152
rect 108356 231140 108362 231192
rect 139118 231140 139124 231192
rect 139176 231180 139182 231192
rect 156874 231180 156880 231192
rect 139176 231152 156880 231180
rect 139176 231140 139182 231152
rect 156874 231140 156880 231152
rect 156932 231140 156938 231192
rect 65886 231072 65892 231124
rect 65944 231112 65950 231124
rect 139210 231112 139216 231124
rect 65944 231084 139216 231112
rect 65944 231072 65950 231084
rect 139210 231072 139216 231084
rect 139268 231072 139274 231124
rect 164142 231072 164148 231124
rect 164200 231112 164206 231124
rect 197262 231112 197268 231124
rect 164200 231084 197268 231112
rect 164200 231072 164206 231084
rect 197262 231072 197268 231084
rect 197320 231072 197326 231124
rect 198550 231072 198556 231124
rect 198608 231112 198614 231124
rect 266354 231112 266360 231124
rect 198608 231084 266360 231112
rect 198608 231072 198614 231084
rect 266354 231072 266360 231084
rect 266412 231072 266418 231124
rect 180058 230460 180064 230512
rect 180116 230500 180122 230512
rect 181622 230500 181628 230512
rect 180116 230472 181628 230500
rect 180116 230460 180122 230472
rect 181622 230460 181628 230472
rect 181680 230460 181686 230512
rect 143350 230392 143356 230444
rect 143408 230432 143414 230444
rect 160094 230432 160100 230444
rect 143408 230404 160100 230432
rect 143408 230392 143414 230404
rect 160094 230392 160100 230404
rect 160152 230392 160158 230444
rect 184658 230392 184664 230444
rect 184716 230432 184722 230444
rect 185670 230432 185676 230444
rect 184716 230404 185676 230432
rect 184716 230392 184722 230404
rect 185670 230392 185676 230404
rect 185728 230392 185734 230444
rect 194226 230392 194232 230444
rect 194284 230432 194290 230444
rect 214742 230432 214748 230444
rect 194284 230404 214748 230432
rect 194284 230392 194290 230404
rect 214742 230392 214748 230404
rect 214800 230392 214806 230444
rect 233050 230392 233056 230444
rect 233108 230432 233114 230444
rect 233418 230432 233424 230444
rect 233108 230404 233424 230432
rect 233108 230392 233114 230404
rect 233418 230392 233424 230404
rect 233476 230392 233482 230444
rect 270402 230392 270408 230444
rect 270460 230432 270466 230444
rect 271138 230432 271144 230444
rect 270460 230404 271144 230432
rect 270460 230392 270466 230404
rect 271138 230392 271144 230404
rect 271196 230392 271202 230444
rect 139486 230324 139492 230376
rect 139544 230364 139550 230376
rect 152734 230364 152740 230376
rect 139544 230336 152740 230364
rect 139544 230324 139550 230336
rect 152734 230324 152740 230336
rect 152792 230324 152798 230376
rect 197262 230324 197268 230376
rect 197320 230364 197326 230376
rect 204990 230364 204996 230376
rect 197320 230336 204996 230364
rect 197320 230324 197326 230336
rect 204990 230324 204996 230336
rect 205048 230324 205054 230376
rect 86954 229780 86960 229832
rect 87012 229820 87018 229832
rect 105538 229820 105544 229832
rect 87012 229792 105544 229820
rect 87012 229780 87018 229792
rect 105538 229780 105544 229792
rect 105596 229780 105602 229832
rect 249794 229820 249800 229832
rect 229066 229792 249800 229820
rect 81250 229712 81256 229764
rect 81308 229752 81314 229764
rect 97258 229752 97264 229764
rect 81308 229724 97264 229752
rect 81308 229712 81314 229724
rect 97258 229712 97264 229724
rect 97316 229712 97322 229764
rect 100754 229712 100760 229764
rect 100812 229752 100818 229764
rect 140774 229752 140780 229764
rect 100812 229724 140780 229752
rect 100812 229712 100818 229724
rect 140774 229712 140780 229724
rect 140832 229712 140838 229764
rect 177390 229712 177396 229764
rect 177448 229752 177454 229764
rect 194226 229752 194232 229764
rect 177448 229724 194232 229752
rect 177448 229712 177454 229724
rect 194226 229712 194232 229724
rect 194284 229712 194290 229764
rect 217318 229712 217324 229764
rect 217376 229752 217382 229764
rect 227254 229752 227260 229764
rect 217376 229724 227260 229752
rect 217376 229712 217382 229724
rect 227254 229712 227260 229724
rect 227312 229752 227318 229764
rect 229066 229752 229094 229792
rect 249794 229780 249800 229792
rect 249852 229780 249858 229832
rect 266354 229780 266360 229832
rect 266412 229820 266418 229832
rect 270402 229820 270408 229832
rect 266412 229792 270408 229820
rect 266412 229780 266418 229792
rect 270402 229780 270408 229792
rect 270460 229780 270466 229832
rect 227312 229724 229094 229752
rect 227312 229712 227318 229724
rect 230382 229712 230388 229764
rect 230440 229752 230446 229764
rect 231118 229752 231124 229764
rect 230440 229724 231124 229752
rect 230440 229712 230446 229724
rect 231118 229712 231124 229724
rect 231176 229712 231182 229764
rect 233418 229712 233424 229764
rect 233476 229752 233482 229764
rect 295334 229752 295340 229764
rect 233476 229724 295340 229752
rect 233476 229712 233482 229724
rect 295334 229712 295340 229724
rect 295392 229712 295398 229764
rect 206830 229100 206836 229152
rect 206888 229140 206894 229152
rect 211798 229140 211804 229152
rect 206888 229112 211804 229140
rect 206888 229100 206894 229112
rect 211798 229100 211804 229112
rect 211856 229100 211862 229152
rect 95326 229032 95332 229084
rect 95384 229072 95390 229084
rect 244274 229072 244280 229084
rect 95384 229044 244280 229072
rect 95384 229032 95390 229044
rect 244274 229032 244280 229044
rect 244332 229032 244338 229084
rect 194226 228964 194232 229016
rect 194284 229004 194290 229016
rect 220078 229004 220084 229016
rect 194284 228976 220084 229004
rect 194284 228964 194290 228976
rect 220078 228964 220084 228976
rect 220136 228964 220142 229016
rect 244274 228760 244280 228812
rect 244332 228800 244338 228812
rect 245010 228800 245016 228812
rect 244332 228772 245016 228800
rect 244332 228760 244338 228772
rect 245010 228760 245016 228772
rect 245068 228760 245074 228812
rect 64506 228352 64512 228404
rect 64564 228392 64570 228404
rect 115014 228392 115020 228404
rect 64564 228364 115020 228392
rect 64564 228352 64570 228364
rect 115014 228352 115020 228364
rect 115072 228352 115078 228404
rect 115842 228352 115848 228404
rect 115900 228392 115906 228404
rect 115900 228364 122834 228392
rect 115900 228352 115906 228364
rect 122806 228324 122834 228364
rect 144730 228352 144736 228404
rect 144788 228392 144794 228404
rect 178034 228392 178040 228404
rect 144788 228364 178040 228392
rect 144788 228352 144794 228364
rect 178034 228352 178040 228364
rect 178092 228352 178098 228404
rect 224402 228352 224408 228404
rect 224460 228392 224466 228404
rect 327810 228392 327816 228404
rect 224460 228364 327816 228392
rect 224460 228352 224466 228364
rect 327810 228352 327816 228364
rect 327868 228352 327874 228404
rect 144086 228324 144092 228336
rect 122806 228296 144092 228324
rect 144086 228284 144092 228296
rect 144144 228284 144150 228336
rect 77202 227672 77208 227724
rect 77260 227712 77266 227724
rect 165154 227712 165160 227724
rect 77260 227684 165160 227712
rect 77260 227672 77266 227684
rect 165154 227672 165160 227684
rect 165212 227672 165218 227724
rect 190454 227672 190460 227724
rect 190512 227712 190518 227724
rect 268378 227712 268384 227724
rect 190512 227684 268384 227712
rect 190512 227672 190518 227684
rect 268378 227672 268384 227684
rect 268436 227672 268442 227724
rect 111702 227604 111708 227656
rect 111760 227644 111766 227656
rect 142154 227644 142160 227656
rect 111760 227616 142160 227644
rect 111760 227604 111766 227616
rect 142154 227604 142160 227616
rect 142212 227604 142218 227656
rect 221642 227604 221648 227656
rect 221700 227644 221706 227656
rect 276014 227644 276020 227656
rect 221700 227616 276020 227644
rect 221700 227604 221706 227616
rect 276014 227604 276020 227616
rect 276072 227604 276078 227656
rect 147674 226992 147680 227044
rect 147732 227032 147738 227044
rect 155218 227032 155224 227044
rect 147732 227004 155224 227032
rect 147732 226992 147738 227004
rect 155218 226992 155224 227004
rect 155276 226992 155282 227044
rect 177482 226992 177488 227044
rect 177540 227032 177546 227044
rect 221550 227032 221556 227044
rect 177540 227004 221556 227032
rect 177540 226992 177546 227004
rect 221550 226992 221556 227004
rect 221608 226992 221614 227044
rect 276014 226992 276020 227044
rect 276072 227032 276078 227044
rect 290090 227032 290096 227044
rect 276072 227004 290096 227032
rect 276072 226992 276078 227004
rect 290090 226992 290096 227004
rect 290148 226992 290154 227044
rect 154574 226312 154580 226364
rect 154632 226352 154638 226364
rect 156782 226352 156788 226364
rect 154632 226324 156788 226352
rect 154632 226312 154638 226324
rect 156782 226312 156788 226324
rect 156840 226312 156846 226364
rect 74534 226244 74540 226296
rect 74592 226284 74598 226296
rect 139118 226284 139124 226296
rect 74592 226256 139124 226284
rect 74592 226244 74598 226256
rect 139118 226244 139124 226256
rect 139176 226244 139182 226296
rect 139210 226244 139216 226296
rect 139268 226284 139274 226296
rect 147674 226284 147680 226296
rect 139268 226256 147680 226284
rect 139268 226244 139274 226256
rect 147674 226244 147680 226256
rect 147732 226244 147738 226296
rect 147766 226244 147772 226296
rect 147824 226284 147830 226296
rect 164878 226284 164884 226296
rect 147824 226256 164884 226284
rect 147824 226244 147830 226256
rect 164878 226244 164884 226256
rect 164936 226244 164942 226296
rect 181714 226244 181720 226296
rect 181772 226284 181778 226296
rect 247126 226284 247132 226296
rect 181772 226256 247132 226284
rect 181772 226244 181778 226256
rect 247126 226244 247132 226256
rect 247184 226244 247190 226296
rect 249794 225632 249800 225684
rect 249852 225672 249858 225684
rect 280154 225672 280160 225684
rect 249852 225644 280160 225672
rect 249852 225632 249858 225644
rect 280154 225632 280160 225644
rect 280212 225672 280218 225684
rect 290458 225672 290464 225684
rect 280212 225644 290464 225672
rect 280212 225632 280218 225644
rect 290458 225632 290464 225644
rect 290516 225632 290522 225684
rect 77294 225564 77300 225616
rect 77352 225604 77358 225616
rect 215938 225604 215944 225616
rect 77352 225576 215944 225604
rect 77352 225564 77358 225576
rect 215938 225564 215944 225576
rect 215996 225564 216002 225616
rect 238018 225564 238024 225616
rect 238076 225604 238082 225616
rect 296806 225604 296812 225616
rect 238076 225576 296812 225604
rect 238076 225564 238082 225576
rect 296806 225564 296812 225576
rect 296864 225604 296870 225616
rect 297358 225604 297364 225616
rect 296864 225576 297364 225604
rect 296864 225564 296870 225576
rect 297358 225564 297364 225576
rect 297416 225564 297422 225616
rect 305638 225564 305644 225616
rect 305696 225604 305702 225616
rect 334618 225604 334624 225616
rect 305696 225576 334624 225604
rect 305696 225564 305702 225576
rect 334618 225564 334624 225576
rect 334676 225564 334682 225616
rect 298462 224952 298468 225004
rect 298520 224992 298526 225004
rect 436094 224992 436100 225004
rect 298520 224964 436100 224992
rect 298520 224952 298526 224964
rect 436094 224952 436100 224964
rect 436152 224952 436158 225004
rect 140774 224272 140780 224324
rect 140832 224312 140838 224324
rect 211062 224312 211068 224324
rect 140832 224284 211068 224312
rect 140832 224272 140838 224284
rect 211062 224272 211068 224284
rect 211120 224312 211126 224324
rect 211430 224312 211436 224324
rect 211120 224284 211436 224312
rect 211120 224272 211126 224284
rect 211430 224272 211436 224284
rect 211488 224272 211494 224324
rect 67818 224204 67824 224256
rect 67876 224244 67882 224256
rect 142798 224244 142804 224256
rect 67876 224216 142804 224244
rect 67876 224204 67882 224216
rect 142798 224204 142804 224216
rect 142856 224204 142862 224256
rect 151722 224204 151728 224256
rect 151780 224244 151786 224256
rect 195238 224244 195244 224256
rect 151780 224216 195244 224244
rect 151780 224204 151786 224216
rect 195238 224204 195244 224216
rect 195296 224204 195302 224256
rect 200758 224204 200764 224256
rect 200816 224244 200822 224256
rect 202230 224244 202236 224256
rect 200816 224216 202236 224244
rect 200816 224204 200822 224216
rect 202230 224204 202236 224216
rect 202288 224204 202294 224256
rect 212442 224204 212448 224256
rect 212500 224244 212506 224256
rect 246114 224244 246120 224256
rect 212500 224216 246120 224244
rect 212500 224204 212506 224216
rect 246114 224204 246120 224216
rect 246172 224204 246178 224256
rect 148318 223524 148324 223576
rect 148376 223564 148382 223576
rect 154574 223564 154580 223576
rect 148376 223536 154580 223564
rect 148376 223524 148382 223536
rect 154574 223524 154580 223536
rect 154632 223564 154638 223576
rect 155218 223564 155224 223576
rect 154632 223536 155224 223564
rect 154632 223524 154638 223536
rect 155218 223524 155224 223536
rect 155276 223524 155282 223576
rect 174538 223524 174544 223576
rect 174596 223564 174602 223576
rect 224310 223564 224316 223576
rect 174596 223536 224316 223564
rect 174596 223524 174602 223536
rect 224310 223524 224316 223536
rect 224368 223564 224374 223576
rect 224862 223564 224868 223576
rect 224368 223536 224868 223564
rect 224368 223524 224374 223536
rect 224862 223524 224868 223536
rect 224920 223524 224926 223576
rect 132310 223456 132316 223508
rect 132368 223496 132374 223508
rect 181530 223496 181536 223508
rect 132368 223468 181536 223496
rect 132368 223456 132374 223468
rect 181530 223456 181536 223468
rect 181588 223456 181594 223508
rect 191190 223456 191196 223508
rect 191248 223496 191254 223508
rect 195698 223496 195704 223508
rect 191248 223468 195704 223496
rect 191248 223456 191254 223468
rect 195698 223456 195704 223468
rect 195756 223456 195762 223508
rect 297910 222844 297916 222896
rect 297968 222884 297974 222896
rect 349798 222884 349804 222896
rect 297968 222856 349804 222884
rect 297968 222844 297974 222856
rect 349798 222844 349804 222856
rect 349856 222844 349862 222896
rect 195422 222164 195428 222216
rect 195480 222204 195486 222216
rect 207934 222204 207940 222216
rect 195480 222176 207940 222204
rect 195480 222164 195486 222176
rect 207934 222164 207940 222176
rect 207992 222164 207998 222216
rect 130930 222096 130936 222148
rect 130988 222136 130994 222148
rect 163498 222136 163504 222148
rect 130988 222108 163504 222136
rect 130988 222096 130994 222108
rect 163498 222096 163504 222108
rect 163556 222136 163562 222148
rect 164142 222136 164148 222148
rect 163556 222108 164148 222136
rect 163556 222096 163562 222108
rect 164142 222096 164148 222108
rect 164200 222096 164206 222148
rect 195238 222096 195244 222148
rect 195296 222136 195302 222148
rect 240870 222136 240876 222148
rect 195296 222108 240876 222136
rect 195296 222096 195302 222108
rect 240870 222096 240876 222108
rect 240928 222096 240934 222148
rect 164142 221484 164148 221536
rect 164200 221524 164206 221536
rect 195238 221524 195244 221536
rect 164200 221496 195244 221524
rect 164200 221484 164206 221496
rect 195238 221484 195244 221496
rect 195296 221484 195302 221536
rect 269022 221484 269028 221536
rect 269080 221524 269086 221536
rect 342898 221524 342904 221536
rect 269080 221496 342904 221524
rect 269080 221484 269086 221496
rect 342898 221484 342904 221496
rect 342956 221484 342962 221536
rect 194318 221416 194324 221468
rect 194376 221456 194382 221468
rect 273898 221456 273904 221468
rect 194376 221428 273904 221456
rect 194376 221416 194382 221428
rect 273898 221416 273904 221428
rect 273956 221416 273962 221468
rect 320634 221416 320640 221468
rect 320692 221456 320698 221468
rect 454034 221456 454040 221468
rect 320692 221428 454040 221456
rect 320692 221416 320698 221428
rect 454034 221416 454040 221428
rect 454092 221416 454098 221468
rect 276750 220804 276756 220856
rect 276808 220844 276814 220856
rect 277394 220844 277400 220856
rect 276808 220816 277400 220844
rect 276808 220804 276814 220816
rect 277394 220804 277400 220816
rect 277452 220804 277458 220856
rect 59170 220736 59176 220788
rect 59228 220776 59234 220788
rect 217134 220776 217140 220788
rect 59228 220748 217140 220776
rect 59228 220736 59234 220748
rect 217134 220736 217140 220748
rect 217192 220736 217198 220788
rect 195698 220668 195704 220720
rect 195756 220708 195762 220720
rect 212442 220708 212448 220720
rect 195756 220680 212448 220708
rect 195756 220668 195762 220680
rect 212442 220668 212448 220680
rect 212500 220668 212506 220720
rect 60458 220056 60464 220108
rect 60516 220096 60522 220108
rect 60516 220068 142154 220096
rect 60516 220056 60522 220068
rect 142126 220028 142154 220068
rect 156506 220056 156512 220108
rect 156564 220096 156570 220108
rect 192938 220096 192944 220108
rect 156564 220068 192944 220096
rect 156564 220056 156570 220068
rect 192938 220056 192944 220068
rect 192996 220056 193002 220108
rect 238754 220056 238760 220108
rect 238812 220096 238818 220108
rect 272702 220096 272708 220108
rect 238812 220068 272708 220096
rect 238812 220056 238818 220068
rect 272702 220056 272708 220068
rect 272760 220056 272766 220108
rect 156690 220028 156696 220040
rect 142126 220000 156696 220028
rect 156690 219988 156696 220000
rect 156748 219988 156754 220040
rect 211982 219444 211988 219496
rect 212040 219484 212046 219496
rect 325050 219484 325056 219496
rect 212040 219456 325056 219484
rect 212040 219444 212046 219456
rect 325050 219444 325056 219456
rect 325108 219444 325114 219496
rect 73798 219376 73804 219428
rect 73856 219416 73862 219428
rect 184290 219416 184296 219428
rect 73856 219388 184296 219416
rect 73856 219376 73862 219388
rect 184290 219376 184296 219388
rect 184348 219376 184354 219428
rect 195882 219376 195888 219428
rect 195940 219416 195946 219428
rect 270494 219416 270500 219428
rect 195940 219388 270500 219416
rect 195940 219376 195946 219388
rect 270494 219376 270500 219388
rect 270552 219376 270558 219428
rect 126974 219308 126980 219360
rect 127032 219348 127038 219360
rect 217318 219348 217324 219360
rect 127032 219320 217324 219348
rect 127032 219308 127038 219320
rect 217318 219308 217324 219320
rect 217376 219308 217382 219360
rect 221366 219308 221372 219360
rect 221424 219348 221430 219360
rect 263778 219348 263784 219360
rect 221424 219320 263784 219348
rect 221424 219308 221430 219320
rect 263778 219308 263784 219320
rect 263836 219308 263842 219360
rect 267090 218696 267096 218748
rect 267148 218736 267154 218748
rect 275370 218736 275376 218748
rect 267148 218708 275376 218736
rect 267148 218696 267154 218708
rect 275370 218696 275376 218708
rect 275428 218696 275434 218748
rect 192662 218016 192668 218068
rect 192720 218056 192726 218068
rect 195238 218056 195244 218068
rect 192720 218028 195244 218056
rect 192720 218016 192726 218028
rect 195238 218016 195244 218028
rect 195296 218016 195302 218068
rect 270494 218016 270500 218068
rect 270552 218056 270558 218068
rect 271138 218056 271144 218068
rect 270552 218028 271144 218056
rect 270552 218016 270558 218028
rect 271138 218016 271144 218028
rect 271196 218016 271202 218068
rect 83550 217948 83556 218000
rect 83608 217988 83614 218000
rect 201494 217988 201500 218000
rect 83608 217960 201500 217988
rect 83608 217948 83614 217960
rect 201494 217948 201500 217960
rect 201552 217988 201558 218000
rect 202046 217988 202052 218000
rect 201552 217960 202052 217988
rect 201552 217948 201558 217960
rect 202046 217948 202052 217960
rect 202104 217948 202110 218000
rect 202322 217948 202328 218000
rect 202380 217988 202386 218000
rect 231118 217988 231124 218000
rect 202380 217960 231124 217988
rect 202380 217948 202386 217960
rect 231118 217948 231124 217960
rect 231176 217948 231182 218000
rect 193030 217676 193036 217728
rect 193088 217716 193094 217728
rect 198090 217716 198096 217728
rect 193088 217688 198096 217716
rect 193088 217676 193094 217688
rect 198090 217676 198096 217688
rect 198148 217676 198154 217728
rect 202046 217336 202052 217388
rect 202104 217376 202110 217388
rect 285674 217376 285680 217388
rect 202104 217348 285680 217376
rect 202104 217336 202110 217348
rect 285674 217336 285680 217348
rect 285732 217336 285738 217388
rect 82722 217268 82728 217320
rect 82780 217308 82786 217320
rect 158714 217308 158720 217320
rect 82780 217280 158720 217308
rect 82780 217268 82786 217280
rect 158714 217268 158720 217280
rect 158772 217268 158778 217320
rect 235350 217268 235356 217320
rect 235408 217308 235414 217320
rect 388530 217308 388536 217320
rect 235408 217280 388536 217308
rect 235408 217268 235414 217280
rect 388530 217268 388536 217280
rect 388588 217268 388594 217320
rect 197998 216656 198004 216708
rect 198056 216696 198062 216708
rect 198734 216696 198740 216708
rect 198056 216668 198740 216696
rect 198056 216656 198062 216668
rect 198734 216656 198740 216668
rect 198792 216656 198798 216708
rect 69750 216588 69756 216640
rect 69808 216628 69814 216640
rect 233510 216628 233516 216640
rect 69808 216600 233516 216628
rect 69808 216588 69814 216600
rect 233510 216588 233516 216600
rect 233568 216588 233574 216640
rect 132402 216520 132408 216572
rect 132460 216560 132466 216572
rect 195330 216560 195336 216572
rect 132460 216532 195336 216560
rect 132460 216520 132466 216532
rect 195330 216520 195336 216532
rect 195388 216520 195394 216572
rect 214558 216520 214564 216572
rect 214616 216560 214622 216572
rect 248966 216560 248972 216572
rect 214616 216532 248972 216560
rect 214616 216520 214622 216532
rect 248966 216520 248972 216532
rect 249024 216560 249030 216572
rect 249702 216560 249708 216572
rect 249024 216532 249708 216560
rect 249024 216520 249030 216532
rect 249702 216520 249708 216532
rect 249760 216520 249766 216572
rect 233510 216044 233516 216096
rect 233568 216084 233574 216096
rect 234430 216084 234436 216096
rect 233568 216056 234436 216084
rect 233568 216044 233574 216056
rect 234430 216044 234436 216056
rect 234488 216044 234494 216096
rect 249702 215908 249708 215960
rect 249760 215948 249766 215960
rect 456794 215948 456800 215960
rect 249760 215920 456800 215948
rect 249760 215908 249766 215920
rect 456794 215908 456800 215920
rect 456852 215908 456858 215960
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 39298 215268 39304 215280
rect 3384 215240 39304 215268
rect 3384 215228 3390 215240
rect 39298 215228 39304 215240
rect 39356 215228 39362 215280
rect 124214 215228 124220 215280
rect 124272 215268 124278 215280
rect 222378 215268 222384 215280
rect 124272 215240 222384 215268
rect 124272 215228 124278 215240
rect 222378 215228 222384 215240
rect 222436 215268 222442 215280
rect 223390 215268 223396 215280
rect 222436 215240 223396 215268
rect 222436 215228 222442 215240
rect 223390 215228 223396 215240
rect 223448 215228 223454 215280
rect 141970 215160 141976 215212
rect 142028 215200 142034 215212
rect 168374 215200 168380 215212
rect 142028 215172 168380 215200
rect 142028 215160 142034 215172
rect 168374 215160 168380 215172
rect 168432 215160 168438 215212
rect 67634 214548 67640 214600
rect 67692 214588 67698 214600
rect 133138 214588 133144 214600
rect 67692 214560 133144 214588
rect 67692 214548 67698 214560
rect 133138 214548 133144 214560
rect 133196 214548 133202 214600
rect 168374 214548 168380 214600
rect 168432 214588 168438 214600
rect 169570 214588 169576 214600
rect 168432 214560 169576 214588
rect 168432 214548 168438 214560
rect 169570 214548 169576 214560
rect 169628 214588 169634 214600
rect 217410 214588 217416 214600
rect 169628 214560 217416 214588
rect 169628 214548 169634 214560
rect 217410 214548 217416 214560
rect 217468 214548 217474 214600
rect 431862 214548 431868 214600
rect 431920 214588 431926 214600
rect 434714 214588 434720 214600
rect 431920 214560 434720 214588
rect 431920 214548 431926 214560
rect 434714 214548 434720 214560
rect 434772 214548 434778 214600
rect 223390 213936 223396 213988
rect 223448 213976 223454 213988
rect 231946 213976 231952 213988
rect 223448 213948 231952 213976
rect 223448 213936 223454 213948
rect 231946 213936 231952 213948
rect 232004 213936 232010 213988
rect 81434 213868 81440 213920
rect 81492 213908 81498 213920
rect 191098 213908 191104 213920
rect 81492 213880 191104 213908
rect 81492 213868 81498 213880
rect 191098 213868 191104 213880
rect 191156 213868 191162 213920
rect 213454 213868 213460 213920
rect 213512 213908 213518 213920
rect 299566 213908 299572 213920
rect 213512 213880 299572 213908
rect 213512 213868 213518 213880
rect 299566 213868 299572 213880
rect 299624 213908 299630 213920
rect 300210 213908 300216 213920
rect 299624 213880 300216 213908
rect 299624 213868 299630 213880
rect 300210 213868 300216 213880
rect 300268 213868 300274 213920
rect 147490 213800 147496 213852
rect 147548 213840 147554 213852
rect 244458 213840 244464 213852
rect 147548 213812 244464 213840
rect 147548 213800 147554 213812
rect 244458 213800 244464 213812
rect 244516 213800 244522 213852
rect 196710 213188 196716 213240
rect 196768 213228 196774 213240
rect 212534 213228 212540 213240
rect 196768 213200 212540 213228
rect 196768 213188 196774 213200
rect 212534 213188 212540 213200
rect 212592 213228 212598 213240
rect 213454 213228 213460 213240
rect 212592 213200 213460 213228
rect 212592 213188 212598 213200
rect 213454 213188 213460 213200
rect 213512 213188 213518 213240
rect 254026 213188 254032 213240
rect 254084 213228 254090 213240
rect 389818 213228 389824 213240
rect 254084 213200 389824 213228
rect 254084 213188 254090 213200
rect 389818 213188 389824 213200
rect 389876 213188 389882 213240
rect 64598 212440 64604 212492
rect 64656 212480 64662 212492
rect 206462 212480 206468 212492
rect 64656 212452 206468 212480
rect 64656 212440 64662 212452
rect 206462 212440 206468 212452
rect 206520 212440 206526 212492
rect 136634 212372 136640 212424
rect 136692 212412 136698 212424
rect 240134 212412 240140 212424
rect 136692 212384 240140 212412
rect 136692 212372 136698 212384
rect 240134 212372 240140 212384
rect 240192 212412 240198 212424
rect 240778 212412 240784 212424
rect 240192 212384 240784 212412
rect 240192 212372 240198 212384
rect 240778 212372 240784 212384
rect 240836 212372 240842 212424
rect 162762 211080 162768 211132
rect 162820 211120 162826 211132
rect 163682 211120 163688 211132
rect 162820 211092 163688 211120
rect 162820 211080 162826 211092
rect 163682 211080 163688 211092
rect 163740 211080 163746 211132
rect 192478 211080 192484 211132
rect 192536 211120 192542 211132
rect 259454 211120 259460 211132
rect 192536 211092 259460 211120
rect 192536 211080 192542 211092
rect 259454 211080 259460 211092
rect 259512 211120 259518 211132
rect 260742 211120 260748 211132
rect 259512 211092 260748 211120
rect 259512 211080 259518 211092
rect 260742 211080 260748 211092
rect 260800 211080 260806 211132
rect 212534 211012 212540 211064
rect 212592 211052 212598 211064
rect 213638 211052 213644 211064
rect 212592 211024 213644 211052
rect 212592 211012 212598 211024
rect 213638 211012 213644 211024
rect 213696 211012 213702 211064
rect 218422 211012 218428 211064
rect 218480 211052 218486 211064
rect 218790 211052 218796 211064
rect 218480 211024 218796 211052
rect 218480 211012 218486 211024
rect 218790 211012 218796 211024
rect 218848 211052 218854 211064
rect 274634 211052 274640 211064
rect 218848 211024 274640 211052
rect 218848 211012 218854 211024
rect 274634 211012 274640 211024
rect 274692 211012 274698 211064
rect 124306 210468 124312 210520
rect 124364 210508 124370 210520
rect 162762 210508 162768 210520
rect 124364 210480 162768 210508
rect 124364 210468 124370 210480
rect 162762 210468 162768 210480
rect 162820 210468 162826 210520
rect 274634 210468 274640 210520
rect 274692 210508 274698 210520
rect 289998 210508 290004 210520
rect 274692 210480 290004 210508
rect 274692 210468 274698 210480
rect 289998 210468 290004 210480
rect 290056 210468 290062 210520
rect 72510 210400 72516 210452
rect 72568 210440 72574 210452
rect 182174 210440 182180 210452
rect 72568 210412 182180 210440
rect 72568 210400 72574 210412
rect 182174 210400 182180 210412
rect 182232 210400 182238 210452
rect 187050 210400 187056 210452
rect 187108 210440 187114 210452
rect 212534 210440 212540 210452
rect 187108 210412 212540 210440
rect 187108 210400 187114 210412
rect 212534 210400 212540 210412
rect 212592 210400 212598 210452
rect 260742 210400 260748 210452
rect 260800 210440 260806 210452
rect 356698 210440 356704 210452
rect 260800 210412 356704 210440
rect 260800 210400 260806 210412
rect 356698 210400 356704 210412
rect 356756 210400 356762 210452
rect 106182 209720 106188 209772
rect 106240 209760 106246 209772
rect 216766 209760 216772 209772
rect 106240 209732 216772 209760
rect 106240 209720 106246 209732
rect 216766 209720 216772 209732
rect 216824 209720 216830 209772
rect 63402 209652 63408 209704
rect 63460 209692 63466 209704
rect 173802 209692 173808 209704
rect 63460 209664 173808 209692
rect 63460 209652 63466 209664
rect 173802 209652 173808 209664
rect 173860 209652 173866 209704
rect 223390 209108 223396 209160
rect 223448 209148 223454 209160
rect 282270 209148 282276 209160
rect 223448 209120 282276 209148
rect 223448 209108 223454 209120
rect 282270 209108 282276 209120
rect 282328 209108 282334 209160
rect 217410 209040 217416 209092
rect 217468 209080 217474 209092
rect 237466 209080 237472 209092
rect 217468 209052 237472 209080
rect 217468 209040 217474 209052
rect 237466 209040 237472 209052
rect 237524 209040 237530 209092
rect 242158 209040 242164 209092
rect 242216 209080 242222 209092
rect 251910 209080 251916 209092
rect 242216 209052 251916 209080
rect 242216 209040 242222 209052
rect 251910 209040 251916 209052
rect 251968 209040 251974 209092
rect 272702 209040 272708 209092
rect 272760 209080 272766 209092
rect 438118 209080 438124 209092
rect 272760 209052 438124 209080
rect 272760 209040 272766 209052
rect 438118 209040 438124 209052
rect 438176 209040 438182 209092
rect 95142 208292 95148 208344
rect 95200 208332 95206 208344
rect 193858 208332 193864 208344
rect 95200 208304 193864 208332
rect 95200 208292 95206 208304
rect 193858 208292 193864 208304
rect 193916 208292 193922 208344
rect 203518 208020 203524 208072
rect 203576 208060 203582 208072
rect 211890 208060 211896 208072
rect 203576 208032 211896 208060
rect 203576 208020 203582 208032
rect 211890 208020 211896 208032
rect 211948 208020 211954 208072
rect 212442 207680 212448 207732
rect 212500 207720 212506 207732
rect 235258 207720 235264 207732
rect 212500 207692 235264 207720
rect 212500 207680 212506 207692
rect 235258 207680 235264 207692
rect 235316 207680 235322 207732
rect 93946 207612 93952 207664
rect 94004 207652 94010 207664
rect 95142 207652 95148 207664
rect 94004 207624 95148 207652
rect 94004 207612 94010 207624
rect 95142 207612 95148 207624
rect 95200 207612 95206 207664
rect 133782 207612 133788 207664
rect 133840 207652 133846 207664
rect 229186 207652 229192 207664
rect 133840 207624 229192 207652
rect 133840 207612 133846 207624
rect 229186 207612 229192 207624
rect 229244 207652 229250 207664
rect 245838 207652 245844 207664
rect 229244 207624 245844 207652
rect 229244 207612 229250 207624
rect 245838 207612 245844 207624
rect 245896 207612 245902 207664
rect 250530 207612 250536 207664
rect 250588 207652 250594 207664
rect 308398 207652 308404 207664
rect 250588 207624 308404 207652
rect 250588 207612 250594 207624
rect 308398 207612 308404 207624
rect 308456 207612 308462 207664
rect 114462 206932 114468 206984
rect 114520 206972 114526 206984
rect 242894 206972 242900 206984
rect 114520 206944 242900 206972
rect 114520 206932 114526 206944
rect 242894 206932 242900 206944
rect 242952 206932 242958 206984
rect 440234 206932 440240 206984
rect 440292 206972 440298 206984
rect 440878 206972 440884 206984
rect 440292 206944 440884 206972
rect 440292 206932 440298 206944
rect 440878 206932 440884 206944
rect 440936 206972 440942 206984
rect 582742 206972 582748 206984
rect 440936 206944 582748 206972
rect 440936 206932 440942 206944
rect 582742 206932 582748 206944
rect 582800 206932 582806 206984
rect 105538 206864 105544 206916
rect 105596 206904 105602 206916
rect 214466 206904 214472 206916
rect 105596 206876 214472 206904
rect 105596 206864 105602 206876
rect 214466 206864 214472 206876
rect 214524 206864 214530 206916
rect 264974 206252 264980 206304
rect 265032 206292 265038 206304
rect 371878 206292 371884 206304
rect 265032 206264 371884 206292
rect 265032 206252 265038 206264
rect 371878 206252 371884 206264
rect 371936 206252 371942 206304
rect 242894 206116 242900 206168
rect 242952 206156 242958 206168
rect 243906 206156 243912 206168
rect 242952 206128 243912 206156
rect 242952 206116 242958 206128
rect 243906 206116 243912 206128
rect 243964 206116 243970 206168
rect 214466 205640 214472 205692
rect 214524 205680 214530 205692
rect 216030 205680 216036 205692
rect 214524 205652 216036 205680
rect 214524 205640 214530 205652
rect 216030 205640 216036 205652
rect 216088 205640 216094 205692
rect 216122 205640 216128 205692
rect 216180 205680 216186 205692
rect 216490 205680 216496 205692
rect 216180 205652 216496 205680
rect 216180 205640 216186 205652
rect 216490 205640 216496 205652
rect 216548 205680 216554 205692
rect 245838 205680 245844 205692
rect 216548 205652 245844 205680
rect 216548 205640 216554 205652
rect 245838 205640 245844 205652
rect 245896 205640 245902 205692
rect 97258 205572 97264 205624
rect 97316 205612 97322 205624
rect 205818 205612 205824 205624
rect 97316 205584 205824 205612
rect 97316 205572 97322 205584
rect 205818 205572 205824 205584
rect 205876 205572 205882 205624
rect 205818 205096 205824 205148
rect 205876 205136 205882 205148
rect 206554 205136 206560 205148
rect 205876 205108 206560 205136
rect 205876 205096 205882 205108
rect 206554 205096 206560 205108
rect 206612 205096 206618 205148
rect 87138 204892 87144 204944
rect 87196 204932 87202 204944
rect 184658 204932 184664 204944
rect 87196 204904 184664 204932
rect 87196 204892 87202 204904
rect 184658 204892 184664 204904
rect 184716 204932 184722 204944
rect 185578 204932 185584 204944
rect 184716 204904 185584 204932
rect 184716 204892 184722 204904
rect 185578 204892 185584 204904
rect 185636 204892 185642 204944
rect 207290 204892 207296 204944
rect 207348 204932 207354 204944
rect 280890 204932 280896 204944
rect 207348 204904 280896 204932
rect 207348 204892 207354 204904
rect 280890 204892 280896 204904
rect 280948 204892 280954 204944
rect 207014 204280 207020 204332
rect 207072 204320 207078 204332
rect 207382 204320 207388 204332
rect 207072 204292 207388 204320
rect 207072 204280 207078 204292
rect 207382 204280 207388 204292
rect 207440 204320 207446 204332
rect 215294 204320 215300 204332
rect 207440 204292 215300 204320
rect 207440 204280 207446 204292
rect 215294 204280 215300 204292
rect 215352 204280 215358 204332
rect 70394 204212 70400 204264
rect 70452 204252 70458 204264
rect 216122 204252 216128 204264
rect 70452 204224 216128 204252
rect 70452 204212 70458 204224
rect 216122 204212 216128 204224
rect 216180 204212 216186 204264
rect 184750 203600 184756 203652
rect 184808 203640 184814 203652
rect 227714 203640 227720 203652
rect 184808 203612 227720 203640
rect 184808 203600 184814 203612
rect 227714 203600 227720 203612
rect 227772 203600 227778 203652
rect 102042 203532 102048 203584
rect 102100 203572 102106 203584
rect 171778 203572 171784 203584
rect 102100 203544 171784 203572
rect 102100 203532 102106 203544
rect 171778 203532 171784 203544
rect 171836 203532 171842 203584
rect 215294 203532 215300 203584
rect 215352 203572 215358 203584
rect 284938 203572 284944 203584
rect 215352 203544 284944 203572
rect 215352 203532 215358 203544
rect 284938 203532 284944 203544
rect 284996 203532 285002 203584
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 128998 202824 129004 202836
rect 3108 202796 129004 202824
rect 3108 202784 3114 202796
rect 128998 202784 129004 202796
rect 129056 202784 129062 202836
rect 156690 202784 156696 202836
rect 156748 202824 156754 202836
rect 177758 202824 177764 202836
rect 156748 202796 177764 202824
rect 156748 202784 156754 202796
rect 177758 202784 177764 202796
rect 177816 202824 177822 202836
rect 207014 202824 207020 202836
rect 177816 202796 207020 202824
rect 177816 202784 177822 202796
rect 207014 202784 207020 202796
rect 207072 202784 207078 202836
rect 126882 202716 126888 202768
rect 126940 202756 126946 202768
rect 248506 202756 248512 202768
rect 126940 202728 248512 202756
rect 126940 202716 126946 202728
rect 248506 202716 248512 202728
rect 248564 202716 248570 202768
rect 211062 202104 211068 202156
rect 211120 202144 211126 202156
rect 240226 202144 240232 202156
rect 211120 202116 240232 202144
rect 211120 202104 211126 202116
rect 240226 202104 240232 202116
rect 240284 202104 240290 202156
rect 273990 201764 273996 201816
rect 274048 201804 274054 201816
rect 278222 201804 278228 201816
rect 274048 201776 278228 201804
rect 274048 201764 274054 201776
rect 278222 201764 278228 201776
rect 278280 201764 278286 201816
rect 97902 201424 97908 201476
rect 97960 201464 97966 201476
rect 165062 201464 165068 201476
rect 97960 201436 165068 201464
rect 97960 201424 97966 201436
rect 165062 201424 165068 201436
rect 165120 201424 165126 201476
rect 168282 201424 168288 201476
rect 168340 201464 168346 201476
rect 211982 201464 211988 201476
rect 168340 201436 211988 201464
rect 168340 201424 168346 201436
rect 211982 201424 211988 201436
rect 212040 201424 212046 201476
rect 195330 200812 195336 200864
rect 195388 200852 195394 200864
rect 218698 200852 218704 200864
rect 195388 200824 218704 200852
rect 195388 200812 195394 200824
rect 218698 200812 218704 200824
rect 218756 200812 218762 200864
rect 224310 200812 224316 200864
rect 224368 200852 224374 200864
rect 235994 200852 236000 200864
rect 224368 200824 236000 200852
rect 224368 200812 224374 200824
rect 235994 200812 236000 200824
rect 236052 200812 236058 200864
rect 122742 200744 122748 200796
rect 122800 200784 122806 200796
rect 178770 200784 178776 200796
rect 122800 200756 178776 200784
rect 122800 200744 122806 200756
rect 178770 200744 178776 200756
rect 178828 200744 178834 200796
rect 214650 200744 214656 200796
rect 214708 200784 214714 200796
rect 306466 200784 306472 200796
rect 214708 200756 306472 200784
rect 214708 200744 214714 200756
rect 306466 200744 306472 200756
rect 306524 200744 306530 200796
rect 323670 200744 323676 200796
rect 323728 200784 323734 200796
rect 431218 200784 431224 200796
rect 323728 200756 431224 200784
rect 323728 200744 323734 200756
rect 431218 200744 431224 200756
rect 431276 200744 431282 200796
rect 79962 200064 79968 200116
rect 80020 200104 80026 200116
rect 194502 200104 194508 200116
rect 80020 200076 194508 200104
rect 80020 200064 80026 200076
rect 194502 200064 194508 200076
rect 194560 200064 194566 200116
rect 194410 199452 194416 199504
rect 194468 199492 194474 199504
rect 287238 199492 287244 199504
rect 194468 199464 287244 199492
rect 194468 199452 194474 199464
rect 287238 199452 287244 199464
rect 287296 199452 287302 199504
rect 54938 199384 54944 199436
rect 54996 199424 55002 199436
rect 177850 199424 177856 199436
rect 54996 199396 177856 199424
rect 54996 199384 55002 199396
rect 177850 199384 177856 199396
rect 177908 199424 177914 199436
rect 178862 199424 178868 199436
rect 177908 199396 178868 199424
rect 177908 199384 177914 199396
rect 178862 199384 178868 199396
rect 178920 199384 178926 199436
rect 194502 199384 194508 199436
rect 194560 199424 194566 199436
rect 217318 199424 217324 199436
rect 194560 199396 217324 199424
rect 194560 199384 194566 199396
rect 217318 199384 217324 199396
rect 217376 199384 217382 199436
rect 239398 199384 239404 199436
rect 239456 199424 239462 199436
rect 385770 199424 385776 199436
rect 239456 199396 385776 199424
rect 239456 199384 239462 199396
rect 385770 199384 385776 199396
rect 385828 199384 385834 199436
rect 53558 198636 53564 198688
rect 53616 198676 53622 198688
rect 168282 198676 168288 198688
rect 53616 198648 168288 198676
rect 53616 198636 53622 198648
rect 168282 198636 168288 198648
rect 168340 198636 168346 198688
rect 178954 198636 178960 198688
rect 179012 198676 179018 198688
rect 195238 198676 195244 198688
rect 179012 198648 195244 198676
rect 179012 198636 179018 198648
rect 195238 198636 195244 198648
rect 195296 198636 195302 198688
rect 139394 198568 139400 198620
rect 139452 198608 139458 198620
rect 166902 198608 166908 198620
rect 139452 198580 166908 198608
rect 139452 198568 139458 198580
rect 166902 198568 166908 198580
rect 166960 198568 166966 198620
rect 195422 198024 195428 198076
rect 195480 198064 195486 198076
rect 206278 198064 206284 198076
rect 195480 198036 206284 198064
rect 195480 198024 195486 198036
rect 206278 198024 206284 198036
rect 206336 198024 206342 198076
rect 206554 198024 206560 198076
rect 206612 198064 206618 198076
rect 288618 198064 288624 198076
rect 206612 198036 288624 198064
rect 206612 198024 206618 198036
rect 288618 198024 288624 198036
rect 288676 198024 288682 198076
rect 166166 197956 166172 198008
rect 166224 197996 166230 198008
rect 218790 197996 218796 198008
rect 166224 197968 218796 197996
rect 166224 197956 166230 197968
rect 218790 197956 218796 197968
rect 218848 197956 218854 198008
rect 220354 197956 220360 198008
rect 220412 197996 220418 198008
rect 407114 197996 407120 198008
rect 220412 197968 407120 197996
rect 220412 197956 220418 197968
rect 407114 197956 407120 197968
rect 407172 197956 407178 198008
rect 64782 197276 64788 197328
rect 64840 197316 64846 197328
rect 221642 197316 221648 197328
rect 64840 197288 221648 197316
rect 64840 197276 64846 197288
rect 221642 197276 221648 197288
rect 221700 197276 221706 197328
rect 221550 196664 221556 196716
rect 221608 196704 221614 196716
rect 244366 196704 244372 196716
rect 221608 196676 244372 196704
rect 221608 196664 221614 196676
rect 244366 196664 244372 196676
rect 244424 196664 244430 196716
rect 135162 196596 135168 196648
rect 135220 196636 135226 196648
rect 181622 196636 181628 196648
rect 135220 196608 181628 196636
rect 135220 196596 135226 196608
rect 181622 196596 181628 196608
rect 181680 196596 181686 196648
rect 189718 196596 189724 196648
rect 189776 196636 189782 196648
rect 250438 196636 250444 196648
rect 189776 196608 250444 196636
rect 189776 196596 189782 196608
rect 250438 196596 250444 196608
rect 250496 196596 250502 196648
rect 251910 196596 251916 196648
rect 251968 196636 251974 196648
rect 300302 196636 300308 196648
rect 251968 196608 300308 196636
rect 251968 196596 251974 196608
rect 300302 196596 300308 196608
rect 300360 196596 300366 196648
rect 155218 195916 155224 195968
rect 155276 195956 155282 195968
rect 163498 195956 163504 195968
rect 155276 195928 163504 195956
rect 155276 195916 155282 195928
rect 163498 195916 163504 195928
rect 163556 195916 163562 195968
rect 163590 195304 163596 195356
rect 163648 195344 163654 195356
rect 176010 195344 176016 195356
rect 163648 195316 176016 195344
rect 163648 195304 163654 195316
rect 176010 195304 176016 195316
rect 176068 195304 176074 195356
rect 177850 195304 177856 195356
rect 177908 195344 177914 195356
rect 206554 195344 206560 195356
rect 177908 195316 206560 195344
rect 177908 195304 177914 195316
rect 206554 195304 206560 195316
rect 206612 195304 206618 195356
rect 280798 195304 280804 195356
rect 280856 195344 280862 195356
rect 303890 195344 303896 195356
rect 280856 195316 303896 195344
rect 280856 195304 280862 195316
rect 303890 195304 303896 195316
rect 303948 195304 303954 195356
rect 89622 195236 89628 195288
rect 89680 195276 89686 195288
rect 166350 195276 166356 195288
rect 89680 195248 166356 195276
rect 89680 195236 89686 195248
rect 166350 195236 166356 195248
rect 166408 195236 166414 195288
rect 206462 195236 206468 195288
rect 206520 195276 206526 195288
rect 241606 195276 241612 195288
rect 206520 195248 241612 195276
rect 206520 195236 206526 195248
rect 241606 195236 241612 195248
rect 241664 195236 241670 195288
rect 270402 195236 270408 195288
rect 270460 195276 270466 195288
rect 302234 195276 302240 195288
rect 270460 195248 302240 195276
rect 270460 195236 270466 195248
rect 302234 195236 302240 195248
rect 302292 195236 302298 195288
rect 61838 194488 61844 194540
rect 61896 194528 61902 194540
rect 220170 194528 220176 194540
rect 61896 194500 220176 194528
rect 61896 194488 61902 194500
rect 220170 194488 220176 194500
rect 220228 194488 220234 194540
rect 223482 193876 223488 193928
rect 223540 193916 223546 193928
rect 238754 193916 238760 193928
rect 223540 193888 238760 193916
rect 223540 193876 223546 193888
rect 238754 193876 238760 193888
rect 238812 193876 238818 193928
rect 144822 193808 144828 193860
rect 144880 193848 144886 193860
rect 163590 193848 163596 193860
rect 144880 193820 163596 193848
rect 144880 193808 144886 193820
rect 163590 193808 163596 193820
rect 163648 193808 163654 193860
rect 198090 193808 198096 193860
rect 198148 193848 198154 193860
rect 227070 193848 227076 193860
rect 198148 193820 227076 193848
rect 198148 193808 198154 193820
rect 227070 193808 227076 193820
rect 227128 193808 227134 193860
rect 395890 193808 395896 193860
rect 395948 193848 395954 193860
rect 582926 193848 582932 193860
rect 395948 193820 582932 193848
rect 395948 193808 395954 193820
rect 582926 193808 582932 193820
rect 582984 193808 582990 193860
rect 226334 193196 226340 193248
rect 226392 193236 226398 193248
rect 432690 193236 432696 193248
rect 226392 193208 432696 193236
rect 226392 193196 226398 193208
rect 432690 193196 432696 193208
rect 432748 193196 432754 193248
rect 57606 193128 57612 193180
rect 57664 193168 57670 193180
rect 166166 193168 166172 193180
rect 57664 193140 166172 193168
rect 57664 193128 57670 193140
rect 166166 193128 166172 193140
rect 166224 193128 166230 193180
rect 93118 193060 93124 193112
rect 93176 193100 93182 193112
rect 196710 193100 196716 193112
rect 93176 193072 196716 193100
rect 93176 193060 93182 193072
rect 196710 193060 196716 193072
rect 196768 193060 196774 193112
rect 202138 192516 202144 192568
rect 202196 192556 202202 192568
rect 239398 192556 239404 192568
rect 202196 192528 239404 192556
rect 202196 192516 202202 192528
rect 239398 192516 239404 192528
rect 239456 192516 239462 192568
rect 185670 192448 185676 192500
rect 185728 192488 185734 192500
rect 230658 192488 230664 192500
rect 185728 192460 230664 192488
rect 185728 192448 185734 192460
rect 230658 192448 230664 192460
rect 230716 192448 230722 192500
rect 400858 192448 400864 192500
rect 400916 192488 400922 192500
rect 415394 192488 415400 192500
rect 400916 192460 415400 192488
rect 400916 192448 400922 192460
rect 415394 192448 415400 192460
rect 415452 192448 415458 192500
rect 200022 192380 200028 192432
rect 200080 192420 200086 192432
rect 201494 192420 201500 192432
rect 200080 192392 201500 192420
rect 200080 192380 200086 192392
rect 201494 192380 201500 192392
rect 201552 192380 201558 192432
rect 156598 191768 156604 191820
rect 156656 191808 156662 191820
rect 226334 191808 226340 191820
rect 156656 191780 226340 191808
rect 156656 191768 156662 191780
rect 226334 191768 226340 191780
rect 226392 191768 226398 191820
rect 221458 191088 221464 191140
rect 221516 191128 221522 191140
rect 447318 191128 447324 191140
rect 221516 191100 447324 191128
rect 221516 191088 221522 191100
rect 447318 191088 447324 191100
rect 447376 191088 447382 191140
rect 118602 190476 118608 190528
rect 118660 190516 118666 190528
rect 170490 190516 170496 190528
rect 118660 190488 170496 190516
rect 118660 190476 118666 190488
rect 170490 190476 170496 190488
rect 170548 190476 170554 190528
rect 159358 190408 159364 190460
rect 159416 190448 159422 190460
rect 225598 190448 225604 190460
rect 159416 190420 225604 190448
rect 159416 190408 159422 190420
rect 225598 190408 225604 190420
rect 225656 190408 225662 190460
rect 264238 189728 264244 189780
rect 264296 189768 264302 189780
rect 281626 189768 281632 189780
rect 264296 189740 281632 189768
rect 264296 189728 264302 189740
rect 281626 189728 281632 189740
rect 281684 189728 281690 189780
rect 122742 189048 122748 189100
rect 122800 189088 122806 189100
rect 174538 189088 174544 189100
rect 122800 189060 174544 189088
rect 122800 189048 122806 189060
rect 174538 189048 174544 189060
rect 174596 189048 174602 189100
rect 224218 189048 224224 189100
rect 224276 189088 224282 189100
rect 243078 189088 243084 189100
rect 224276 189060 243084 189088
rect 224276 189048 224282 189060
rect 243078 189048 243084 189060
rect 243136 189048 243142 189100
rect 2774 188844 2780 188896
rect 2832 188884 2838 188896
rect 4798 188884 4804 188896
rect 2832 188856 4804 188884
rect 2832 188844 2838 188856
rect 4798 188844 4804 188856
rect 4856 188844 4862 188896
rect 188430 188368 188436 188420
rect 188488 188408 188494 188420
rect 204530 188408 204536 188420
rect 188488 188380 204536 188408
rect 188488 188368 188494 188380
rect 204530 188368 204536 188380
rect 204588 188368 204594 188420
rect 206370 188368 206376 188420
rect 206428 188408 206434 188420
rect 233418 188408 233424 188420
rect 206428 188380 233424 188408
rect 206428 188368 206434 188380
rect 233418 188368 233424 188380
rect 233476 188368 233482 188420
rect 32398 188300 32404 188352
rect 32456 188340 32462 188352
rect 159358 188340 159364 188352
rect 32456 188312 159364 188340
rect 32456 188300 32462 188312
rect 159358 188300 159364 188312
rect 159416 188300 159422 188352
rect 162762 188300 162768 188352
rect 162820 188340 162826 188352
rect 177574 188340 177580 188352
rect 162820 188312 177580 188340
rect 162820 188300 162826 188312
rect 177574 188300 177580 188312
rect 177632 188300 177638 188352
rect 201494 188300 201500 188352
rect 201552 188340 201558 188352
rect 249794 188340 249800 188352
rect 201552 188312 249800 188340
rect 201552 188300 201558 188312
rect 249794 188300 249800 188312
rect 249852 188300 249858 188352
rect 268378 188300 268384 188352
rect 268436 188340 268442 188352
rect 296898 188340 296904 188352
rect 268436 188312 296904 188340
rect 268436 188300 268442 188312
rect 296898 188300 296904 188312
rect 296956 188300 296962 188352
rect 300302 188300 300308 188352
rect 300360 188340 300366 188352
rect 310698 188340 310704 188352
rect 300360 188312 310704 188340
rect 300360 188300 300366 188312
rect 310698 188300 310704 188312
rect 310756 188300 310762 188352
rect 125502 187688 125508 187740
rect 125560 187728 125566 187740
rect 202138 187728 202144 187740
rect 125560 187700 202144 187728
rect 125560 187688 125566 187700
rect 202138 187688 202144 187700
rect 202196 187688 202202 187740
rect 282178 187144 282184 187196
rect 282236 187184 282242 187196
rect 284570 187184 284576 187196
rect 282236 187156 284576 187184
rect 282236 187144 282242 187156
rect 284570 187144 284576 187156
rect 284628 187144 284634 187196
rect 191742 186940 191748 186992
rect 191800 186980 191806 186992
rect 235350 186980 235356 186992
rect 191800 186952 235356 186980
rect 191800 186940 191806 186952
rect 235350 186940 235356 186952
rect 235408 186940 235414 186992
rect 126882 186396 126888 186448
rect 126940 186436 126946 186448
rect 164878 186436 164884 186448
rect 126940 186408 164884 186436
rect 126940 186396 126946 186408
rect 164878 186396 164884 186408
rect 164936 186396 164942 186448
rect 110322 186328 110328 186380
rect 110380 186368 110386 186380
rect 187142 186368 187148 186380
rect 110380 186340 187148 186368
rect 110380 186328 110386 186340
rect 187142 186328 187148 186340
rect 187200 186328 187206 186380
rect 204530 186260 204536 186312
rect 204588 186300 204594 186312
rect 224218 186300 224224 186312
rect 204588 186272 224224 186300
rect 204588 186260 204594 186272
rect 224218 186260 224224 186272
rect 224276 186260 224282 186312
rect 191098 185648 191104 185700
rect 191156 185688 191162 185700
rect 204990 185688 204996 185700
rect 191156 185660 204996 185688
rect 191156 185648 191162 185660
rect 204990 185648 204996 185660
rect 205048 185648 205054 185700
rect 215294 185648 215300 185700
rect 215352 185688 215358 185700
rect 227806 185688 227812 185700
rect 215352 185660 227812 185688
rect 215352 185648 215358 185660
rect 227806 185648 227812 185660
rect 227864 185648 227870 185700
rect 181530 185580 181536 185632
rect 181588 185620 181594 185632
rect 216030 185620 216036 185632
rect 181588 185592 216036 185620
rect 181588 185580 181594 185592
rect 216030 185580 216036 185592
rect 216088 185580 216094 185632
rect 226334 185580 226340 185632
rect 226392 185620 226398 185632
rect 249886 185620 249892 185632
rect 226392 185592 249892 185620
rect 226392 185580 226398 185592
rect 249886 185580 249892 185592
rect 249944 185580 249950 185632
rect 266998 185580 267004 185632
rect 267056 185620 267062 185632
rect 279142 185620 279148 185632
rect 267056 185592 279148 185620
rect 267056 185580 267062 185592
rect 279142 185580 279148 185592
rect 279200 185580 279206 185632
rect 130930 184968 130936 185020
rect 130988 185008 130994 185020
rect 169202 185008 169208 185020
rect 130988 184980 169208 185008
rect 130988 184968 130994 184980
rect 169202 184968 169208 184980
rect 169260 184968 169266 185020
rect 148870 184900 148876 184952
rect 148928 184940 148934 184952
rect 191098 184940 191104 184952
rect 148928 184912 191104 184940
rect 148928 184900 148934 184912
rect 191098 184900 191104 184912
rect 191156 184900 191162 184952
rect 272426 184900 272432 184952
rect 272484 184940 272490 184952
rect 302418 184940 302424 184952
rect 272484 184912 302424 184940
rect 272484 184900 272490 184912
rect 302418 184900 302424 184912
rect 302476 184900 302482 184952
rect 207014 184832 207020 184884
rect 207072 184872 207078 184884
rect 226334 184872 226340 184884
rect 207072 184844 226340 184872
rect 207072 184832 207078 184844
rect 226334 184832 226340 184844
rect 226392 184832 226398 184884
rect 271230 184832 271236 184884
rect 271288 184872 271294 184884
rect 279602 184872 279608 184884
rect 271288 184844 279608 184872
rect 271288 184832 271294 184844
rect 279602 184832 279608 184844
rect 279660 184832 279666 184884
rect 196618 184152 196624 184204
rect 196676 184192 196682 184204
rect 231118 184192 231124 184204
rect 196676 184164 231124 184192
rect 196676 184152 196682 184164
rect 231118 184152 231124 184164
rect 231176 184152 231182 184204
rect 257430 184152 257436 184204
rect 257488 184192 257494 184204
rect 280246 184192 280252 184204
rect 257488 184164 280252 184192
rect 257488 184152 257494 184164
rect 280246 184152 280252 184164
rect 280304 184152 280310 184204
rect 334802 184152 334808 184204
rect 334860 184192 334866 184204
rect 396902 184192 396908 184204
rect 334860 184164 396908 184192
rect 334860 184152 334866 184164
rect 396902 184152 396908 184164
rect 396960 184152 396966 184204
rect 133782 183608 133788 183660
rect 133840 183648 133846 183660
rect 162118 183648 162124 183660
rect 133840 183620 162124 183648
rect 133840 183608 133846 183620
rect 162118 183608 162124 183620
rect 162176 183608 162182 183660
rect 124858 183540 124864 183592
rect 124916 183580 124922 183592
rect 200758 183580 200764 183592
rect 124916 183552 200764 183580
rect 124916 183540 124922 183552
rect 200758 183540 200764 183552
rect 200816 183540 200822 183592
rect 224310 182860 224316 182912
rect 224368 182900 224374 182912
rect 232038 182900 232044 182912
rect 224368 182872 232044 182900
rect 224368 182860 224374 182872
rect 232038 182860 232044 182872
rect 232096 182860 232102 182912
rect 180702 182792 180708 182844
rect 180760 182832 180766 182844
rect 215110 182832 215116 182844
rect 180760 182804 215116 182832
rect 180760 182792 180766 182804
rect 215110 182792 215116 182804
rect 215168 182792 215174 182844
rect 215938 182792 215944 182844
rect 215996 182832 216002 182844
rect 241514 182832 241520 182844
rect 215996 182804 241520 182832
rect 215996 182792 216002 182804
rect 241514 182792 241520 182804
rect 241572 182792 241578 182844
rect 270310 182792 270316 182844
rect 270368 182832 270374 182844
rect 303798 182832 303804 182844
rect 270368 182804 303804 182832
rect 270368 182792 270374 182804
rect 303798 182792 303804 182804
rect 303856 182792 303862 182844
rect 114370 182248 114376 182300
rect 114428 182288 114434 182300
rect 164970 182288 164976 182300
rect 114428 182260 164976 182288
rect 114428 182248 114434 182260
rect 164970 182248 164976 182260
rect 165028 182248 165034 182300
rect 103330 182180 103336 182232
rect 103388 182220 103394 182232
rect 171870 182220 171876 182232
rect 103388 182192 171876 182220
rect 103388 182180 103394 182192
rect 171870 182180 171876 182192
rect 171928 182180 171934 182232
rect 211890 182112 211896 182164
rect 211948 182152 211954 182164
rect 272426 182152 272432 182164
rect 211948 182124 272432 182152
rect 211948 182112 211954 182124
rect 272426 182112 272432 182124
rect 272484 182112 272490 182164
rect 269850 181500 269856 181552
rect 269908 181540 269914 181552
rect 283098 181540 283104 181552
rect 269908 181512 283104 181540
rect 269908 181500 269914 181512
rect 283098 181500 283104 181512
rect 283156 181500 283162 181552
rect 273898 181432 273904 181484
rect 273956 181472 273962 181484
rect 294046 181472 294052 181484
rect 273956 181444 294052 181472
rect 273956 181432 273962 181444
rect 294046 181432 294052 181444
rect 294104 181432 294110 181484
rect 124030 180888 124036 180940
rect 124088 180928 124094 180940
rect 166534 180928 166540 180940
rect 124088 180900 166540 180928
rect 124088 180888 124094 180900
rect 166534 180888 166540 180900
rect 166592 180888 166598 180940
rect 132402 180820 132408 180872
rect 132460 180860 132466 180872
rect 211798 180860 211804 180872
rect 132460 180832 211804 180860
rect 132460 180820 132466 180832
rect 211798 180820 211804 180832
rect 211856 180820 211862 180872
rect 226978 180820 226984 180872
rect 227036 180860 227042 180872
rect 229278 180860 229284 180872
rect 227036 180832 229284 180860
rect 227036 180820 227042 180832
rect 229278 180820 229284 180832
rect 229336 180820 229342 180872
rect 204990 180752 204996 180804
rect 205048 180792 205054 180804
rect 218790 180792 218796 180804
rect 205048 180764 218796 180792
rect 205048 180752 205054 180764
rect 218790 180752 218796 180764
rect 218848 180752 218854 180804
rect 260098 180140 260104 180192
rect 260156 180180 260162 180192
rect 285858 180180 285864 180192
rect 260156 180152 285864 180180
rect 260156 180140 260162 180152
rect 285858 180140 285864 180152
rect 285916 180140 285922 180192
rect 220078 180072 220084 180124
rect 220136 180112 220142 180124
rect 234706 180112 234712 180124
rect 220136 180084 234712 180112
rect 220136 180072 220142 180084
rect 234706 180072 234712 180084
rect 234764 180072 234770 180124
rect 262858 180072 262864 180124
rect 262916 180112 262922 180124
rect 291378 180112 291384 180124
rect 262916 180084 291384 180112
rect 262916 180072 262922 180084
rect 291378 180072 291384 180084
rect 291436 180072 291442 180124
rect 119522 179460 119528 179512
rect 119580 179500 119586 179512
rect 198090 179500 198096 179512
rect 119580 179472 198096 179500
rect 119580 179460 119586 179472
rect 198090 179460 198096 179472
rect 198148 179460 198154 179512
rect 129458 179392 129464 179444
rect 129516 179432 129522 179444
rect 214190 179432 214196 179444
rect 129516 179404 214196 179432
rect 129516 179392 129522 179404
rect 214190 179392 214196 179404
rect 214248 179392 214254 179444
rect 215938 179392 215944 179444
rect 215996 179432 216002 179444
rect 230842 179432 230848 179444
rect 215996 179404 230848 179432
rect 215996 179392 216002 179404
rect 230842 179392 230848 179404
rect 230900 179392 230906 179444
rect 230382 179324 230388 179376
rect 230440 179364 230446 179376
rect 258074 179364 258080 179376
rect 230440 179336 258080 179364
rect 230440 179324 230446 179336
rect 258074 179324 258080 179336
rect 258132 179364 258138 179376
rect 259270 179364 259276 179376
rect 258132 179336 259276 179364
rect 258132 179324 258138 179336
rect 259270 179324 259276 179336
rect 259328 179324 259334 179376
rect 215110 178712 215116 178764
rect 215168 178752 215174 178764
rect 240318 178752 240324 178764
rect 215168 178724 240324 178752
rect 215168 178712 215174 178724
rect 240318 178712 240324 178724
rect 240376 178712 240382 178764
rect 271138 178712 271144 178764
rect 271196 178752 271202 178764
rect 283006 178752 283012 178764
rect 271196 178724 283012 178752
rect 271196 178712 271202 178724
rect 283006 178712 283012 178724
rect 283064 178712 283070 178764
rect 283558 178712 283564 178764
rect 283616 178752 283622 178764
rect 298186 178752 298192 178764
rect 283616 178724 298192 178752
rect 283616 178712 283622 178724
rect 298186 178712 298192 178724
rect 298244 178712 298250 178764
rect 177942 178644 177948 178696
rect 178000 178684 178006 178696
rect 229554 178684 229560 178696
rect 178000 178656 229560 178684
rect 178000 178644 178006 178656
rect 229554 178644 229560 178656
rect 229612 178644 229618 178696
rect 262122 178644 262128 178696
rect 262180 178684 262186 178696
rect 280338 178684 280344 178696
rect 262180 178656 280344 178684
rect 262180 178644 262186 178656
rect 280338 178644 280344 178656
rect 280396 178644 280402 178696
rect 280890 178644 280896 178696
rect 280948 178684 280954 178696
rect 299566 178684 299572 178696
rect 280948 178656 299572 178684
rect 280948 178644 280954 178656
rect 299566 178644 299572 178656
rect 299624 178644 299630 178696
rect 115842 178100 115848 178152
rect 115900 178140 115906 178152
rect 170582 178140 170588 178152
rect 115900 178112 170588 178140
rect 115900 178100 115906 178112
rect 170582 178100 170588 178112
rect 170640 178100 170646 178152
rect 113726 178032 113732 178084
rect 113784 178072 113790 178084
rect 177482 178072 177488 178084
rect 113784 178044 177488 178072
rect 113784 178032 113790 178044
rect 177482 178032 177488 178044
rect 177540 178032 177546 178084
rect 120810 177964 120816 178016
rect 120868 178004 120874 178016
rect 124858 178004 124864 178016
rect 120868 177976 124864 178004
rect 120868 177964 120874 177976
rect 124858 177964 124864 177976
rect 124916 177964 124922 178016
rect 275462 177964 275468 178016
rect 275520 178004 275526 178016
rect 284294 178004 284300 178016
rect 275520 177976 284300 178004
rect 275520 177964 275526 177976
rect 284294 177964 284300 177976
rect 284352 177964 284358 178016
rect 282270 177896 282276 177948
rect 282328 177936 282334 177948
rect 288710 177936 288716 177948
rect 282328 177908 288716 177936
rect 282328 177896 282334 177908
rect 288710 177896 288716 177908
rect 288768 177896 288774 177948
rect 226334 177556 226340 177608
rect 226392 177596 226398 177608
rect 230566 177596 230572 177608
rect 226392 177568 230572 177596
rect 226392 177556 226398 177568
rect 230566 177556 230572 177568
rect 230624 177556 230630 177608
rect 181622 177352 181628 177404
rect 181680 177392 181686 177404
rect 207658 177392 207664 177404
rect 181680 177364 207664 177392
rect 181680 177352 181686 177364
rect 207658 177352 207664 177364
rect 207716 177352 207722 177404
rect 284938 177352 284944 177404
rect 284996 177392 285002 177404
rect 289814 177392 289820 177404
rect 284996 177364 289820 177392
rect 284996 177352 285002 177364
rect 289814 177352 289820 177364
rect 289872 177352 289878 177404
rect 181438 177284 181444 177336
rect 181496 177324 181502 177336
rect 234614 177324 234620 177336
rect 181496 177296 234620 177324
rect 181496 177284 181502 177296
rect 234614 177284 234620 177296
rect 234672 177284 234678 177336
rect 235258 177284 235264 177336
rect 235316 177324 235322 177336
rect 243170 177324 243176 177336
rect 235316 177296 243176 177324
rect 235316 177284 235322 177296
rect 243170 177284 243176 177296
rect 243228 177284 243234 177336
rect 276750 177284 276756 177336
rect 276808 177324 276814 177336
rect 280798 177324 280804 177336
rect 276808 177296 280804 177324
rect 276808 177284 276814 177296
rect 280798 177284 280804 177296
rect 280856 177284 280862 177336
rect 298738 177284 298744 177336
rect 298796 177324 298802 177336
rect 371970 177324 371976 177336
rect 298796 177296 371976 177324
rect 298796 177284 298802 177296
rect 371970 177284 371976 177296
rect 372028 177284 372034 177336
rect 158990 176740 158996 176792
rect 159048 176780 159054 176792
rect 166258 176780 166264 176792
rect 159048 176752 166264 176780
rect 159048 176740 159054 176752
rect 166258 176740 166264 176752
rect 166316 176740 166322 176792
rect 127066 176672 127072 176724
rect 127124 176712 127130 176724
rect 165430 176712 165436 176724
rect 127124 176684 165436 176712
rect 127124 176672 127130 176684
rect 165430 176672 165436 176684
rect 165488 176672 165494 176724
rect 231118 176672 231124 176724
rect 231176 176712 231182 176724
rect 231854 176712 231860 176724
rect 231176 176684 231860 176712
rect 231176 176672 231182 176684
rect 231854 176672 231860 176684
rect 231912 176672 231918 176724
rect 135714 176604 135720 176656
rect 135772 176644 135778 176656
rect 213914 176644 213920 176656
rect 135772 176616 213920 176644
rect 135772 176604 135778 176616
rect 213914 176604 213920 176616
rect 213972 176604 213978 176656
rect 228358 175992 228364 176044
rect 228416 176032 228422 176044
rect 234798 176032 234804 176044
rect 228416 176004 234804 176032
rect 228416 175992 228422 176004
rect 234798 175992 234804 176004
rect 234856 175992 234862 176044
rect 134426 175924 134432 175976
rect 134484 175964 134490 175976
rect 165522 175964 165528 175976
rect 134484 175936 165528 175964
rect 134484 175924 134490 175936
rect 165522 175924 165528 175936
rect 165580 175924 165586 175976
rect 218698 175924 218704 175976
rect 218756 175964 218762 175976
rect 233234 175964 233240 175976
rect 218756 175936 233240 175964
rect 218756 175924 218762 175936
rect 233234 175924 233240 175936
rect 233292 175924 233298 175976
rect 239398 175924 239404 175976
rect 239456 175964 239462 175976
rect 281902 175964 281908 175976
rect 239456 175936 281908 175964
rect 239456 175924 239462 175936
rect 281902 175924 281908 175936
rect 281960 175924 281966 175976
rect 305178 175924 305184 175976
rect 305236 175964 305242 175976
rect 316126 175964 316132 175976
rect 305236 175936 316132 175964
rect 305236 175924 305242 175936
rect 316126 175924 316132 175936
rect 316184 175924 316190 175976
rect 333882 175924 333888 175976
rect 333940 175964 333946 175976
rect 401686 175964 401692 175976
rect 333940 175936 401692 175964
rect 333940 175924 333946 175936
rect 401686 175924 401692 175936
rect 401744 175924 401750 175976
rect 278222 175788 278228 175840
rect 278280 175828 278286 175840
rect 279326 175828 279332 175840
rect 278280 175800 279332 175828
rect 278280 175788 278286 175800
rect 279326 175788 279332 175800
rect 279384 175788 279390 175840
rect 215386 175244 215392 175296
rect 215444 175284 215450 175296
rect 229002 175284 229008 175296
rect 215444 175256 229008 175284
rect 215444 175244 215450 175256
rect 229002 175244 229008 175256
rect 229060 175244 229066 175296
rect 239490 175244 239496 175296
rect 239548 175284 239554 175296
rect 264974 175284 264980 175296
rect 239548 175256 264980 175284
rect 239548 175244 239554 175256
rect 264974 175244 264980 175256
rect 265032 175244 265038 175296
rect 281534 175244 281540 175296
rect 281592 175284 281598 175296
rect 305178 175284 305184 175296
rect 281592 175256 305184 175284
rect 281592 175244 281598 175256
rect 305178 175244 305184 175256
rect 305236 175284 305242 175296
rect 305638 175284 305644 175296
rect 305236 175256 305644 175284
rect 305236 175244 305242 175256
rect 305638 175244 305644 175256
rect 305696 175244 305702 175296
rect 162118 175176 162124 175228
rect 162176 175216 162182 175228
rect 214006 175216 214012 175228
rect 162176 175188 214012 175216
rect 162176 175176 162182 175188
rect 214006 175176 214012 175188
rect 214064 175176 214070 175228
rect 230474 175176 230480 175228
rect 230532 175216 230538 175228
rect 244918 175216 244924 175228
rect 230532 175188 244924 175216
rect 230532 175176 230538 175188
rect 244918 175176 244924 175188
rect 244976 175176 244982 175228
rect 281810 175176 281816 175228
rect 281868 175216 281874 175228
rect 305270 175216 305276 175228
rect 281868 175188 305276 175216
rect 281868 175176 281874 175188
rect 305270 175176 305276 175188
rect 305328 175176 305334 175228
rect 165522 175108 165528 175160
rect 165580 175148 165586 175160
rect 213914 175148 213920 175160
rect 165580 175120 213920 175148
rect 165580 175108 165586 175120
rect 213914 175108 213920 175120
rect 213972 175108 213978 175160
rect 229094 174564 229100 174616
rect 229152 174604 229158 174616
rect 229278 174604 229284 174616
rect 229152 174576 229284 174604
rect 229152 174564 229158 174576
rect 229278 174564 229284 174576
rect 229336 174564 229342 174616
rect 229002 173992 229008 174004
rect 219406 173964 229008 173992
rect 215294 173884 215300 173936
rect 215352 173924 215358 173936
rect 219406 173924 219434 173964
rect 229002 173952 229008 173964
rect 229060 173952 229066 174004
rect 230014 173952 230020 174004
rect 230072 173992 230078 174004
rect 230934 173992 230940 174004
rect 230072 173964 230940 173992
rect 230072 173952 230078 173964
rect 230934 173952 230940 173964
rect 230992 173952 230998 174004
rect 245010 173952 245016 174004
rect 245068 173992 245074 174004
rect 264974 173992 264980 174004
rect 245068 173964 264980 173992
rect 245068 173952 245074 173964
rect 264974 173952 264980 173964
rect 265032 173952 265038 174004
rect 215352 173896 219434 173924
rect 215352 173884 215358 173896
rect 238202 173884 238208 173936
rect 238260 173924 238266 173936
rect 265066 173924 265072 173936
rect 238260 173896 265072 173924
rect 238260 173884 238266 173896
rect 265066 173884 265072 173896
rect 265124 173884 265130 173936
rect 169202 173816 169208 173868
rect 169260 173856 169266 173868
rect 213914 173856 213920 173868
rect 169260 173828 213920 173856
rect 169260 173816 169266 173828
rect 213914 173816 213920 173828
rect 213972 173816 213978 173868
rect 211798 173748 211804 173800
rect 211856 173788 211862 173800
rect 214466 173788 214472 173800
rect 211856 173760 214472 173788
rect 211856 173748 211862 173760
rect 214466 173748 214472 173760
rect 214524 173748 214530 173800
rect 231670 173136 231676 173188
rect 231728 173176 231734 173188
rect 244458 173176 244464 173188
rect 231728 173148 244464 173176
rect 231728 173136 231734 173148
rect 244458 173136 244464 173148
rect 244516 173136 244522 173188
rect 300118 173136 300124 173188
rect 300176 173176 300182 173188
rect 419626 173176 419632 173188
rect 300176 173148 419632 173176
rect 300176 173136 300182 173148
rect 419626 173136 419632 173148
rect 419684 173136 419690 173188
rect 250530 172592 250536 172644
rect 250588 172632 250594 172644
rect 265066 172632 265072 172644
rect 250588 172604 265072 172632
rect 250588 172592 250594 172604
rect 265066 172592 265072 172604
rect 265124 172592 265130 172644
rect 236914 172524 236920 172576
rect 236972 172564 236978 172576
rect 264974 172564 264980 172576
rect 236972 172536 264980 172564
rect 236972 172524 236978 172536
rect 264974 172524 264980 172536
rect 265032 172524 265038 172576
rect 166350 172456 166356 172508
rect 166408 172496 166414 172508
rect 215294 172496 215300 172508
rect 166408 172468 215300 172496
rect 166408 172456 166414 172468
rect 215294 172456 215300 172468
rect 215352 172456 215358 172508
rect 231394 172456 231400 172508
rect 231452 172496 231458 172508
rect 248598 172496 248604 172508
rect 231452 172468 248604 172496
rect 231452 172456 231458 172468
rect 248598 172456 248604 172468
rect 248656 172456 248662 172508
rect 190362 172388 190368 172440
rect 190420 172428 190426 172440
rect 216766 172428 216772 172440
rect 190420 172400 216772 172428
rect 190420 172388 190426 172400
rect 216766 172388 216772 172400
rect 216824 172388 216830 172440
rect 231762 172388 231768 172440
rect 231820 172428 231826 172440
rect 242986 172428 242992 172440
rect 231820 172400 242992 172428
rect 231820 172388 231826 172400
rect 242986 172388 242992 172400
rect 243044 172388 243050 172440
rect 289814 171816 289820 171828
rect 282886 171788 289820 171816
rect 254578 171164 254584 171216
rect 254636 171204 254642 171216
rect 265066 171204 265072 171216
rect 254636 171176 265072 171204
rect 254636 171164 254642 171176
rect 265066 171164 265072 171176
rect 265124 171164 265130 171216
rect 249334 171096 249340 171148
rect 249392 171136 249398 171148
rect 264974 171136 264980 171148
rect 249392 171108 264980 171136
rect 249392 171096 249398 171108
rect 264974 171096 264980 171108
rect 265032 171096 265038 171148
rect 282886 171136 282914 171788
rect 289814 171776 289820 171788
rect 289872 171776 289878 171828
rect 354122 171776 354128 171828
rect 354180 171816 354186 171828
rect 417418 171816 417424 171828
rect 354180 171788 417424 171816
rect 354180 171776 354186 171788
rect 417418 171776 417424 171788
rect 417476 171776 417482 171828
rect 280080 171108 282914 171136
rect 164878 171028 164884 171080
rect 164936 171068 164942 171080
rect 213914 171068 213920 171080
rect 164936 171040 213920 171068
rect 164936 171028 164942 171040
rect 213914 171028 213920 171040
rect 213972 171028 213978 171080
rect 210510 170960 210516 171012
rect 210568 171000 210574 171012
rect 214006 171000 214012 171012
rect 210568 170972 214012 171000
rect 210568 170960 210574 170972
rect 214006 170960 214012 170972
rect 214064 170960 214070 171012
rect 280080 170944 280108 171108
rect 280062 170892 280068 170944
rect 280120 170892 280126 170944
rect 230750 170620 230756 170672
rect 230808 170660 230814 170672
rect 233234 170660 233240 170672
rect 230808 170632 233240 170660
rect 230808 170620 230814 170632
rect 233234 170620 233240 170632
rect 233292 170620 233298 170672
rect 231118 170348 231124 170400
rect 231176 170388 231182 170400
rect 247034 170388 247040 170400
rect 231176 170360 247040 170388
rect 231176 170348 231182 170360
rect 247034 170348 247040 170360
rect 247092 170348 247098 170400
rect 342990 170348 342996 170400
rect 343048 170388 343054 170400
rect 392762 170388 392768 170400
rect 343048 170360 392768 170388
rect 343048 170348 343054 170360
rect 392762 170348 392768 170360
rect 392820 170348 392826 170400
rect 247678 169804 247684 169856
rect 247736 169844 247742 169856
rect 264974 169844 264980 169856
rect 247736 169816 264980 169844
rect 247736 169804 247742 169816
rect 264974 169804 264980 169816
rect 265032 169804 265038 169856
rect 240870 169736 240876 169788
rect 240928 169776 240934 169788
rect 265066 169776 265072 169788
rect 240928 169748 265072 169776
rect 240928 169736 240934 169748
rect 265066 169736 265072 169748
rect 265124 169736 265130 169788
rect 166534 169668 166540 169720
rect 166592 169708 166598 169720
rect 214006 169708 214012 169720
rect 166592 169680 214012 169708
rect 166592 169668 166598 169680
rect 214006 169668 214012 169680
rect 214064 169668 214070 169720
rect 281534 169668 281540 169720
rect 281592 169708 281598 169720
rect 284662 169708 284668 169720
rect 281592 169680 284668 169708
rect 281592 169668 281598 169680
rect 284662 169668 284668 169680
rect 284720 169668 284726 169720
rect 202138 169600 202144 169652
rect 202196 169640 202202 169652
rect 213914 169640 213920 169652
rect 202196 169612 213920 169640
rect 202196 169600 202202 169612
rect 213914 169600 213920 169612
rect 213972 169600 213978 169652
rect 231762 169532 231768 169584
rect 231820 169572 231826 169584
rect 235994 169572 236000 169584
rect 231820 169544 236000 169572
rect 231820 169532 231826 169544
rect 235994 169532 236000 169544
rect 236052 169532 236058 169584
rect 231762 169124 231768 169176
rect 231820 169164 231826 169176
rect 234706 169164 234712 169176
rect 231820 169136 234712 169164
rect 231820 169124 231826 169136
rect 234706 169124 234712 169136
rect 234764 169124 234770 169176
rect 242250 168444 242256 168496
rect 242308 168484 242314 168496
rect 264974 168484 264980 168496
rect 242308 168456 264980 168484
rect 242308 168444 242314 168456
rect 264974 168444 264980 168456
rect 265032 168444 265038 168496
rect 235258 168376 235264 168428
rect 235316 168416 235322 168428
rect 265066 168416 265072 168428
rect 235316 168388 265072 168416
rect 235316 168376 235322 168388
rect 265066 168376 265072 168388
rect 265124 168376 265130 168428
rect 174538 168308 174544 168360
rect 174596 168348 174602 168360
rect 213914 168348 213920 168360
rect 174596 168320 213920 168348
rect 174596 168308 174602 168320
rect 213914 168308 213920 168320
rect 213972 168308 213978 168360
rect 231486 168308 231492 168360
rect 231544 168348 231550 168360
rect 234798 168348 234804 168360
rect 231544 168320 234804 168348
rect 231544 168308 231550 168320
rect 234798 168308 234804 168320
rect 234856 168308 234862 168360
rect 200758 168240 200764 168292
rect 200816 168280 200822 168292
rect 214006 168280 214012 168292
rect 200816 168252 214012 168280
rect 200816 168240 200822 168252
rect 214006 168240 214012 168252
rect 214064 168240 214070 168292
rect 234706 167968 234712 168020
rect 234764 168008 234770 168020
rect 237374 168008 237380 168020
rect 234764 167980 237380 168008
rect 234764 167968 234770 167980
rect 237374 167968 237380 167980
rect 237432 167968 237438 168020
rect 308398 167628 308404 167680
rect 308456 167668 308462 167680
rect 434714 167668 434720 167680
rect 308456 167640 434720 167668
rect 308456 167628 308462 167640
rect 434714 167628 434720 167640
rect 434772 167628 434778 167680
rect 262950 167084 262956 167136
rect 263008 167124 263014 167136
rect 265342 167124 265348 167136
rect 263008 167096 265348 167124
rect 263008 167084 263014 167096
rect 265342 167084 265348 167096
rect 265400 167084 265406 167136
rect 233970 167016 233976 167068
rect 234028 167056 234034 167068
rect 264974 167056 264980 167068
rect 234028 167028 264980 167056
rect 234028 167016 234034 167028
rect 264974 167016 264980 167028
rect 265032 167016 265038 167068
rect 170490 166948 170496 167000
rect 170548 166988 170554 167000
rect 214006 166988 214012 167000
rect 170548 166960 214012 166988
rect 170548 166948 170554 166960
rect 214006 166948 214012 166960
rect 214064 166948 214070 167000
rect 281902 166948 281908 167000
rect 281960 166988 281966 167000
rect 291470 166988 291476 167000
rect 281960 166960 291476 166988
rect 281960 166948 281966 166960
rect 291470 166948 291476 166960
rect 291528 166948 291534 167000
rect 198090 166880 198096 166932
rect 198148 166920 198154 166932
rect 213914 166920 213920 166932
rect 198148 166892 213920 166920
rect 198148 166880 198154 166892
rect 213914 166880 213920 166892
rect 213972 166880 213978 166932
rect 231302 166880 231308 166932
rect 231360 166920 231366 166932
rect 234614 166920 234620 166932
rect 231360 166892 234620 166920
rect 231360 166880 231366 166892
rect 234614 166880 234620 166892
rect 234672 166880 234678 166932
rect 231762 166676 231768 166728
rect 231820 166716 231826 166728
rect 234706 166716 234712 166728
rect 231820 166688 234712 166716
rect 231820 166676 231826 166688
rect 234706 166676 234712 166688
rect 234764 166676 234770 166728
rect 249058 165656 249064 165708
rect 249116 165696 249122 165708
rect 265066 165696 265072 165708
rect 249116 165668 265072 165696
rect 249116 165656 249122 165668
rect 265066 165656 265072 165668
rect 265124 165656 265130 165708
rect 237006 165588 237012 165640
rect 237064 165628 237070 165640
rect 264974 165628 264980 165640
rect 237064 165600 264980 165628
rect 237064 165588 237070 165600
rect 264974 165588 264980 165600
rect 265032 165588 265038 165640
rect 170582 165520 170588 165572
rect 170640 165560 170646 165572
rect 213914 165560 213920 165572
rect 170640 165532 213920 165560
rect 170640 165520 170646 165532
rect 213914 165520 213920 165532
rect 213972 165520 213978 165572
rect 231486 165180 231492 165232
rect 231544 165220 231550 165232
rect 234614 165220 234620 165232
rect 231544 165192 234620 165220
rect 231544 165180 231550 165192
rect 234614 165180 234620 165192
rect 234672 165180 234678 165232
rect 230934 165112 230940 165164
rect 230992 165152 230998 165164
rect 233326 165152 233332 165164
rect 230992 165124 233332 165152
rect 230992 165112 230998 165124
rect 233326 165112 233332 165124
rect 233384 165112 233390 165164
rect 282178 164908 282184 164960
rect 282236 164948 282242 164960
rect 310698 164948 310704 164960
rect 282236 164920 310704 164948
rect 282236 164908 282242 164920
rect 310698 164908 310704 164920
rect 310756 164908 310762 164960
rect 300210 164840 300216 164892
rect 300268 164880 300274 164892
rect 381722 164880 381728 164892
rect 300268 164852 381728 164880
rect 300268 164840 300274 164852
rect 381722 164840 381728 164852
rect 381780 164840 381786 164892
rect 257338 164296 257344 164348
rect 257396 164336 257402 164348
rect 264974 164336 264980 164348
rect 257396 164308 264980 164336
rect 257396 164296 257402 164308
rect 264974 164296 264980 164308
rect 265032 164296 265038 164348
rect 247770 164228 247776 164280
rect 247828 164268 247834 164280
rect 265066 164268 265072 164280
rect 247828 164240 265072 164268
rect 247828 164228 247834 164240
rect 265066 164228 265072 164240
rect 265124 164228 265130 164280
rect 282822 164228 282828 164280
rect 282880 164268 282886 164280
rect 287238 164268 287244 164280
rect 282880 164240 287244 164268
rect 282880 164228 282886 164240
rect 287238 164228 287244 164240
rect 287296 164228 287302 164280
rect 3326 164160 3332 164212
rect 3384 164200 3390 164212
rect 29638 164200 29644 164212
rect 3384 164172 29644 164200
rect 3384 164160 3390 164172
rect 29638 164160 29644 164172
rect 29696 164160 29702 164212
rect 176102 164160 176108 164212
rect 176160 164200 176166 164212
rect 214006 164200 214012 164212
rect 176160 164172 214012 164200
rect 176160 164160 176166 164172
rect 214006 164160 214012 164172
rect 214064 164160 214070 164212
rect 231026 164160 231032 164212
rect 231084 164200 231090 164212
rect 248414 164200 248420 164212
rect 231084 164172 248420 164200
rect 231084 164160 231090 164172
rect 248414 164160 248420 164172
rect 248472 164160 248478 164212
rect 177482 164092 177488 164144
rect 177540 164132 177546 164144
rect 213914 164132 213920 164144
rect 177540 164104 213920 164132
rect 177540 164092 177546 164104
rect 213914 164092 213920 164104
rect 213972 164092 213978 164144
rect 167822 163480 167828 163532
rect 167880 163520 167886 163532
rect 175918 163520 175924 163532
rect 167880 163492 175924 163520
rect 167880 163480 167886 163492
rect 175918 163480 175924 163492
rect 175976 163480 175982 163532
rect 245102 163480 245108 163532
rect 245160 163520 245166 163532
rect 265434 163520 265440 163532
rect 245160 163492 265440 163520
rect 245160 163480 245166 163492
rect 265434 163480 265440 163492
rect 265492 163480 265498 163532
rect 281810 163480 281816 163532
rect 281868 163520 281874 163532
rect 295334 163520 295340 163532
rect 281868 163492 295340 163520
rect 281868 163480 281874 163492
rect 295334 163480 295340 163492
rect 295392 163480 295398 163532
rect 341610 163480 341616 163532
rect 341668 163520 341674 163532
rect 444558 163520 444564 163532
rect 341668 163492 444564 163520
rect 341668 163480 341674 163492
rect 444558 163480 444564 163492
rect 444616 163480 444622 163532
rect 282822 163072 282828 163124
rect 282880 163112 282886 163124
rect 288710 163112 288716 163124
rect 282880 163084 288716 163112
rect 282880 163072 282886 163084
rect 288710 163072 288716 163084
rect 288768 163072 288774 163124
rect 252186 162868 252192 162920
rect 252244 162908 252250 162920
rect 265066 162908 265072 162920
rect 252244 162880 265072 162908
rect 252244 162868 252250 162880
rect 265066 162868 265072 162880
rect 265124 162868 265130 162920
rect 166442 162800 166448 162852
rect 166500 162840 166506 162852
rect 213914 162840 213920 162852
rect 166500 162812 213920 162840
rect 166500 162800 166506 162812
rect 213914 162800 213920 162812
rect 213972 162800 213978 162852
rect 242434 162800 242440 162852
rect 242492 162840 242498 162852
rect 243078 162840 243084 162852
rect 242492 162812 243084 162840
rect 242492 162800 242498 162812
rect 243078 162800 243084 162812
rect 243136 162800 243142 162852
rect 243538 162800 243544 162852
rect 243596 162840 243602 162852
rect 244366 162840 244372 162852
rect 243596 162812 244372 162840
rect 243596 162800 243602 162812
rect 244366 162800 244372 162812
rect 244424 162800 244430 162852
rect 281626 162800 281632 162852
rect 281684 162840 281690 162852
rect 303890 162840 303896 162852
rect 281684 162812 303896 162840
rect 281684 162800 281690 162812
rect 303890 162800 303896 162812
rect 303948 162800 303954 162852
rect 187142 162732 187148 162784
rect 187200 162772 187206 162784
rect 214006 162772 214012 162784
rect 187200 162744 214012 162772
rect 187200 162732 187206 162744
rect 214006 162732 214012 162744
rect 214064 162732 214070 162784
rect 231670 162732 231676 162784
rect 231728 162772 231734 162784
rect 241606 162772 241612 162784
rect 231728 162744 241612 162772
rect 231728 162732 231734 162744
rect 241606 162732 241612 162744
rect 241664 162732 241670 162784
rect 256142 162120 256148 162172
rect 256200 162160 256206 162172
rect 264974 162160 264980 162172
rect 256200 162132 264980 162160
rect 256200 162120 256206 162132
rect 264974 162120 264980 162132
rect 265032 162120 265038 162172
rect 281902 161780 281908 161832
rect 281960 161820 281966 161832
rect 286318 161820 286324 161832
rect 281960 161792 286324 161820
rect 281960 161780 281966 161792
rect 286318 161780 286324 161792
rect 286376 161780 286382 161832
rect 235534 161440 235540 161492
rect 235592 161480 235598 161492
rect 265066 161480 265072 161492
rect 235592 161452 265072 161480
rect 235592 161440 235598 161452
rect 265066 161440 265072 161452
rect 265124 161440 265130 161492
rect 165522 161372 165528 161424
rect 165580 161412 165586 161424
rect 214006 161412 214012 161424
rect 165580 161384 214012 161412
rect 165580 161372 165586 161384
rect 214006 161372 214012 161384
rect 214064 161372 214070 161424
rect 282822 161372 282828 161424
rect 282880 161412 282886 161424
rect 317506 161412 317512 161424
rect 282880 161384 317512 161412
rect 282880 161372 282886 161384
rect 317506 161372 317512 161384
rect 317564 161372 317570 161424
rect 173342 161304 173348 161356
rect 173400 161344 173406 161356
rect 213914 161344 213920 161356
rect 173400 161316 213920 161344
rect 173400 161304 173406 161316
rect 213914 161304 213920 161316
rect 213972 161304 213978 161356
rect 231026 161032 231032 161084
rect 231084 161072 231090 161084
rect 233510 161072 233516 161084
rect 231084 161044 233516 161072
rect 231084 161032 231090 161044
rect 233510 161032 233516 161044
rect 233568 161032 233574 161084
rect 249702 160692 249708 160744
rect 249760 160732 249766 160744
rect 262950 160732 262956 160744
rect 249760 160704 262956 160732
rect 249760 160692 249766 160704
rect 262950 160692 262956 160704
rect 263008 160692 263014 160744
rect 356790 160692 356796 160744
rect 356848 160732 356854 160744
rect 395430 160732 395436 160744
rect 356848 160704 395436 160732
rect 356848 160692 356854 160704
rect 395430 160692 395436 160704
rect 395488 160692 395494 160744
rect 282822 160420 282828 160472
rect 282880 160460 282886 160472
rect 287330 160460 287336 160472
rect 282880 160432 287336 160460
rect 282880 160420 282886 160432
rect 287330 160420 287336 160432
rect 287388 160420 287394 160472
rect 263042 160148 263048 160200
rect 263100 160188 263106 160200
rect 265434 160188 265440 160200
rect 263100 160160 265440 160188
rect 263100 160148 263106 160160
rect 265434 160148 265440 160160
rect 265492 160148 265498 160200
rect 229738 160080 229744 160132
rect 229796 160120 229802 160132
rect 231946 160120 231952 160132
rect 229796 160092 231952 160120
rect 229796 160080 229802 160092
rect 231946 160080 231952 160092
rect 232004 160080 232010 160132
rect 245194 160080 245200 160132
rect 245252 160120 245258 160132
rect 264974 160120 264980 160132
rect 245252 160092 264980 160120
rect 245252 160080 245258 160092
rect 264974 160080 264980 160092
rect 265032 160080 265038 160132
rect 167638 160012 167644 160064
rect 167696 160052 167702 160064
rect 213914 160052 213920 160064
rect 167696 160024 213920 160052
rect 167696 160012 167702 160024
rect 213914 160012 213920 160024
rect 213972 160012 213978 160064
rect 282822 160012 282828 160064
rect 282880 160052 282886 160064
rect 293954 160052 293960 160064
rect 282880 160024 293960 160052
rect 282880 160012 282886 160024
rect 293954 160012 293960 160024
rect 294012 160012 294018 160064
rect 230566 159400 230572 159452
rect 230624 159440 230630 159452
rect 240226 159440 240232 159452
rect 230624 159412 240232 159440
rect 230624 159400 230630 159412
rect 240226 159400 240232 159412
rect 240284 159400 240290 159452
rect 232682 159332 232688 159384
rect 232740 159372 232746 159384
rect 265250 159372 265256 159384
rect 232740 159344 265256 159372
rect 232740 159332 232746 159344
rect 265250 159332 265256 159344
rect 265308 159332 265314 159384
rect 307110 159332 307116 159384
rect 307168 159372 307174 159384
rect 409966 159372 409972 159384
rect 307168 159344 409972 159372
rect 307168 159332 307174 159344
rect 409966 159332 409972 159344
rect 410024 159332 410030 159384
rect 241054 158720 241060 158772
rect 241112 158760 241118 158772
rect 264974 158760 264980 158772
rect 241112 158732 264980 158760
rect 241112 158720 241118 158732
rect 264974 158720 264980 158732
rect 265032 158720 265038 158772
rect 171870 158652 171876 158704
rect 171928 158692 171934 158704
rect 213914 158692 213920 158704
rect 171928 158664 213920 158692
rect 171928 158652 171934 158664
rect 213914 158652 213920 158664
rect 213972 158652 213978 158704
rect 231762 158652 231768 158704
rect 231820 158692 231826 158704
rect 241698 158692 241704 158704
rect 231820 158664 241704 158692
rect 231820 158652 231826 158664
rect 241698 158652 241704 158664
rect 241756 158652 241762 158704
rect 282086 158652 282092 158704
rect 282144 158692 282150 158704
rect 292758 158692 292764 158704
rect 282144 158664 292764 158692
rect 282144 158652 282150 158664
rect 292758 158652 292764 158664
rect 292816 158652 292822 158704
rect 180242 158584 180248 158636
rect 180300 158624 180306 158636
rect 214006 158624 214012 158636
rect 180300 158596 214012 158624
rect 180300 158584 180306 158596
rect 214006 158584 214012 158596
rect 214064 158584 214070 158636
rect 231486 158584 231492 158636
rect 231544 158624 231550 158636
rect 234246 158624 234252 158636
rect 231544 158596 234252 158624
rect 231544 158584 231550 158596
rect 234246 158584 234252 158596
rect 234304 158584 234310 158636
rect 322290 157972 322296 158024
rect 322348 158012 322354 158024
rect 430574 158012 430580 158024
rect 322348 157984 430580 158012
rect 322348 157972 322354 157984
rect 430574 157972 430580 157984
rect 430632 157972 430638 158024
rect 242158 157428 242164 157480
rect 242216 157468 242222 157480
rect 264974 157468 264980 157480
rect 242216 157440 264980 157468
rect 242216 157428 242222 157440
rect 264974 157428 264980 157440
rect 265032 157428 265038 157480
rect 238294 157360 238300 157412
rect 238352 157400 238358 157412
rect 265066 157400 265072 157412
rect 238352 157372 265072 157400
rect 238352 157360 238358 157372
rect 265066 157360 265072 157372
rect 265124 157360 265130 157412
rect 281534 157360 281540 157412
rect 281592 157400 281598 157412
rect 283190 157400 283196 157412
rect 281592 157372 283196 157400
rect 281592 157360 281598 157372
rect 283190 157360 283196 157372
rect 283248 157360 283254 157412
rect 169110 157292 169116 157344
rect 169168 157332 169174 157344
rect 213914 157332 213920 157344
rect 169168 157304 213920 157332
rect 169168 157292 169174 157304
rect 213914 157292 213920 157304
rect 213972 157292 213978 157344
rect 231762 157292 231768 157344
rect 231820 157332 231826 157344
rect 244274 157332 244280 157344
rect 231820 157304 244280 157332
rect 231820 157292 231826 157304
rect 244274 157292 244280 157304
rect 244332 157292 244338 157344
rect 180150 157224 180156 157276
rect 180208 157264 180214 157276
rect 214006 157264 214012 157276
rect 180208 157236 214012 157264
rect 180208 157224 180214 157236
rect 214006 157224 214012 157236
rect 214064 157224 214070 157276
rect 318058 156612 318064 156664
rect 318116 156652 318122 156664
rect 422294 156652 422300 156664
rect 318116 156624 422300 156652
rect 318116 156612 318122 156624
rect 422294 156612 422300 156624
rect 422352 156612 422358 156664
rect 250622 156000 250628 156052
rect 250680 156040 250686 156052
rect 265066 156040 265072 156052
rect 250680 156012 265072 156040
rect 250680 156000 250686 156012
rect 265066 156000 265072 156012
rect 265124 156000 265130 156052
rect 246298 155932 246304 155984
rect 246356 155972 246362 155984
rect 264974 155972 264980 155984
rect 246356 155944 264980 155972
rect 246356 155932 246362 155944
rect 264974 155932 264980 155944
rect 265032 155932 265038 155984
rect 170398 155864 170404 155916
rect 170456 155904 170462 155916
rect 214006 155904 214012 155916
rect 170456 155876 214012 155904
rect 170456 155864 170462 155876
rect 214006 155864 214012 155876
rect 214064 155864 214070 155916
rect 231762 155864 231768 155916
rect 231820 155904 231826 155916
rect 238754 155904 238760 155916
rect 231820 155876 238760 155904
rect 231820 155864 231826 155876
rect 238754 155864 238760 155876
rect 238812 155864 238818 155916
rect 282270 155864 282276 155916
rect 282328 155904 282334 155916
rect 311986 155904 311992 155916
rect 282328 155876 311992 155904
rect 282328 155864 282334 155876
rect 311986 155864 311992 155876
rect 312044 155864 312050 155916
rect 178862 155796 178868 155848
rect 178920 155836 178926 155848
rect 213914 155836 213920 155848
rect 178920 155808 213920 155836
rect 178920 155796 178926 155808
rect 213914 155796 213920 155808
rect 213972 155796 213978 155848
rect 239674 155184 239680 155236
rect 239732 155224 239738 155236
rect 249702 155224 249708 155236
rect 239732 155196 249708 155224
rect 239732 155184 239738 155196
rect 249702 155184 249708 155196
rect 249760 155184 249766 155236
rect 358078 155184 358084 155236
rect 358136 155224 358142 155236
rect 436830 155224 436836 155236
rect 358136 155196 436836 155224
rect 358136 155184 358142 155196
rect 436830 155184 436836 155196
rect 436888 155184 436894 155236
rect 250438 154640 250444 154692
rect 250496 154680 250502 154692
rect 264974 154680 264980 154692
rect 250496 154652 264980 154680
rect 250496 154640 250502 154652
rect 264974 154640 264980 154652
rect 265032 154640 265038 154692
rect 233878 154572 233884 154624
rect 233936 154612 233942 154624
rect 265066 154612 265072 154624
rect 233936 154584 265072 154612
rect 233936 154572 233942 154584
rect 265066 154572 265072 154584
rect 265124 154572 265130 154624
rect 282822 154504 282828 154556
rect 282880 154544 282886 154556
rect 306466 154544 306472 154556
rect 282880 154516 306472 154544
rect 282880 154504 282886 154516
rect 306466 154504 306472 154516
rect 306524 154504 306530 154556
rect 282086 154436 282092 154488
rect 282144 154476 282150 154488
rect 302234 154476 302240 154488
rect 282144 154448 302240 154476
rect 282144 154436 282150 154448
rect 302234 154436 302240 154448
rect 302292 154436 302298 154488
rect 230658 153824 230664 153876
rect 230716 153864 230722 153876
rect 245838 153864 245844 153876
rect 230716 153836 245844 153864
rect 230716 153824 230722 153836
rect 245838 153824 245844 153836
rect 245896 153824 245902 153876
rect 309778 153824 309784 153876
rect 309836 153864 309842 153876
rect 423030 153864 423036 153876
rect 309836 153836 423036 153864
rect 309836 153824 309842 153836
rect 423030 153824 423036 153836
rect 423088 153824 423094 153876
rect 231210 153688 231216 153740
rect 231268 153728 231274 153740
rect 233418 153728 233424 153740
rect 231268 153700 233424 153728
rect 231268 153688 231274 153700
rect 233418 153688 233424 153700
rect 233476 153688 233482 153740
rect 211890 153280 211896 153332
rect 211948 153320 211954 153332
rect 214006 153320 214012 153332
rect 211948 153292 214012 153320
rect 211948 153280 211954 153292
rect 214006 153280 214012 153292
rect 214064 153280 214070 153332
rect 195422 153212 195428 153264
rect 195480 153252 195486 153264
rect 213914 153252 213920 153264
rect 195480 153224 213920 153252
rect 195480 153212 195486 153224
rect 213914 153212 213920 153224
rect 213972 153212 213978 153264
rect 253198 153212 253204 153264
rect 253256 153252 253262 153264
rect 264974 153252 264980 153264
rect 253256 153224 264980 153252
rect 253256 153212 253262 153224
rect 264974 153212 264980 153224
rect 265032 153212 265038 153264
rect 230474 152464 230480 152516
rect 230532 152504 230538 152516
rect 238846 152504 238852 152516
rect 230532 152476 238852 152504
rect 230532 152464 230538 152476
rect 238846 152464 238852 152476
rect 238904 152464 238910 152516
rect 319438 152464 319444 152516
rect 319496 152504 319502 152516
rect 441798 152504 441804 152516
rect 319496 152476 441804 152504
rect 319496 152464 319502 152476
rect 441798 152464 441804 152476
rect 441856 152464 441862 152516
rect 211982 152056 211988 152108
rect 212040 152096 212046 152108
rect 214006 152096 214012 152108
rect 212040 152068 214012 152096
rect 212040 152056 212046 152068
rect 214006 152056 214012 152068
rect 214064 152056 214070 152108
rect 249242 151852 249248 151904
rect 249300 151892 249306 151904
rect 265066 151892 265072 151904
rect 249300 151864 265072 151892
rect 249300 151852 249306 151864
rect 265066 151852 265072 151864
rect 265124 151852 265130 151904
rect 202230 151784 202236 151836
rect 202288 151824 202294 151836
rect 213914 151824 213920 151836
rect 202288 151796 213920 151824
rect 202288 151784 202294 151796
rect 213914 151784 213920 151796
rect 213972 151784 213978 151836
rect 238110 151784 238116 151836
rect 238168 151824 238174 151836
rect 264974 151824 264980 151836
rect 238168 151796 264980 151824
rect 238168 151784 238174 151796
rect 264974 151784 264980 151796
rect 265032 151784 265038 151836
rect 281902 151716 281908 151768
rect 281960 151756 281966 151768
rect 300854 151756 300860 151768
rect 281960 151728 300860 151756
rect 281960 151716 281966 151728
rect 300854 151716 300860 151728
rect 300912 151716 300918 151768
rect 230474 151580 230480 151632
rect 230532 151620 230538 151632
rect 232130 151620 232136 151632
rect 230532 151592 232136 151620
rect 230532 151580 230538 151592
rect 232130 151580 232136 151592
rect 232188 151580 232194 151632
rect 238386 151104 238392 151156
rect 238444 151144 238450 151156
rect 263042 151144 263048 151156
rect 238444 151116 263048 151144
rect 238444 151104 238450 151116
rect 263042 151104 263048 151116
rect 263100 151104 263106 151156
rect 374730 151104 374736 151156
rect 374788 151144 374794 151156
rect 429930 151144 429936 151156
rect 374788 151116 429936 151144
rect 374788 151104 374794 151116
rect 429930 151104 429936 151116
rect 429988 151104 429994 151156
rect 436738 151104 436744 151156
rect 436796 151144 436802 151156
rect 448606 151144 448612 151156
rect 436796 151116 448612 151144
rect 436796 151104 436802 151116
rect 448606 151104 448612 151116
rect 448664 151104 448670 151156
rect 229922 151036 229928 151088
rect 229980 151076 229986 151088
rect 265710 151076 265716 151088
rect 229980 151048 265716 151076
rect 229980 151036 229986 151048
rect 265710 151036 265716 151048
rect 265768 151036 265774 151088
rect 282270 151036 282276 151088
rect 282328 151076 282334 151088
rect 289906 151076 289912 151088
rect 282328 151048 289912 151076
rect 282328 151036 282334 151048
rect 289906 151036 289912 151048
rect 289964 151036 289970 151088
rect 398742 151036 398748 151088
rect 398800 151076 398806 151088
rect 583018 151076 583024 151088
rect 398800 151048 583024 151076
rect 398800 151036 398806 151048
rect 583018 151036 583024 151048
rect 583076 151036 583082 151088
rect 198090 150492 198096 150544
rect 198148 150532 198154 150544
rect 214006 150532 214012 150544
rect 198148 150504 214012 150532
rect 198148 150492 198154 150504
rect 214006 150492 214012 150504
rect 214064 150492 214070 150544
rect 180334 150424 180340 150476
rect 180392 150464 180398 150476
rect 213914 150464 213920 150476
rect 180392 150436 213920 150464
rect 180392 150424 180398 150436
rect 213914 150424 213920 150436
rect 213972 150424 213978 150476
rect 262950 150424 262956 150476
rect 263008 150464 263014 150476
rect 265342 150464 265348 150476
rect 263008 150436 265348 150464
rect 263008 150424 263014 150436
rect 265342 150424 265348 150436
rect 265400 150424 265406 150476
rect 3602 150356 3608 150408
rect 3660 150396 3666 150408
rect 11698 150396 11704 150408
rect 3660 150368 11704 150396
rect 3660 150356 3666 150368
rect 11698 150356 11704 150368
rect 11756 150356 11762 150408
rect 175918 150356 175924 150408
rect 175976 150396 175982 150408
rect 214006 150396 214012 150408
rect 175976 150368 214012 150396
rect 175976 150356 175982 150368
rect 214006 150356 214012 150368
rect 214064 150356 214070 150408
rect 282730 150356 282736 150408
rect 282788 150396 282794 150408
rect 307846 150396 307852 150408
rect 282788 150368 307852 150396
rect 282788 150356 282794 150368
rect 307846 150356 307852 150368
rect 307904 150356 307910 150408
rect 191098 150288 191104 150340
rect 191156 150328 191162 150340
rect 213914 150328 213920 150340
rect 191156 150300 213920 150328
rect 191156 150288 191162 150300
rect 213914 150288 213920 150300
rect 213972 150288 213978 150340
rect 282822 150288 282828 150340
rect 282880 150328 282886 150340
rect 302418 150328 302424 150340
rect 282880 150300 302424 150328
rect 282880 150288 282886 150300
rect 302418 150288 302424 150300
rect 302476 150288 302482 150340
rect 239398 149676 239404 149728
rect 239456 149716 239462 149728
rect 265618 149716 265624 149728
rect 239456 149688 265624 149716
rect 239456 149676 239462 149688
rect 265618 149676 265624 149688
rect 265676 149676 265682 149728
rect 367738 149676 367744 149728
rect 367796 149716 367802 149728
rect 439590 149716 439596 149728
rect 367796 149688 439596 149716
rect 367796 149676 367802 149688
rect 439590 149676 439596 149688
rect 439648 149676 439654 149728
rect 235442 149064 235448 149116
rect 235500 149104 235506 149116
rect 264974 149104 264980 149116
rect 235500 149076 264980 149104
rect 235500 149064 235506 149076
rect 264974 149064 264980 149076
rect 265032 149064 265038 149116
rect 166258 148996 166264 149048
rect 166316 149036 166322 149048
rect 213914 149036 213920 149048
rect 166316 149008 213920 149036
rect 166316 148996 166322 149008
rect 213914 148996 213920 149008
rect 213972 148996 213978 149048
rect 282822 148996 282828 149048
rect 282880 149036 282886 149048
rect 310606 149036 310612 149048
rect 282880 149008 310612 149036
rect 282880 148996 282886 149008
rect 310606 148996 310612 149008
rect 310664 148996 310670 149048
rect 449894 148996 449900 149048
rect 449952 149036 449958 149048
rect 582834 149036 582840 149048
rect 449952 149008 582840 149036
rect 449952 148996 449958 149008
rect 582834 148996 582840 149008
rect 582892 148996 582898 149048
rect 282178 148928 282184 148980
rect 282236 148968 282242 148980
rect 288526 148968 288532 148980
rect 282236 148940 288532 148968
rect 282236 148928 282242 148940
rect 288526 148928 288532 148940
rect 288584 148928 288590 148980
rect 429838 148384 429844 148436
rect 429896 148424 429902 148436
rect 440418 148424 440424 148436
rect 429896 148396 440424 148424
rect 429896 148384 429902 148396
rect 440418 148384 440424 148396
rect 440476 148384 440482 148436
rect 231118 148316 231124 148368
rect 231176 148356 231182 148368
rect 240870 148356 240876 148368
rect 231176 148328 240876 148356
rect 231176 148316 231182 148328
rect 240870 148316 240876 148328
rect 240928 148316 240934 148368
rect 437658 148316 437664 148368
rect 437716 148356 437722 148368
rect 449894 148356 449900 148368
rect 437716 148328 449900 148356
rect 437716 148316 437722 148328
rect 449894 148316 449900 148328
rect 449952 148316 449958 148368
rect 240962 147704 240968 147756
rect 241020 147744 241026 147756
rect 264974 147744 264980 147756
rect 241020 147716 264980 147744
rect 241020 147704 241026 147716
rect 264974 147704 264980 147716
rect 265032 147704 265038 147756
rect 209222 147636 209228 147688
rect 209280 147676 209286 147688
rect 213914 147676 213920 147688
rect 209280 147648 213920 147676
rect 209280 147636 209286 147648
rect 213914 147636 213920 147648
rect 213972 147636 213978 147688
rect 234062 147636 234068 147688
rect 234120 147676 234126 147688
rect 265066 147676 265072 147688
rect 234120 147648 265072 147676
rect 234120 147636 234126 147648
rect 265066 147636 265072 147648
rect 265124 147636 265130 147688
rect 281718 147568 281724 147620
rect 281776 147608 281782 147620
rect 299566 147608 299572 147620
rect 281776 147580 299572 147608
rect 281776 147568 281782 147580
rect 299566 147568 299572 147580
rect 299624 147568 299630 147620
rect 282822 147500 282828 147552
rect 282880 147540 282886 147552
rect 291378 147540 291384 147552
rect 282880 147512 291384 147540
rect 282880 147500 282886 147512
rect 291378 147500 291384 147512
rect 291436 147500 291442 147552
rect 432690 146956 432696 147008
rect 432748 146996 432754 147008
rect 443270 146996 443276 147008
rect 432748 146968 443276 146996
rect 432748 146956 432754 146968
rect 443270 146956 443276 146968
rect 443328 146956 443334 147008
rect 580902 146956 580908 147008
rect 580960 146996 580966 147008
rect 582742 146996 582748 147008
rect 580960 146968 582748 146996
rect 580960 146956 580966 146968
rect 582742 146956 582748 146968
rect 582800 146956 582806 147008
rect 169018 146888 169024 146940
rect 169076 146928 169082 146940
rect 204990 146928 204996 146940
rect 169076 146900 204996 146928
rect 169076 146888 169082 146900
rect 204990 146888 204996 146900
rect 205048 146888 205054 146940
rect 231854 146888 231860 146940
rect 231912 146928 231918 146940
rect 248506 146928 248512 146940
rect 231912 146900 248512 146928
rect 231912 146888 231918 146900
rect 248506 146888 248512 146900
rect 248564 146888 248570 146940
rect 298830 146888 298836 146940
rect 298888 146928 298894 146940
rect 404722 146928 404728 146940
rect 298888 146900 404728 146928
rect 298888 146888 298894 146900
rect 404722 146888 404728 146900
rect 404780 146888 404786 146940
rect 414658 146888 414664 146940
rect 414716 146928 414722 146940
rect 436370 146928 436376 146940
rect 414716 146900 436376 146928
rect 414716 146888 414722 146900
rect 436370 146888 436376 146900
rect 436428 146888 436434 146940
rect 441798 146820 441804 146872
rect 441856 146860 441862 146872
rect 441982 146860 441988 146872
rect 441856 146832 441988 146860
rect 441856 146820 441862 146832
rect 441982 146820 441988 146832
rect 442040 146820 442046 146872
rect 263042 146344 263048 146396
rect 263100 146384 263106 146396
rect 265158 146384 265164 146396
rect 263100 146356 265164 146384
rect 263100 146344 263106 146356
rect 265158 146344 265164 146356
rect 265216 146344 265222 146396
rect 169110 146276 169116 146328
rect 169168 146316 169174 146328
rect 213914 146316 213920 146328
rect 169168 146288 213920 146316
rect 169168 146276 169174 146288
rect 213914 146276 213920 146288
rect 213972 146276 213978 146328
rect 240870 146276 240876 146328
rect 240928 146316 240934 146328
rect 265066 146316 265072 146328
rect 240928 146288 265072 146316
rect 240928 146276 240934 146288
rect 265066 146276 265072 146288
rect 265124 146276 265130 146328
rect 282822 146208 282828 146260
rect 282880 146248 282886 146260
rect 302326 146248 302332 146260
rect 282880 146220 302332 146248
rect 282880 146208 282886 146220
rect 302326 146208 302332 146220
rect 302384 146208 302390 146260
rect 403618 146208 403624 146260
rect 403676 146248 403682 146260
rect 411898 146248 411904 146260
rect 403676 146220 411904 146248
rect 403676 146208 403682 146220
rect 411898 146208 411904 146220
rect 411956 146208 411962 146260
rect 412542 146208 412548 146260
rect 412600 146248 412606 146260
rect 414474 146248 414480 146260
rect 412600 146220 414480 146248
rect 412600 146208 412606 146220
rect 414474 146208 414480 146220
rect 414532 146208 414538 146260
rect 392578 145528 392584 145580
rect 392636 145568 392642 145580
rect 407298 145568 407304 145580
rect 392636 145540 407304 145568
rect 392636 145528 392642 145540
rect 407298 145528 407304 145540
rect 407356 145528 407362 145580
rect 421466 145528 421472 145580
rect 421524 145568 421530 145580
rect 582558 145568 582564 145580
rect 421524 145540 582564 145568
rect 421524 145528 421530 145540
rect 582558 145528 582564 145540
rect 582616 145528 582622 145580
rect 235350 144984 235356 145036
rect 235408 145024 235414 145036
rect 264974 145024 264980 145036
rect 235408 144996 264980 145024
rect 235408 144984 235414 144996
rect 264974 144984 264980 144996
rect 265032 144984 265038 145036
rect 185670 144916 185676 144968
rect 185728 144956 185734 144968
rect 213914 144956 213920 144968
rect 185728 144928 213920 144956
rect 185728 144916 185734 144928
rect 213914 144916 213920 144928
rect 213972 144916 213978 144968
rect 232866 144916 232872 144968
rect 232924 144956 232930 144968
rect 265066 144956 265072 144968
rect 232924 144928 265072 144956
rect 232924 144916 232930 144928
rect 265066 144916 265072 144928
rect 265124 144916 265130 144968
rect 295978 144916 295984 144968
rect 296036 144956 296042 144968
rect 403434 144956 403440 144968
rect 296036 144928 403440 144956
rect 296036 144916 296042 144928
rect 403434 144916 403440 144928
rect 403492 144916 403498 144968
rect 231762 144848 231768 144900
rect 231820 144888 231826 144900
rect 240778 144888 240784 144900
rect 231820 144860 240784 144888
rect 231820 144848 231826 144860
rect 240778 144848 240784 144860
rect 240836 144848 240842 144900
rect 282822 144848 282828 144900
rect 282880 144888 282886 144900
rect 294046 144888 294052 144900
rect 282880 144860 294052 144888
rect 282880 144848 282886 144860
rect 294046 144848 294052 144860
rect 294104 144848 294110 144900
rect 417418 144848 417424 144900
rect 417476 144888 417482 144900
rect 418062 144888 418068 144900
rect 417476 144860 418068 144888
rect 417476 144848 417482 144860
rect 418062 144848 418068 144860
rect 418120 144888 418126 144900
rect 583294 144888 583300 144900
rect 418120 144860 583300 144888
rect 418120 144848 418126 144860
rect 583294 144848 583300 144860
rect 583352 144848 583358 144900
rect 170398 144168 170404 144220
rect 170456 144208 170462 144220
rect 214006 144208 214012 144220
rect 170456 144180 214012 144208
rect 170456 144168 170462 144180
rect 214006 144168 214012 144180
rect 214064 144168 214070 144220
rect 247862 144168 247868 144220
rect 247920 144208 247926 144220
rect 265158 144208 265164 144220
rect 247920 144180 265164 144208
rect 247920 144168 247926 144180
rect 265158 144168 265164 144180
rect 265216 144168 265222 144220
rect 280890 144168 280896 144220
rect 280948 144208 280954 144220
rect 296806 144208 296812 144220
rect 280948 144180 296812 144208
rect 280948 144168 280954 144180
rect 296806 144168 296812 144180
rect 296864 144168 296870 144220
rect 338758 144168 338764 144220
rect 338816 144208 338822 144220
rect 441706 144208 441712 144220
rect 338816 144180 441712 144208
rect 338816 144168 338822 144180
rect 441706 144168 441712 144180
rect 441764 144168 441770 144220
rect 171870 143556 171876 143608
rect 171928 143596 171934 143608
rect 213914 143596 213920 143608
rect 171928 143568 213920 143596
rect 171928 143556 171934 143568
rect 213914 143556 213920 143568
rect 213972 143556 213978 143608
rect 249150 143556 249156 143608
rect 249208 143596 249214 143608
rect 264974 143596 264980 143608
rect 249208 143568 264980 143596
rect 249208 143556 249214 143568
rect 264974 143556 264980 143568
rect 265032 143556 265038 143608
rect 300854 143488 300860 143540
rect 300912 143528 300918 143540
rect 301498 143528 301504 143540
rect 300912 143500 301504 143528
rect 300912 143488 300918 143500
rect 301498 143488 301504 143500
rect 301556 143488 301562 143540
rect 404998 143488 405004 143540
rect 405056 143528 405062 143540
rect 409046 143528 409052 143540
rect 405056 143500 409052 143528
rect 405056 143488 405062 143500
rect 409046 143488 409052 143500
rect 409104 143488 409110 143540
rect 418890 143488 418896 143540
rect 418948 143528 418954 143540
rect 419994 143528 420000 143540
rect 418948 143500 420000 143528
rect 418948 143488 418954 143500
rect 419994 143488 420000 143500
rect 420052 143488 420058 143540
rect 436830 143488 436836 143540
rect 436888 143528 436894 143540
rect 439314 143528 439320 143540
rect 436888 143500 439320 143528
rect 436888 143488 436894 143500
rect 439314 143488 439320 143500
rect 439372 143488 439378 143540
rect 231762 142808 231768 142860
rect 231820 142848 231826 142860
rect 241514 142848 241520 142860
rect 231820 142820 241520 142848
rect 231820 142808 231826 142820
rect 241514 142808 241520 142820
rect 241572 142808 241578 142860
rect 244274 142808 244280 142860
rect 244332 142848 244338 142860
rect 264974 142848 264980 142860
rect 244332 142820 264980 142848
rect 244332 142808 244338 142820
rect 264974 142808 264980 142820
rect 265032 142808 265038 142860
rect 422938 142808 422944 142860
rect 422996 142848 423002 142860
rect 432230 142848 432236 142860
rect 422996 142820 432236 142848
rect 422996 142808 423002 142820
rect 432230 142808 432236 142820
rect 432288 142808 432294 142860
rect 191098 142196 191104 142248
rect 191156 142236 191162 142248
rect 214006 142236 214012 142248
rect 191156 142208 214012 142236
rect 191156 142196 191162 142208
rect 214006 142196 214012 142208
rect 214064 142196 214070 142248
rect 396718 142196 396724 142248
rect 396776 142236 396782 142248
rect 414198 142236 414204 142248
rect 396776 142208 414204 142236
rect 396776 142196 396782 142208
rect 414198 142196 414204 142208
rect 414256 142196 414262 142248
rect 173250 142128 173256 142180
rect 173308 142168 173314 142180
rect 213914 142168 213920 142180
rect 173308 142140 213920 142168
rect 173308 142128 173314 142140
rect 213914 142128 213920 142140
rect 213972 142128 213978 142180
rect 257614 142128 257620 142180
rect 257672 142168 257678 142180
rect 265066 142168 265072 142180
rect 257672 142140 265072 142168
rect 257672 142128 257678 142140
rect 265066 142128 265072 142140
rect 265124 142128 265130 142180
rect 300854 142128 300860 142180
rect 300912 142168 300918 142180
rect 402606 142168 402612 142180
rect 300912 142140 402612 142168
rect 300912 142128 300918 142140
rect 402606 142128 402612 142140
rect 402664 142128 402670 142180
rect 428458 142128 428464 142180
rect 428516 142168 428522 142180
rect 432874 142168 432880 142180
rect 428516 142140 432880 142168
rect 428516 142128 428522 142140
rect 432874 142128 432880 142140
rect 432932 142168 432938 142180
rect 583018 142168 583024 142180
rect 432932 142140 583024 142168
rect 432932 142128 432938 142140
rect 583018 142128 583024 142140
rect 583076 142128 583082 142180
rect 282822 142060 282828 142112
rect 282880 142100 282886 142112
rect 295518 142100 295524 142112
rect 282880 142072 295524 142100
rect 282880 142060 282886 142072
rect 295518 142060 295524 142072
rect 295576 142060 295582 142112
rect 281902 141720 281908 141772
rect 281960 141760 281966 141772
rect 285858 141760 285864 141772
rect 281960 141732 285864 141760
rect 281960 141720 281966 141732
rect 285858 141720 285864 141732
rect 285916 141720 285922 141772
rect 247954 141448 247960 141500
rect 248012 141488 248018 141500
rect 265802 141488 265808 141500
rect 248012 141460 265808 141488
rect 248012 141448 248018 141460
rect 265802 141448 265808 141460
rect 265860 141448 265866 141500
rect 173158 141380 173164 141432
rect 173216 141420 173222 141432
rect 184290 141420 184296 141432
rect 173216 141392 184296 141420
rect 173216 141380 173222 141392
rect 184290 141380 184296 141392
rect 184348 141380 184354 141432
rect 232590 141380 232596 141432
rect 232648 141420 232654 141432
rect 265158 141420 265164 141432
rect 232648 141392 265164 141420
rect 232648 141380 232654 141392
rect 265158 141380 265164 141392
rect 265216 141380 265222 141432
rect 319438 141380 319444 141432
rect 319496 141420 319502 141432
rect 416774 141420 416780 141432
rect 319496 141392 416780 141420
rect 319496 141380 319502 141392
rect 416774 141380 416780 141392
rect 416832 141380 416838 141432
rect 431218 141380 431224 141432
rect 431276 141420 431282 141432
rect 440326 141420 440332 141432
rect 431276 141392 440332 141420
rect 431276 141380 431282 141392
rect 440326 141380 440332 141392
rect 440384 141380 440390 141432
rect 198182 140836 198188 140888
rect 198240 140876 198246 140888
rect 213914 140876 213920 140888
rect 198240 140848 213920 140876
rect 198240 140836 198246 140848
rect 213914 140836 213920 140848
rect 213972 140836 213978 140888
rect 317414 140836 317420 140888
rect 317472 140876 317478 140888
rect 317472 140848 412634 140876
rect 317472 140836 317478 140848
rect 191282 140768 191288 140820
rect 191340 140808 191346 140820
rect 214006 140808 214012 140820
rect 191340 140780 214012 140808
rect 191340 140768 191346 140780
rect 214006 140768 214012 140780
rect 214064 140768 214070 140820
rect 412606 140808 412634 140848
rect 422570 140836 422576 140888
rect 422628 140876 422634 140888
rect 423030 140876 423036 140888
rect 422628 140848 423036 140876
rect 422628 140836 422634 140848
rect 423030 140836 423036 140848
rect 423088 140876 423094 140888
rect 423088 140848 431954 140876
rect 423088 140836 423094 140848
rect 423674 140808 423680 140820
rect 412606 140780 423680 140808
rect 423674 140768 423680 140780
rect 423732 140808 423738 140820
rect 424502 140808 424508 140820
rect 423732 140780 424508 140808
rect 423732 140768 423738 140780
rect 424502 140768 424508 140780
rect 424560 140768 424566 140820
rect 431926 140808 431954 140848
rect 580258 140808 580264 140820
rect 431926 140780 580264 140808
rect 580258 140768 580264 140780
rect 580316 140768 580322 140820
rect 282730 140700 282736 140752
rect 282788 140740 282794 140752
rect 318794 140740 318800 140752
rect 282788 140712 318800 140740
rect 282788 140700 282794 140712
rect 318794 140700 318800 140712
rect 318852 140700 318858 140752
rect 400214 140700 400220 140752
rect 400272 140740 400278 140752
rect 400950 140740 400956 140752
rect 400272 140712 400956 140740
rect 400272 140700 400278 140712
rect 400950 140700 400956 140712
rect 401008 140700 401014 140752
rect 434714 140700 434720 140752
rect 434772 140740 434778 140752
rect 435174 140740 435180 140752
rect 434772 140712 435180 140740
rect 434772 140700 434778 140712
rect 435174 140700 435180 140712
rect 435232 140700 435238 140752
rect 436094 140700 436100 140752
rect 436152 140740 436158 140752
rect 437014 140740 437020 140752
rect 436152 140712 437020 140740
rect 436152 140700 436158 140712
rect 437014 140700 437020 140712
rect 437072 140700 437078 140752
rect 192478 140020 192484 140072
rect 192536 140060 192542 140072
rect 214190 140060 214196 140072
rect 192536 140032 214196 140060
rect 192536 140020 192542 140032
rect 214190 140020 214196 140032
rect 214248 140020 214254 140072
rect 307110 140020 307116 140072
rect 307168 140060 307174 140072
rect 317690 140060 317696 140072
rect 307168 140032 317696 140060
rect 307168 140020 307174 140032
rect 317690 140020 317696 140032
rect 317748 140060 317754 140072
rect 318702 140060 318708 140072
rect 317748 140032 318708 140060
rect 317748 140020 317754 140032
rect 318702 140020 318708 140032
rect 318760 140020 318766 140072
rect 420270 140020 420276 140072
rect 420328 140060 420334 140072
rect 440234 140060 440240 140072
rect 420328 140032 440240 140060
rect 420328 140020 420334 140032
rect 440234 140020 440240 140032
rect 440292 140020 440298 140072
rect 282822 139544 282828 139596
rect 282880 139584 282886 139596
rect 288434 139584 288440 139596
rect 282880 139556 288440 139584
rect 282880 139544 282886 139556
rect 288434 139544 288440 139556
rect 288492 139544 288498 139596
rect 399846 139544 399852 139596
rect 399904 139584 399910 139596
rect 400398 139584 400404 139596
rect 399904 139556 400404 139584
rect 399904 139544 399910 139556
rect 400398 139544 400404 139556
rect 400456 139544 400462 139596
rect 231210 139476 231216 139528
rect 231268 139516 231274 139528
rect 236914 139516 236920 139528
rect 231268 139488 236920 139516
rect 231268 139476 231274 139488
rect 236914 139476 236920 139488
rect 236972 139476 236978 139528
rect 398006 139476 398012 139528
rect 398064 139516 398070 139528
rect 404354 139516 404360 139528
rect 398064 139488 404360 139516
rect 398064 139476 398070 139488
rect 404354 139476 404360 139488
rect 404412 139476 404418 139528
rect 174538 139408 174544 139460
rect 174596 139448 174602 139460
rect 213914 139448 213920 139460
rect 174596 139420 213920 139448
rect 174596 139408 174602 139420
rect 213914 139408 213920 139420
rect 213972 139408 213978 139460
rect 231394 139408 231400 139460
rect 231452 139448 231458 139460
rect 235258 139448 235264 139460
rect 231452 139420 235264 139448
rect 231452 139408 231458 139420
rect 235258 139408 235264 139420
rect 235316 139408 235322 139460
rect 248046 139408 248052 139460
rect 248104 139448 248110 139460
rect 264974 139448 264980 139460
rect 248104 139420 264980 139448
rect 248104 139408 248110 139420
rect 264974 139408 264980 139420
rect 265032 139408 265038 139460
rect 318702 139408 318708 139460
rect 318760 139448 318766 139460
rect 417142 139448 417148 139460
rect 318760 139420 417148 139448
rect 318760 139408 318766 139420
rect 417142 139408 417148 139420
rect 417200 139408 417206 139460
rect 426802 139408 426808 139460
rect 426860 139448 426866 139460
rect 582650 139448 582656 139460
rect 426860 139420 582656 139448
rect 426860 139408 426866 139420
rect 582650 139408 582656 139420
rect 582708 139408 582714 139460
rect 231762 139340 231768 139392
rect 231820 139380 231826 139392
rect 255406 139380 255412 139392
rect 231820 139352 255412 139380
rect 231820 139340 231826 139352
rect 255406 139340 255412 139352
rect 255464 139340 255470 139392
rect 282822 139340 282828 139392
rect 282880 139380 282886 139392
rect 296898 139380 296904 139392
rect 282880 139352 296904 139380
rect 282880 139340 282886 139352
rect 296898 139340 296904 139352
rect 296956 139340 296962 139392
rect 398098 139340 398104 139392
rect 398156 139380 398162 139392
rect 412726 139380 412732 139392
rect 398156 139352 412732 139380
rect 398156 139340 398162 139352
rect 412726 139340 412732 139352
rect 412784 139340 412790 139392
rect 438210 139340 438216 139392
rect 438268 139380 438274 139392
rect 439498 139380 439504 139392
rect 438268 139352 439504 139380
rect 438268 139340 438274 139352
rect 439498 139340 439504 139352
rect 439556 139340 439562 139392
rect 231302 138796 231308 138848
rect 231360 138836 231366 138848
rect 238202 138836 238208 138848
rect 231360 138808 238208 138836
rect 231360 138796 231366 138808
rect 238202 138796 238208 138808
rect 238260 138796 238266 138848
rect 178770 138660 178776 138712
rect 178828 138700 178834 138712
rect 200758 138700 200764 138712
rect 178828 138672 200764 138700
rect 178828 138660 178834 138672
rect 200758 138660 200764 138672
rect 200816 138660 200822 138712
rect 263134 138048 263140 138100
rect 263192 138088 263198 138100
rect 265066 138088 265072 138100
rect 263192 138060 265072 138088
rect 263192 138048 263198 138060
rect 265066 138048 265072 138060
rect 265124 138048 265130 138100
rect 322290 138048 322296 138100
rect 322348 138088 322354 138100
rect 398098 138088 398104 138100
rect 322348 138060 398104 138088
rect 322348 138048 322354 138060
rect 398098 138048 398104 138060
rect 398156 138048 398162 138100
rect 175918 137980 175924 138032
rect 175976 138020 175982 138032
rect 213914 138020 213920 138032
rect 175976 137992 213920 138020
rect 175976 137980 175982 137992
rect 213914 137980 213920 137992
rect 213972 137980 213978 138032
rect 238018 137980 238024 138032
rect 238076 138020 238082 138032
rect 264974 138020 264980 138032
rect 238076 137992 264980 138020
rect 238076 137980 238082 137992
rect 264974 137980 264980 137992
rect 265032 137980 265038 138032
rect 398650 137980 398656 138032
rect 398708 138020 398714 138032
rect 580166 138020 580172 138032
rect 398708 137992 580172 138020
rect 398708 137980 398714 137992
rect 580166 137980 580172 137992
rect 580224 137980 580230 138032
rect 3326 137912 3332 137964
rect 3384 137952 3390 137964
rect 21358 137952 21364 137964
rect 3384 137924 21364 137952
rect 3384 137912 3390 137924
rect 21358 137912 21364 137924
rect 21416 137912 21422 137964
rect 231578 137912 231584 137964
rect 231636 137952 231642 137964
rect 249794 137952 249800 137964
rect 231636 137924 249800 137952
rect 231636 137912 231642 137924
rect 249794 137912 249800 137924
rect 249852 137912 249858 137964
rect 281626 137912 281632 137964
rect 281684 137952 281690 137964
rect 300946 137952 300952 137964
rect 281684 137924 300952 137952
rect 281684 137912 281690 137924
rect 300946 137912 300952 137924
rect 301004 137912 301010 137964
rect 327718 137912 327724 137964
rect 327776 137952 327782 137964
rect 397546 137952 397552 137964
rect 327776 137924 397552 137952
rect 327776 137912 327782 137924
rect 397546 137912 397552 137924
rect 397604 137912 397610 137964
rect 170674 137232 170680 137284
rect 170732 137272 170738 137284
rect 214374 137272 214380 137284
rect 170732 137244 214380 137272
rect 170732 137232 170738 137244
rect 214374 137232 214380 137244
rect 214432 137232 214438 137284
rect 264514 137232 264520 137284
rect 264572 137272 264578 137284
rect 265618 137272 265624 137284
rect 264572 137244 265624 137272
rect 264572 137232 264578 137244
rect 265618 137232 265624 137244
rect 265676 137232 265682 137284
rect 442902 136688 442908 136740
rect 442960 136728 442966 136740
rect 452746 136728 452752 136740
rect 442960 136700 452752 136728
rect 442960 136688 442966 136700
rect 452746 136688 452752 136700
rect 452804 136688 452810 136740
rect 229738 136620 229744 136672
rect 229796 136660 229802 136672
rect 264974 136660 264980 136672
rect 229796 136632 264980 136660
rect 229796 136620 229802 136632
rect 264974 136620 264980 136632
rect 265032 136620 265038 136672
rect 388438 136620 388444 136672
rect 388496 136660 388502 136672
rect 397546 136660 397552 136672
rect 388496 136632 397552 136660
rect 388496 136620 388502 136632
rect 397546 136620 397552 136632
rect 397604 136620 397610 136672
rect 440418 136620 440424 136672
rect 440476 136660 440482 136672
rect 582558 136660 582564 136672
rect 440476 136632 582564 136660
rect 440476 136620 440482 136632
rect 582558 136620 582564 136632
rect 582616 136620 582622 136672
rect 231486 136552 231492 136604
rect 231544 136592 231550 136604
rect 245010 136592 245016 136604
rect 231544 136564 245016 136592
rect 231544 136552 231550 136564
rect 245010 136552 245016 136564
rect 245068 136552 245074 136604
rect 395430 136552 395436 136604
rect 395488 136592 395494 136604
rect 397638 136592 397644 136604
rect 395488 136564 397644 136592
rect 395488 136552 395494 136564
rect 397638 136552 397644 136564
rect 397696 136552 397702 136604
rect 441982 136552 441988 136604
rect 442040 136592 442046 136604
rect 583386 136592 583392 136604
rect 442040 136564 583392 136592
rect 442040 136552 442046 136564
rect 583386 136552 583392 136564
rect 583444 136552 583450 136604
rect 231762 136484 231768 136536
rect 231820 136524 231826 136536
rect 242986 136524 242992 136536
rect 231820 136496 242992 136524
rect 231820 136484 231826 136496
rect 242986 136484 242992 136496
rect 243044 136484 243050 136536
rect 282270 136008 282276 136060
rect 282328 136048 282334 136060
rect 285674 136048 285680 136060
rect 282328 136020 285680 136048
rect 282328 136008 282334 136020
rect 285674 136008 285680 136020
rect 285732 136008 285738 136060
rect 328362 135872 328368 135924
rect 328420 135912 328426 135924
rect 398006 135912 398012 135924
rect 328420 135884 398012 135912
rect 328420 135872 328426 135884
rect 398006 135872 398012 135884
rect 398064 135872 398070 135924
rect 182910 135328 182916 135380
rect 182968 135368 182974 135380
rect 213914 135368 213920 135380
rect 182968 135340 213920 135368
rect 182968 135328 182974 135340
rect 213914 135328 213920 135340
rect 213972 135328 213978 135380
rect 250806 135328 250812 135380
rect 250864 135368 250870 135380
rect 265066 135368 265072 135380
rect 250864 135340 265072 135368
rect 250864 135328 250870 135340
rect 265066 135328 265072 135340
rect 265124 135328 265130 135380
rect 177482 135260 177488 135312
rect 177540 135300 177546 135312
rect 214006 135300 214012 135312
rect 177540 135272 214012 135300
rect 177540 135260 177546 135272
rect 214006 135260 214012 135272
rect 214064 135260 214070 135312
rect 243538 135260 243544 135312
rect 243596 135300 243602 135312
rect 264974 135300 264980 135312
rect 243596 135272 264980 135300
rect 243596 135260 243602 135272
rect 264974 135260 264980 135272
rect 265032 135260 265038 135312
rect 231486 135192 231492 135244
rect 231544 135232 231550 135244
rect 250530 135232 250536 135244
rect 231544 135204 250536 135232
rect 231544 135192 231550 135204
rect 250530 135192 250536 135204
rect 250588 135192 250594 135244
rect 363598 135192 363604 135244
rect 363656 135232 363662 135244
rect 398650 135232 398656 135244
rect 363656 135204 398656 135232
rect 363656 135192 363662 135204
rect 398650 135192 398656 135204
rect 398708 135192 398714 135244
rect 230750 135056 230756 135108
rect 230808 135096 230814 135108
rect 237006 135096 237012 135108
rect 230808 135068 237012 135096
rect 230808 135056 230814 135068
rect 237006 135056 237012 135068
rect 237064 135056 237070 135108
rect 178678 134580 178684 134632
rect 178736 134620 178742 134632
rect 199470 134620 199476 134632
rect 178736 134592 199476 134620
rect 178736 134580 178742 134592
rect 199470 134580 199476 134592
rect 199528 134580 199534 134632
rect 185578 134512 185584 134564
rect 185636 134552 185642 134564
rect 214098 134552 214104 134564
rect 185636 134524 214104 134552
rect 185636 134512 185642 134524
rect 214098 134512 214104 134524
rect 214156 134512 214162 134564
rect 250714 134512 250720 134564
rect 250772 134552 250778 134564
rect 265250 134552 265256 134564
rect 250772 134524 265256 134552
rect 250772 134512 250778 134524
rect 265250 134512 265256 134524
rect 265308 134512 265314 134564
rect 442902 134512 442908 134564
rect 442960 134552 442966 134564
rect 443086 134552 443092 134564
rect 442960 134524 443092 134552
rect 442960 134512 442966 134524
rect 443086 134512 443092 134524
rect 443144 134552 443150 134564
rect 456886 134552 456892 134564
rect 443144 134524 456892 134552
rect 443144 134512 443150 134524
rect 456886 134512 456892 134524
rect 456944 134512 456950 134564
rect 202138 133900 202144 133952
rect 202196 133940 202202 133952
rect 213914 133940 213920 133952
rect 202196 133912 213920 133940
rect 202196 133900 202202 133912
rect 213914 133900 213920 133912
rect 213972 133900 213978 133952
rect 260190 133900 260196 133952
rect 260248 133940 260254 133952
rect 264974 133940 264980 133952
rect 260248 133912 264980 133940
rect 260248 133900 260254 133912
rect 264974 133900 264980 133912
rect 265032 133900 265038 133952
rect 376110 133900 376116 133952
rect 376168 133940 376174 133952
rect 397546 133940 397552 133952
rect 376168 133912 397552 133940
rect 376168 133900 376174 133912
rect 397546 133900 397552 133912
rect 397604 133900 397610 133952
rect 231670 133832 231676 133884
rect 231728 133872 231734 133884
rect 254578 133872 254584 133884
rect 231728 133844 254584 133872
rect 231728 133832 231734 133844
rect 254578 133832 254584 133844
rect 254636 133832 254642 133884
rect 282822 133832 282828 133884
rect 282880 133872 282886 133884
rect 313366 133872 313372 133884
rect 282880 133844 313372 133872
rect 282880 133832 282886 133844
rect 313366 133832 313372 133844
rect 313424 133832 313430 133884
rect 342898 133832 342904 133884
rect 342956 133872 342962 133884
rect 397638 133872 397644 133884
rect 342956 133844 397644 133872
rect 342956 133832 342962 133844
rect 397638 133832 397644 133844
rect 397696 133832 397702 133884
rect 442902 133832 442908 133884
rect 442960 133872 442966 133884
rect 582466 133872 582472 133884
rect 442960 133844 582472 133872
rect 442960 133832 442966 133844
rect 582466 133832 582472 133844
rect 582524 133832 582530 133884
rect 231762 133764 231768 133816
rect 231820 133804 231826 133816
rect 253290 133804 253296 133816
rect 231820 133776 253296 133804
rect 231820 133764 231826 133776
rect 253290 133764 253296 133776
rect 253348 133764 253354 133816
rect 171778 133152 171784 133204
rect 171836 133192 171842 133204
rect 206462 133192 206468 133204
rect 171836 133164 206468 133192
rect 171836 133152 171842 133164
rect 206462 133152 206468 133164
rect 206520 133152 206526 133204
rect 211798 132540 211804 132592
rect 211856 132580 211862 132592
rect 214466 132580 214472 132592
rect 211856 132552 214472 132580
rect 211856 132540 211862 132552
rect 214466 132540 214472 132552
rect 214524 132540 214530 132592
rect 196802 132472 196808 132524
rect 196860 132512 196866 132524
rect 213914 132512 213920 132524
rect 196860 132484 213920 132512
rect 196860 132472 196866 132484
rect 213914 132472 213920 132484
rect 213972 132472 213978 132524
rect 253566 132472 253572 132524
rect 253624 132512 253630 132524
rect 264974 132512 264980 132524
rect 253624 132484 264980 132512
rect 253624 132472 253630 132484
rect 264974 132472 264980 132484
rect 265032 132472 265038 132524
rect 231762 132404 231768 132456
rect 231820 132444 231826 132456
rect 249334 132444 249340 132456
rect 231820 132416 249340 132444
rect 231820 132404 231826 132416
rect 249334 132404 249340 132416
rect 249392 132404 249398 132456
rect 282638 132404 282644 132456
rect 282696 132444 282702 132456
rect 325694 132444 325700 132456
rect 282696 132416 325700 132444
rect 282696 132404 282702 132416
rect 325694 132404 325700 132416
rect 325752 132404 325758 132456
rect 369118 132404 369124 132456
rect 369176 132444 369182 132456
rect 397546 132444 397552 132456
rect 369176 132416 397552 132444
rect 369176 132404 369182 132416
rect 397546 132404 397552 132416
rect 397604 132404 397610 132456
rect 281718 132336 281724 132388
rect 281776 132376 281782 132388
rect 303614 132376 303620 132388
rect 281776 132348 303620 132376
rect 281776 132336 281782 132348
rect 303614 132336 303620 132348
rect 303672 132336 303678 132388
rect 178770 131724 178776 131776
rect 178828 131764 178834 131776
rect 211982 131764 211988 131776
rect 178828 131736 211988 131764
rect 178828 131724 178834 131736
rect 211982 131724 211988 131736
rect 212040 131724 212046 131776
rect 231670 131724 231676 131776
rect 231728 131764 231734 131776
rect 239674 131764 239680 131776
rect 231728 131736 239680 131764
rect 231728 131724 231734 131736
rect 239674 131724 239680 131736
rect 239732 131724 239738 131776
rect 256694 131724 256700 131776
rect 256752 131764 256758 131776
rect 265158 131764 265164 131776
rect 256752 131736 265164 131764
rect 256752 131724 256758 131736
rect 265158 131724 265164 131736
rect 265216 131724 265222 131776
rect 180242 131112 180248 131164
rect 180300 131152 180306 131164
rect 213914 131152 213920 131164
rect 180300 131124 213920 131152
rect 180300 131112 180306 131124
rect 213914 131112 213920 131124
rect 213972 131112 213978 131164
rect 252002 131112 252008 131164
rect 252060 131152 252066 131164
rect 264974 131152 264980 131164
rect 252060 131124 264980 131152
rect 252060 131112 252066 131124
rect 264974 131112 264980 131124
rect 265032 131112 265038 131164
rect 231762 131044 231768 131096
rect 231820 131084 231826 131096
rect 260098 131084 260104 131096
rect 231820 131056 260104 131084
rect 231820 131044 231826 131056
rect 260098 131044 260104 131056
rect 260156 131044 260162 131096
rect 282270 131044 282276 131096
rect 282328 131084 282334 131096
rect 316034 131084 316040 131096
rect 282328 131056 316040 131084
rect 282328 131044 282334 131056
rect 316034 131044 316040 131056
rect 316092 131044 316098 131096
rect 231394 130976 231400 131028
rect 231452 131016 231458 131028
rect 247678 131016 247684 131028
rect 231452 130988 247684 131016
rect 231452 130976 231458 130988
rect 247678 130976 247684 130988
rect 247736 130976 247742 131028
rect 282822 130976 282828 131028
rect 282880 131016 282886 131028
rect 303798 131016 303804 131028
rect 282880 130988 303804 131016
rect 282880 130976 282886 130988
rect 303798 130976 303804 130988
rect 303856 130976 303862 131028
rect 442902 130772 442908 130824
rect 442960 130812 442966 130824
rect 444374 130812 444380 130824
rect 442960 130784 444380 130812
rect 442960 130772 442966 130784
rect 444374 130772 444380 130784
rect 444432 130772 444438 130824
rect 192570 130432 192576 130484
rect 192628 130472 192634 130484
rect 214466 130472 214472 130484
rect 192628 130444 214472 130472
rect 192628 130432 192634 130444
rect 214466 130432 214472 130444
rect 214524 130432 214530 130484
rect 180150 130364 180156 130416
rect 180208 130404 180214 130416
rect 209222 130404 209228 130416
rect 180208 130376 209228 130404
rect 180208 130364 180214 130376
rect 209222 130364 209228 130376
rect 209280 130364 209286 130416
rect 345750 130364 345756 130416
rect 345808 130404 345814 130416
rect 391198 130404 391204 130416
rect 345808 130376 391204 130404
rect 345808 130364 345814 130376
rect 391198 130364 391204 130376
rect 391256 130364 391262 130416
rect 209130 129752 209136 129804
rect 209188 129792 209194 129804
rect 213914 129792 213920 129804
rect 209188 129764 213920 129792
rect 209188 129752 209194 129764
rect 213914 129752 213920 129764
rect 213972 129752 213978 129804
rect 256050 129752 256056 129804
rect 256108 129792 256114 129804
rect 264974 129792 264980 129804
rect 256108 129764 264980 129792
rect 256108 129752 256114 129764
rect 264974 129752 264980 129764
rect 265032 129752 265038 129804
rect 355318 129752 355324 129804
rect 355376 129792 355382 129804
rect 358814 129792 358820 129804
rect 355376 129764 358820 129792
rect 355376 129752 355382 129764
rect 358814 129752 358820 129764
rect 358872 129792 358878 129804
rect 397546 129792 397552 129804
rect 358872 129764 397552 129792
rect 358872 129752 358878 129764
rect 397546 129752 397552 129764
rect 397604 129752 397610 129804
rect 442902 129752 442908 129804
rect 442960 129792 442966 129804
rect 454126 129792 454132 129804
rect 442960 129764 454132 129792
rect 442960 129752 442966 129764
rect 454126 129752 454132 129764
rect 454184 129752 454190 129804
rect 231762 129684 231768 129736
rect 231820 129724 231826 129736
rect 252094 129724 252100 129736
rect 231820 129696 252100 129724
rect 231820 129684 231826 129696
rect 252094 129684 252100 129696
rect 252152 129684 252158 129736
rect 282086 129684 282092 129736
rect 282144 129724 282150 129736
rect 288618 129724 288624 129736
rect 282144 129696 288624 129724
rect 282144 129684 282150 129696
rect 288618 129684 288624 129696
rect 288676 129684 288682 129736
rect 231394 129616 231400 129668
rect 231452 129656 231458 129668
rect 242250 129656 242256 129668
rect 231452 129628 242256 129656
rect 231452 129616 231458 129628
rect 242250 129616 242256 129628
rect 242308 129616 242314 129668
rect 367830 129072 367836 129124
rect 367888 129112 367894 129124
rect 393314 129112 393320 129124
rect 367888 129084 393320 129112
rect 367888 129072 367894 129084
rect 393314 129072 393320 129084
rect 393372 129112 393378 129124
rect 394602 129112 394608 129124
rect 393372 129084 394608 129112
rect 393372 129072 393378 129084
rect 394602 129072 394608 129084
rect 394660 129072 394666 129124
rect 167730 129004 167736 129056
rect 167788 129044 167794 129056
rect 198090 129044 198096 129056
rect 167788 129016 198096 129044
rect 167788 129004 167794 129016
rect 198090 129004 198096 129016
rect 198148 129004 198154 129056
rect 335998 129004 336004 129056
rect 336056 129044 336062 129056
rect 378870 129044 378876 129056
rect 336056 129016 378876 129044
rect 336056 129004 336062 129016
rect 378870 129004 378876 129016
rect 378928 129004 378934 129056
rect 257522 128392 257528 128444
rect 257580 128432 257586 128444
rect 265066 128432 265072 128444
rect 257580 128404 265072 128432
rect 257580 128392 257586 128404
rect 265066 128392 265072 128404
rect 265124 128392 265130 128444
rect 60642 128324 60648 128376
rect 60700 128364 60706 128376
rect 66162 128364 66168 128376
rect 60700 128336 66168 128364
rect 60700 128324 60706 128336
rect 66162 128324 66168 128336
rect 66220 128324 66226 128376
rect 210602 128324 210608 128376
rect 210660 128364 210666 128376
rect 213914 128364 213920 128376
rect 210660 128336 213920 128364
rect 210660 128324 210666 128336
rect 213914 128324 213920 128336
rect 213972 128324 213978 128376
rect 251910 128324 251916 128376
rect 251968 128364 251974 128376
rect 264974 128364 264980 128376
rect 251968 128336 264980 128364
rect 251968 128324 251974 128336
rect 264974 128324 264980 128336
rect 265032 128324 265038 128376
rect 393958 128324 393964 128376
rect 394016 128364 394022 128376
rect 397546 128364 397552 128376
rect 394016 128336 397552 128364
rect 394016 128324 394022 128336
rect 397546 128324 397552 128336
rect 397604 128324 397610 128376
rect 442166 128324 442172 128376
rect 442224 128364 442230 128376
rect 444466 128364 444472 128376
rect 442224 128336 444472 128364
rect 442224 128324 442230 128336
rect 444466 128324 444472 128336
rect 444524 128324 444530 128376
rect 231762 128256 231768 128308
rect 231820 128296 231826 128308
rect 245102 128296 245108 128308
rect 231820 128268 245108 128296
rect 231820 128256 231826 128268
rect 245102 128256 245108 128268
rect 245160 128256 245166 128308
rect 231302 127984 231308 128036
rect 231360 128024 231366 128036
rect 233970 128024 233976 128036
rect 231360 127996 233976 128024
rect 231360 127984 231366 127996
rect 233970 127984 233976 127996
rect 234028 127984 234034 128036
rect 285674 127644 285680 127696
rect 285732 127684 285738 127696
rect 295978 127684 295984 127696
rect 285732 127656 295984 127684
rect 285732 127644 285738 127656
rect 295978 127644 295984 127656
rect 296036 127644 296042 127696
rect 173342 127576 173348 127628
rect 173400 127616 173406 127628
rect 214558 127616 214564 127628
rect 173400 127588 214564 127616
rect 173400 127576 173406 127588
rect 214558 127576 214564 127588
rect 214616 127576 214622 127628
rect 282822 127576 282828 127628
rect 282880 127616 282886 127628
rect 314654 127616 314660 127628
rect 282880 127588 314660 127616
rect 282880 127576 282886 127588
rect 314654 127576 314660 127588
rect 314712 127576 314718 127628
rect 442902 127168 442908 127220
rect 442960 127208 442966 127220
rect 448514 127208 448520 127220
rect 442960 127180 448520 127208
rect 442960 127168 442966 127180
rect 448514 127168 448520 127180
rect 448572 127168 448578 127220
rect 261478 127032 261484 127084
rect 261536 127072 261542 127084
rect 265066 127072 265072 127084
rect 261536 127044 265072 127072
rect 261536 127032 261542 127044
rect 265066 127032 265072 127044
rect 265124 127032 265130 127084
rect 187142 126964 187148 127016
rect 187200 127004 187206 127016
rect 213914 127004 213920 127016
rect 187200 126976 213920 127004
rect 187200 126964 187206 126976
rect 213914 126964 213920 126976
rect 213972 126964 213978 127016
rect 242250 126964 242256 127016
rect 242308 127004 242314 127016
rect 264974 127004 264980 127016
rect 242308 126976 264980 127004
rect 242308 126964 242314 126976
rect 264974 126964 264980 126976
rect 265032 126964 265038 127016
rect 371878 126964 371884 127016
rect 371936 127004 371942 127016
rect 397546 127004 397552 127016
rect 371936 126976 397552 127004
rect 371936 126964 371942 126976
rect 397546 126964 397552 126976
rect 397604 126964 397610 127016
rect 231670 126896 231676 126948
rect 231728 126936 231734 126948
rect 249058 126936 249064 126948
rect 231728 126908 249064 126936
rect 231728 126896 231734 126908
rect 249058 126896 249064 126908
rect 249116 126896 249122 126948
rect 282270 126896 282276 126948
rect 282328 126936 282334 126948
rect 298186 126936 298192 126948
rect 282328 126908 298192 126936
rect 282328 126896 282334 126908
rect 298186 126896 298192 126908
rect 298244 126896 298250 126948
rect 371234 126896 371240 126948
rect 371292 126936 371298 126948
rect 398098 126936 398104 126948
rect 371292 126908 398104 126936
rect 371292 126896 371298 126908
rect 398098 126896 398104 126908
rect 398156 126896 398162 126948
rect 442902 126896 442908 126948
rect 442960 126936 442966 126948
rect 583110 126936 583116 126948
rect 442960 126908 583116 126936
rect 442960 126896 442966 126908
rect 583110 126896 583116 126908
rect 583168 126896 583174 126948
rect 231762 126828 231768 126880
rect 231820 126868 231826 126880
rect 243630 126868 243636 126880
rect 231820 126840 243636 126868
rect 231820 126828 231826 126840
rect 243630 126828 243636 126840
rect 243688 126828 243694 126880
rect 442810 126828 442816 126880
rect 442868 126868 442874 126880
rect 454034 126868 454040 126880
rect 442868 126840 454040 126868
rect 442868 126828 442874 126840
rect 454034 126828 454040 126840
rect 454092 126828 454098 126880
rect 169018 126216 169024 126268
rect 169076 126256 169082 126268
rect 211890 126256 211896 126268
rect 169076 126228 211896 126256
rect 169076 126216 169082 126228
rect 211890 126216 211896 126228
rect 211948 126216 211954 126268
rect 243722 126216 243728 126268
rect 243780 126256 243786 126268
rect 256694 126256 256700 126268
rect 243780 126228 256700 126256
rect 243780 126216 243786 126228
rect 256694 126216 256700 126228
rect 256752 126216 256758 126268
rect 260374 126216 260380 126268
rect 260432 126256 260438 126268
rect 263134 126256 263140 126268
rect 260432 126228 263140 126256
rect 260432 126216 260438 126228
rect 263134 126216 263140 126228
rect 263192 126216 263198 126268
rect 281994 126216 282000 126268
rect 282052 126256 282058 126268
rect 306374 126256 306380 126268
rect 282052 126228 306380 126256
rect 282052 126216 282058 126228
rect 306374 126216 306380 126228
rect 306432 126216 306438 126268
rect 202414 125604 202420 125656
rect 202472 125644 202478 125656
rect 213914 125644 213920 125656
rect 202472 125616 213920 125644
rect 202472 125604 202478 125616
rect 213914 125604 213920 125616
rect 213972 125604 213978 125656
rect 257430 125604 257436 125656
rect 257488 125644 257494 125656
rect 264974 125644 264980 125656
rect 257488 125616 264980 125644
rect 257488 125604 257494 125616
rect 264974 125604 264980 125616
rect 265032 125604 265038 125656
rect 282362 125536 282368 125588
rect 282420 125576 282426 125588
rect 298094 125576 298100 125588
rect 282420 125548 298100 125576
rect 282420 125536 282426 125548
rect 298094 125536 298100 125548
rect 298152 125536 298158 125588
rect 442902 125536 442908 125588
rect 442960 125576 442966 125588
rect 460934 125576 460940 125588
rect 442960 125548 460940 125576
rect 442960 125536 442966 125548
rect 460934 125536 460940 125548
rect 460992 125576 460998 125588
rect 582742 125576 582748 125588
rect 460992 125548 582748 125576
rect 460992 125536 460998 125548
rect 582742 125536 582748 125548
rect 582800 125536 582806 125588
rect 230750 124924 230756 124976
rect 230808 124964 230814 124976
rect 250622 124964 250628 124976
rect 230808 124936 250628 124964
rect 230808 124924 230814 124936
rect 250622 124924 250628 124936
rect 250680 124924 250686 124976
rect 205082 124856 205088 124908
rect 205140 124896 205146 124908
rect 214006 124896 214012 124908
rect 205140 124868 214012 124896
rect 205140 124856 205146 124868
rect 214006 124856 214012 124868
rect 214064 124856 214070 124908
rect 230658 124856 230664 124908
rect 230716 124896 230722 124908
rect 245194 124896 245200 124908
rect 230716 124868 245200 124896
rect 230716 124856 230722 124868
rect 245194 124856 245200 124868
rect 245252 124856 245258 124908
rect 245286 124856 245292 124908
rect 245344 124896 245350 124908
rect 265710 124896 265716 124908
rect 245344 124868 265716 124896
rect 245344 124856 245350 124868
rect 265710 124856 265716 124868
rect 265768 124856 265774 124908
rect 166258 124176 166264 124228
rect 166316 124216 166322 124228
rect 213914 124216 213920 124228
rect 166316 124188 213920 124216
rect 166316 124176 166322 124188
rect 213914 124176 213920 124188
rect 213972 124176 213978 124228
rect 254762 124176 254768 124228
rect 254820 124216 254826 124228
rect 264974 124216 264980 124228
rect 254820 124188 264980 124216
rect 254820 124176 254826 124188
rect 264974 124176 264980 124188
rect 265032 124176 265038 124228
rect 377398 124176 377404 124228
rect 377456 124216 377462 124228
rect 385034 124216 385040 124228
rect 377456 124188 385040 124216
rect 377456 124176 377462 124188
rect 385034 124176 385040 124188
rect 385092 124216 385098 124228
rect 397546 124216 397552 124228
rect 385092 124188 397552 124216
rect 385092 124176 385098 124188
rect 397546 124176 397552 124188
rect 397604 124176 397610 124228
rect 231762 124108 231768 124160
rect 231820 124148 231826 124160
rect 252186 124148 252192 124160
rect 231820 124120 252192 124148
rect 231820 124108 231826 124120
rect 252186 124108 252192 124120
rect 252244 124108 252250 124160
rect 385678 124108 385684 124160
rect 385736 124148 385742 124160
rect 397638 124148 397644 124160
rect 385736 124120 397644 124148
rect 385736 124108 385742 124120
rect 397638 124108 397644 124120
rect 397696 124108 397702 124160
rect 442626 124108 442632 124160
rect 442684 124148 442690 124160
rect 583478 124148 583484 124160
rect 442684 124120 583484 124148
rect 442684 124108 442690 124120
rect 583478 124108 583484 124120
rect 583536 124108 583542 124160
rect 230566 124040 230572 124092
rect 230624 124080 230630 124092
rect 232682 124080 232688 124092
rect 230624 124052 232688 124080
rect 230624 124040 230630 124052
rect 232682 124040 232688 124052
rect 232740 124040 232746 124092
rect 167638 123428 167644 123480
rect 167696 123468 167702 123480
rect 180334 123468 180340 123480
rect 167696 123440 180340 123468
rect 167696 123428 167702 123440
rect 180334 123428 180340 123440
rect 180392 123428 180398 123480
rect 232774 123428 232780 123480
rect 232832 123468 232838 123480
rect 248046 123468 248052 123480
rect 232832 123440 248052 123468
rect 232832 123428 232838 123440
rect 248046 123428 248052 123440
rect 248104 123428 248110 123480
rect 282730 123428 282736 123480
rect 282788 123468 282794 123480
rect 291286 123468 291292 123480
rect 282788 123440 291292 123468
rect 282788 123428 282794 123440
rect 291286 123428 291292 123440
rect 291344 123428 291350 123480
rect 354030 123428 354036 123480
rect 354088 123468 354094 123480
rect 397546 123468 397552 123480
rect 354088 123440 397552 123468
rect 354088 123428 354094 123440
rect 397546 123428 397552 123440
rect 397604 123428 397610 123480
rect 196710 122884 196716 122936
rect 196768 122924 196774 122936
rect 214006 122924 214012 122936
rect 196768 122896 214012 122924
rect 196768 122884 196774 122896
rect 214006 122884 214012 122896
rect 214064 122884 214070 122936
rect 252094 122884 252100 122936
rect 252152 122924 252158 122936
rect 264974 122924 264980 122936
rect 252152 122896 264980 122924
rect 252152 122884 252158 122896
rect 264974 122884 264980 122896
rect 265032 122884 265038 122936
rect 176010 122816 176016 122868
rect 176068 122856 176074 122868
rect 213914 122856 213920 122868
rect 176068 122828 213920 122856
rect 176068 122816 176074 122828
rect 213914 122816 213920 122828
rect 213972 122816 213978 122868
rect 250806 122816 250812 122868
rect 250864 122856 250870 122868
rect 265066 122856 265072 122868
rect 250864 122828 265072 122856
rect 250864 122816 250870 122828
rect 265066 122816 265072 122828
rect 265124 122816 265130 122868
rect 231762 122748 231768 122800
rect 231820 122788 231826 122800
rect 256142 122788 256148 122800
rect 231820 122760 256148 122788
rect 231820 122748 231826 122760
rect 256142 122748 256148 122760
rect 256200 122748 256206 122800
rect 282822 122748 282828 122800
rect 282880 122788 282886 122800
rect 304994 122788 305000 122800
rect 282880 122760 305000 122788
rect 282880 122748 282886 122760
rect 304994 122748 305000 122760
rect 305052 122748 305058 122800
rect 441890 122612 441896 122664
rect 441948 122652 441954 122664
rect 444558 122652 444564 122664
rect 441948 122624 444564 122652
rect 441948 122612 441954 122624
rect 444558 122612 444564 122624
rect 444616 122612 444622 122664
rect 230934 121864 230940 121916
rect 230992 121904 230998 121916
rect 235534 121904 235540 121916
rect 230992 121876 235540 121904
rect 230992 121864 230998 121876
rect 235534 121864 235540 121876
rect 235592 121864 235598 121916
rect 180334 121524 180340 121576
rect 180392 121564 180398 121576
rect 213914 121564 213920 121576
rect 180392 121536 213920 121564
rect 180392 121524 180398 121536
rect 213914 121524 213920 121536
rect 213972 121524 213978 121576
rect 171778 121456 171784 121508
rect 171836 121496 171842 121508
rect 214006 121496 214012 121508
rect 171836 121468 214012 121496
rect 171836 121456 171842 121468
rect 214006 121456 214012 121468
rect 214064 121456 214070 121508
rect 249058 121456 249064 121508
rect 249116 121496 249122 121508
rect 264974 121496 264980 121508
rect 249116 121468 264980 121496
rect 249116 121456 249122 121468
rect 264974 121456 264980 121468
rect 265032 121456 265038 121508
rect 367738 121456 367744 121508
rect 367796 121496 367802 121508
rect 397546 121496 397552 121508
rect 367796 121468 397552 121496
rect 367796 121456 367802 121468
rect 397546 121456 397552 121468
rect 397604 121456 397610 121508
rect 231670 121388 231676 121440
rect 231728 121428 231734 121440
rect 260282 121428 260288 121440
rect 231728 121400 260288 121428
rect 231728 121388 231734 121400
rect 260282 121388 260288 121400
rect 260340 121388 260346 121440
rect 282822 121388 282828 121440
rect 282880 121428 282886 121440
rect 289998 121428 290004 121440
rect 282880 121400 290004 121428
rect 282880 121388 282886 121400
rect 289998 121388 290004 121400
rect 290056 121388 290062 121440
rect 387058 121388 387064 121440
rect 387116 121428 387122 121440
rect 397638 121428 397644 121440
rect 387116 121400 397644 121428
rect 387116 121388 387122 121400
rect 397638 121388 397644 121400
rect 397696 121388 397702 121440
rect 231762 121320 231768 121372
rect 231820 121360 231826 121372
rect 240778 121360 240784 121372
rect 231820 121332 240784 121360
rect 231820 121320 231826 121332
rect 240778 121320 240784 121332
rect 240836 121320 240842 121372
rect 191190 120164 191196 120216
rect 191248 120204 191254 120216
rect 214006 120204 214012 120216
rect 191248 120176 214012 120204
rect 191248 120164 191254 120176
rect 214006 120164 214012 120176
rect 214064 120164 214070 120216
rect 260098 120164 260104 120216
rect 260156 120204 260162 120216
rect 265066 120204 265072 120216
rect 260156 120176 265072 120204
rect 260156 120164 260162 120176
rect 265066 120164 265072 120176
rect 265124 120164 265130 120216
rect 166350 120096 166356 120148
rect 166408 120136 166414 120148
rect 213914 120136 213920 120148
rect 166408 120108 213920 120136
rect 166408 120096 166414 120108
rect 213914 120096 213920 120108
rect 213972 120096 213978 120148
rect 262766 120096 262772 120148
rect 262824 120136 262830 120148
rect 264974 120136 264980 120148
rect 262824 120108 264980 120136
rect 262824 120096 262830 120108
rect 264974 120096 264980 120108
rect 265032 120096 265038 120148
rect 231762 120028 231768 120080
rect 231820 120068 231826 120080
rect 241054 120068 241060 120080
rect 231820 120040 241060 120068
rect 231820 120028 231826 120040
rect 241054 120028 241060 120040
rect 241112 120028 241118 120080
rect 282822 120028 282828 120080
rect 282880 120068 282886 120080
rect 292574 120068 292580 120080
rect 282880 120040 292580 120068
rect 282880 120028 282886 120040
rect 292574 120028 292580 120040
rect 292632 120028 292638 120080
rect 338850 120028 338856 120080
rect 338908 120068 338914 120080
rect 397638 120068 397644 120080
rect 338908 120040 397644 120068
rect 338908 120028 338914 120040
rect 397638 120028 397644 120040
rect 397696 120028 397702 120080
rect 385770 119960 385776 120012
rect 385828 120000 385834 120012
rect 397546 120000 397552 120012
rect 385828 119972 397552 120000
rect 385828 119960 385834 119972
rect 397546 119960 397552 119972
rect 397604 119960 397610 120012
rect 231026 119892 231032 119944
rect 231084 119932 231090 119944
rect 238294 119932 238300 119944
rect 231084 119904 238300 119932
rect 231084 119892 231090 119904
rect 238294 119892 238300 119904
rect 238352 119892 238358 119944
rect 240870 119348 240876 119400
rect 240928 119388 240934 119400
rect 258902 119388 258908 119400
rect 240928 119360 258908 119388
rect 240928 119348 240934 119360
rect 258902 119348 258908 119360
rect 258960 119348 258966 119400
rect 192570 118736 192576 118788
rect 192628 118776 192634 118788
rect 213914 118776 213920 118788
rect 192628 118748 213920 118776
rect 192628 118736 192634 118748
rect 213914 118736 213920 118748
rect 213972 118736 213978 118788
rect 258718 118736 258724 118788
rect 258776 118776 258782 118788
rect 265066 118776 265072 118788
rect 258776 118748 265072 118776
rect 258776 118736 258782 118748
rect 265066 118736 265072 118748
rect 265124 118736 265130 118788
rect 174630 118668 174636 118720
rect 174688 118708 174694 118720
rect 214006 118708 214012 118720
rect 174688 118680 214012 118708
rect 174688 118668 174694 118680
rect 214006 118668 214012 118680
rect 214064 118668 214070 118720
rect 240778 118668 240784 118720
rect 240836 118708 240842 118720
rect 264974 118708 264980 118720
rect 240836 118680 264980 118708
rect 240836 118668 240842 118680
rect 264974 118668 264980 118680
rect 265032 118668 265038 118720
rect 231762 118600 231768 118652
rect 231820 118640 231826 118652
rect 267274 118640 267280 118652
rect 231820 118612 267280 118640
rect 231820 118600 231826 118612
rect 267274 118600 267280 118612
rect 267332 118600 267338 118652
rect 352650 118600 352656 118652
rect 352708 118640 352714 118652
rect 397546 118640 397552 118652
rect 352708 118612 397552 118640
rect 352708 118600 352714 118612
rect 397546 118600 397552 118612
rect 397604 118600 397610 118652
rect 442902 118532 442908 118584
rect 442960 118572 442966 118584
rect 445846 118572 445852 118584
rect 442960 118544 445852 118572
rect 442960 118532 442966 118544
rect 445846 118532 445852 118544
rect 445904 118532 445910 118584
rect 230934 118396 230940 118448
rect 230992 118436 230998 118448
rect 236730 118436 236736 118448
rect 230992 118408 236736 118436
rect 230992 118396 230998 118408
rect 236730 118396 236736 118408
rect 236788 118396 236794 118448
rect 282546 118396 282552 118448
rect 282604 118436 282610 118448
rect 285766 118436 285772 118448
rect 282604 118408 285772 118436
rect 282604 118396 282610 118408
rect 285766 118396 285772 118408
rect 285824 118396 285830 118448
rect 177390 117988 177396 118040
rect 177448 118028 177454 118040
rect 188338 118028 188344 118040
rect 177448 118000 188344 118028
rect 177448 117988 177454 118000
rect 188338 117988 188344 118000
rect 188396 117988 188402 118040
rect 173158 117920 173164 117972
rect 173216 117960 173222 117972
rect 191098 117960 191104 117972
rect 173216 117932 191104 117960
rect 173216 117920 173222 117932
rect 191098 117920 191104 117932
rect 191156 117920 191162 117972
rect 236914 117920 236920 117972
rect 236972 117960 236978 117972
rect 248414 117960 248420 117972
rect 236972 117932 248420 117960
rect 236972 117920 236978 117932
rect 248414 117920 248420 117932
rect 248472 117920 248478 117972
rect 282178 117920 282184 117972
rect 282236 117960 282242 117972
rect 296714 117960 296720 117972
rect 282236 117932 296720 117960
rect 282236 117920 282242 117932
rect 296714 117920 296720 117932
rect 296772 117920 296778 117972
rect 338114 117512 338120 117564
rect 338172 117552 338178 117564
rect 340230 117552 340236 117564
rect 338172 117524 340236 117552
rect 338172 117512 338178 117524
rect 340230 117512 340236 117524
rect 340288 117512 340294 117564
rect 198090 117376 198096 117428
rect 198148 117416 198154 117428
rect 213914 117416 213920 117428
rect 198148 117388 213920 117416
rect 198148 117376 198154 117388
rect 213914 117376 213920 117388
rect 213972 117376 213978 117428
rect 194042 117308 194048 117360
rect 194100 117348 194106 117360
rect 214006 117348 214012 117360
rect 194100 117320 214012 117348
rect 194100 117308 194106 117320
rect 214006 117308 214012 117320
rect 214064 117308 214070 117360
rect 253474 117308 253480 117360
rect 253532 117348 253538 117360
rect 264974 117348 264980 117360
rect 253532 117320 264980 117348
rect 253532 117308 253538 117320
rect 264974 117308 264980 117320
rect 265032 117308 265038 117360
rect 374730 117308 374736 117360
rect 374788 117348 374794 117360
rect 397638 117348 397644 117360
rect 374788 117320 397644 117348
rect 374788 117308 374794 117320
rect 397638 117308 397644 117320
rect 397696 117308 397702 117360
rect 231486 117240 231492 117292
rect 231544 117280 231550 117292
rect 242158 117280 242164 117292
rect 231544 117252 242164 117280
rect 231544 117240 231550 117252
rect 242158 117240 242164 117252
rect 242216 117240 242222 117292
rect 320910 117240 320916 117292
rect 320968 117280 320974 117292
rect 395890 117280 395896 117292
rect 320968 117252 395896 117280
rect 320968 117240 320974 117252
rect 395890 117240 395896 117252
rect 395948 117280 395954 117292
rect 397546 117280 397552 117292
rect 395948 117252 397552 117280
rect 395948 117240 395954 117252
rect 397546 117240 397552 117252
rect 397604 117240 397610 117292
rect 235534 116560 235540 116612
rect 235592 116600 235598 116612
rect 253566 116600 253572 116612
rect 235592 116572 253572 116600
rect 235592 116560 235598 116572
rect 253566 116560 253572 116572
rect 253624 116560 253630 116612
rect 282270 116560 282276 116612
rect 282328 116600 282334 116612
rect 307754 116600 307760 116612
rect 282328 116572 307760 116600
rect 282328 116560 282334 116572
rect 307754 116560 307760 116572
rect 307812 116560 307818 116612
rect 442902 116288 442908 116340
rect 442960 116328 442966 116340
rect 449894 116328 449900 116340
rect 442960 116300 449900 116328
rect 442960 116288 442966 116300
rect 449894 116288 449900 116300
rect 449952 116288 449958 116340
rect 282822 116084 282828 116136
rect 282880 116124 282886 116136
rect 287146 116124 287152 116136
rect 282880 116096 287152 116124
rect 282880 116084 282886 116096
rect 287146 116084 287152 116096
rect 287204 116084 287210 116136
rect 188430 116016 188436 116068
rect 188488 116056 188494 116068
rect 213914 116056 213920 116068
rect 188488 116028 213920 116056
rect 188488 116016 188494 116028
rect 213914 116016 213920 116028
rect 213972 116016 213978 116068
rect 170582 115948 170588 116000
rect 170640 115988 170646 116000
rect 214006 115988 214012 116000
rect 170640 115960 214012 115988
rect 170640 115948 170646 115960
rect 214006 115948 214012 115960
rect 214064 115948 214070 116000
rect 253290 115948 253296 116000
rect 253348 115988 253354 116000
rect 264974 115988 264980 116000
rect 253348 115960 264980 115988
rect 253348 115948 253354 115960
rect 264974 115948 264980 115960
rect 265032 115948 265038 116000
rect 231486 115880 231492 115932
rect 231544 115920 231550 115932
rect 246482 115920 246488 115932
rect 231544 115892 246488 115920
rect 231544 115880 231550 115892
rect 246482 115880 246488 115892
rect 246540 115880 246546 115932
rect 282454 115880 282460 115932
rect 282512 115920 282518 115932
rect 309134 115920 309140 115932
rect 282512 115892 309140 115920
rect 282512 115880 282518 115892
rect 309134 115880 309140 115892
rect 309192 115880 309198 115932
rect 358170 115880 358176 115932
rect 358228 115920 358234 115932
rect 397546 115920 397552 115932
rect 358228 115892 397552 115920
rect 358228 115880 358234 115892
rect 397546 115880 397552 115892
rect 397604 115880 397610 115932
rect 392670 115812 392676 115864
rect 392728 115852 392734 115864
rect 397638 115852 397644 115864
rect 392728 115824 397644 115852
rect 392728 115812 392734 115824
rect 397638 115812 397644 115824
rect 397696 115812 397702 115864
rect 442902 115812 442908 115864
rect 442960 115852 442966 115864
rect 447318 115852 447324 115864
rect 442960 115824 447324 115852
rect 442960 115812 442966 115824
rect 447318 115812 447324 115824
rect 447376 115812 447382 115864
rect 230658 114928 230664 114980
rect 230716 114968 230722 114980
rect 233878 114968 233884 114980
rect 230716 114940 233884 114968
rect 230716 114928 230722 114940
rect 233878 114928 233884 114940
rect 233936 114928 233942 114980
rect 195330 114588 195336 114640
rect 195388 114628 195394 114640
rect 213914 114628 213920 114640
rect 195388 114600 213920 114628
rect 195388 114588 195394 114600
rect 213914 114588 213920 114600
rect 213972 114588 213978 114640
rect 250530 114588 250536 114640
rect 250588 114628 250594 114640
rect 265066 114628 265072 114640
rect 250588 114600 265072 114628
rect 250588 114588 250594 114600
rect 265066 114588 265072 114600
rect 265124 114588 265130 114640
rect 169202 114520 169208 114572
rect 169260 114560 169266 114572
rect 214006 114560 214012 114572
rect 169260 114532 214012 114560
rect 169260 114520 169266 114532
rect 214006 114520 214012 114532
rect 214064 114520 214070 114572
rect 242158 114520 242164 114572
rect 242216 114560 242222 114572
rect 264974 114560 264980 114572
rect 242216 114532 264980 114560
rect 242216 114520 242222 114532
rect 264974 114520 264980 114532
rect 265032 114520 265038 114572
rect 231762 114452 231768 114504
rect 231820 114492 231826 114504
rect 250438 114492 250444 114504
rect 231820 114464 250444 114492
rect 231820 114452 231826 114464
rect 250438 114452 250444 114464
rect 250496 114452 250502 114504
rect 282822 114452 282828 114504
rect 282880 114492 282886 114504
rect 290090 114492 290096 114504
rect 282880 114464 290096 114492
rect 282880 114452 282886 114464
rect 290090 114452 290096 114464
rect 290148 114452 290154 114504
rect 352558 114452 352564 114504
rect 352616 114492 352622 114504
rect 397546 114492 397552 114504
rect 352616 114464 397552 114492
rect 352616 114452 352622 114464
rect 397546 114452 397552 114464
rect 397604 114452 397610 114504
rect 231670 114384 231676 114436
rect 231728 114424 231734 114436
rect 243814 114424 243820 114436
rect 231728 114396 243820 114424
rect 231728 114384 231734 114396
rect 243814 114384 243820 114396
rect 243872 114384 243878 114436
rect 384298 114384 384304 114436
rect 384356 114424 384362 114436
rect 397638 114424 397644 114436
rect 384356 114396 397644 114424
rect 384356 114384 384362 114396
rect 397638 114384 397644 114396
rect 397696 114384 397702 114436
rect 177574 113840 177580 113892
rect 177632 113880 177638 113892
rect 202138 113880 202144 113892
rect 177632 113852 202144 113880
rect 177632 113840 177638 113852
rect 202138 113840 202144 113852
rect 202196 113840 202202 113892
rect 164878 113772 164884 113824
rect 164936 113812 164942 113824
rect 214742 113812 214748 113824
rect 164936 113784 214748 113812
rect 164936 113772 164942 113784
rect 214742 113772 214748 113784
rect 214800 113772 214806 113824
rect 442902 113364 442908 113416
rect 442960 113404 442966 113416
rect 444374 113404 444380 113416
rect 442960 113376 444380 113404
rect 442960 113364 442966 113376
rect 444374 113364 444380 113376
rect 444432 113364 444438 113416
rect 207750 113160 207756 113212
rect 207808 113200 207814 113212
rect 213914 113200 213920 113212
rect 207808 113172 213920 113200
rect 207808 113160 207814 113172
rect 213914 113160 213920 113172
rect 213972 113160 213978 113212
rect 245102 113160 245108 113212
rect 245160 113200 245166 113212
rect 264974 113200 264980 113212
rect 245160 113172 264980 113200
rect 245160 113160 245166 113172
rect 264974 113160 264980 113172
rect 265032 113160 265038 113212
rect 231762 113092 231768 113144
rect 231820 113132 231826 113144
rect 264422 113132 264428 113144
rect 231820 113104 264428 113132
rect 231820 113092 231826 113104
rect 264422 113092 264428 113104
rect 264480 113092 264486 113144
rect 282822 113092 282828 113144
rect 282880 113132 282886 113144
rect 303706 113132 303712 113144
rect 282880 113104 303712 113132
rect 282880 113092 282886 113104
rect 303706 113092 303712 113104
rect 303764 113092 303770 113144
rect 309870 113092 309876 113144
rect 309928 113132 309934 113144
rect 397546 113132 397552 113144
rect 309928 113104 397552 113132
rect 309928 113092 309934 113104
rect 397546 113092 397552 113104
rect 397604 113092 397610 113144
rect 442902 113092 442908 113144
rect 442960 113132 442966 113144
rect 456794 113132 456800 113144
rect 442960 113104 456800 113132
rect 442960 113092 442966 113104
rect 456794 113092 456800 113104
rect 456852 113092 456858 113144
rect 230934 113024 230940 113076
rect 230992 113064 230998 113076
rect 253198 113064 253204 113076
rect 230992 113036 253204 113064
rect 230992 113024 230998 113036
rect 253198 113024 253204 113036
rect 253256 113024 253262 113076
rect 281810 113024 281816 113076
rect 281868 113064 281874 113076
rect 284478 113064 284484 113076
rect 281868 113036 284484 113064
rect 281868 113024 281874 113036
rect 284478 113024 284484 113036
rect 284536 113024 284542 113076
rect 388530 112412 388536 112464
rect 388588 112452 388594 112464
rect 398742 112452 398748 112464
rect 388588 112424 398748 112452
rect 388588 112412 388594 112424
rect 398742 112412 398748 112424
rect 398800 112412 398806 112464
rect 202598 111868 202604 111920
rect 202656 111908 202662 111920
rect 214006 111908 214012 111920
rect 202656 111880 214012 111908
rect 202656 111868 202662 111880
rect 214006 111868 214012 111880
rect 214064 111868 214070 111920
rect 166534 111800 166540 111852
rect 166592 111840 166598 111852
rect 213914 111840 213920 111852
rect 166592 111812 213920 111840
rect 166592 111800 166598 111812
rect 213914 111800 213920 111812
rect 213972 111800 213978 111852
rect 261570 111800 261576 111852
rect 261628 111840 261634 111852
rect 264974 111840 264980 111852
rect 261628 111812 264980 111840
rect 261628 111800 261634 111812
rect 264974 111800 264980 111812
rect 265032 111800 265038 111852
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 32398 111772 32404 111784
rect 3200 111744 32404 111772
rect 3200 111732 3206 111744
rect 32398 111732 32404 111744
rect 32456 111732 32462 111784
rect 231762 111732 231768 111784
rect 231820 111772 231826 111784
rect 249242 111772 249248 111784
rect 231820 111744 249248 111772
rect 231820 111732 231826 111744
rect 249242 111732 249248 111744
rect 249300 111732 249306 111784
rect 378778 111732 378784 111784
rect 378836 111772 378842 111784
rect 397454 111772 397460 111784
rect 378836 111744 397460 111772
rect 378836 111732 378842 111744
rect 397454 111732 397460 111744
rect 397512 111732 397518 111784
rect 282822 111528 282828 111580
rect 282880 111568 282886 111580
rect 287054 111568 287060 111580
rect 282880 111540 287060 111568
rect 282880 111528 282886 111540
rect 287054 111528 287060 111540
rect 287112 111528 287118 111580
rect 281534 111392 281540 111444
rect 281592 111432 281598 111444
rect 284570 111432 284576 111444
rect 281592 111404 284576 111432
rect 281592 111392 281598 111404
rect 284570 111392 284576 111404
rect 284628 111392 284634 111444
rect 230750 110848 230756 110900
rect 230808 110888 230814 110900
rect 238110 110888 238116 110900
rect 230808 110860 238116 110888
rect 230808 110848 230814 110860
rect 238110 110848 238116 110860
rect 238168 110848 238174 110900
rect 181622 110508 181628 110560
rect 181680 110548 181686 110560
rect 213914 110548 213920 110560
rect 181680 110520 213920 110548
rect 181680 110508 181686 110520
rect 213914 110508 213920 110520
rect 213972 110508 213978 110560
rect 256234 110508 256240 110560
rect 256292 110548 256298 110560
rect 264974 110548 264980 110560
rect 256292 110520 264980 110548
rect 256292 110508 256298 110520
rect 264974 110508 264980 110520
rect 265032 110508 265038 110560
rect 170490 110440 170496 110492
rect 170548 110480 170554 110492
rect 214006 110480 214012 110492
rect 170548 110452 214012 110480
rect 170548 110440 170554 110452
rect 214006 110440 214012 110452
rect 214064 110440 214070 110492
rect 247678 110440 247684 110492
rect 247736 110480 247742 110492
rect 265066 110480 265072 110492
rect 247736 110452 265072 110480
rect 247736 110440 247742 110452
rect 265066 110440 265072 110452
rect 265124 110440 265130 110492
rect 231670 110372 231676 110424
rect 231728 110412 231734 110424
rect 262950 110412 262956 110424
rect 231728 110384 262956 110412
rect 231728 110372 231734 110384
rect 262950 110372 262956 110384
rect 263008 110372 263014 110424
rect 282822 110372 282828 110424
rect 282880 110412 282886 110424
rect 295426 110412 295432 110424
rect 282880 110384 295432 110412
rect 282880 110372 282886 110384
rect 295426 110372 295432 110384
rect 295484 110372 295490 110424
rect 231762 110304 231768 110356
rect 231820 110344 231826 110356
rect 244918 110344 244924 110356
rect 231820 110316 244924 110344
rect 231820 110304 231826 110316
rect 244918 110304 244924 110316
rect 244976 110304 244982 110356
rect 177666 109080 177672 109132
rect 177724 109120 177730 109132
rect 214006 109120 214012 109132
rect 177724 109092 214012 109120
rect 177724 109080 177730 109092
rect 214006 109080 214012 109092
rect 214064 109080 214070 109132
rect 167638 109012 167644 109064
rect 167696 109052 167702 109064
rect 213914 109052 213920 109064
rect 167696 109024 213920 109052
rect 167696 109012 167702 109024
rect 213914 109012 213920 109024
rect 213972 109012 213978 109064
rect 260282 109012 260288 109064
rect 260340 109052 260346 109064
rect 265066 109052 265072 109064
rect 260340 109024 265072 109052
rect 260340 109012 260346 109024
rect 265066 109012 265072 109024
rect 265124 109012 265130 109064
rect 354030 109012 354036 109064
rect 354088 109052 354094 109064
rect 397546 109052 397552 109064
rect 354088 109024 397552 109052
rect 354088 109012 354094 109024
rect 397546 109012 397552 109024
rect 397604 109012 397610 109064
rect 442166 109012 442172 109064
rect 442224 109052 442230 109064
rect 443362 109052 443368 109064
rect 442224 109024 443368 109052
rect 442224 109012 442230 109024
rect 443362 109012 443368 109024
rect 443420 109012 443426 109064
rect 167546 108944 167552 108996
rect 167604 108984 167610 108996
rect 170674 108984 170680 108996
rect 167604 108956 170680 108984
rect 167604 108944 167610 108956
rect 170674 108944 170680 108956
rect 170732 108944 170738 108996
rect 231762 108944 231768 108996
rect 231820 108984 231826 108996
rect 242342 108984 242348 108996
rect 231820 108956 242348 108984
rect 231820 108944 231826 108956
rect 242342 108944 242348 108956
rect 242400 108944 242406 108996
rect 282362 108944 282368 108996
rect 282420 108984 282426 108996
rect 305086 108984 305092 108996
rect 282420 108956 305092 108984
rect 282420 108944 282426 108956
rect 305086 108944 305092 108956
rect 305144 108944 305150 108996
rect 389818 108944 389824 108996
rect 389876 108984 389882 108996
rect 397454 108984 397460 108996
rect 389876 108956 397460 108984
rect 389876 108944 389882 108956
rect 397454 108944 397460 108956
rect 397512 108944 397518 108996
rect 442442 108944 442448 108996
rect 442500 108984 442506 108996
rect 443270 108984 443276 108996
rect 442500 108956 443276 108984
rect 442500 108944 442506 108956
rect 443270 108944 443276 108956
rect 443328 108944 443334 108996
rect 231302 108876 231308 108928
rect 231360 108916 231366 108928
rect 235442 108916 235448 108928
rect 231360 108888 235448 108916
rect 231360 108876 231366 108888
rect 235442 108876 235448 108888
rect 235500 108876 235506 108928
rect 378778 108264 378784 108316
rect 378836 108304 378842 108316
rect 397638 108304 397644 108316
rect 378836 108276 397644 108304
rect 378836 108264 378842 108276
rect 397638 108264 397644 108276
rect 397696 108264 397702 108316
rect 203702 107720 203708 107772
rect 203760 107760 203766 107772
rect 213914 107760 213920 107772
rect 203760 107732 213920 107760
rect 203760 107720 203766 107732
rect 213914 107720 213920 107732
rect 213972 107720 213978 107772
rect 170766 107652 170772 107704
rect 170824 107692 170830 107704
rect 214006 107692 214012 107704
rect 170824 107664 214012 107692
rect 170824 107652 170830 107664
rect 214006 107652 214012 107664
rect 214064 107652 214070 107704
rect 253198 107652 253204 107704
rect 253256 107692 253262 107704
rect 264974 107692 264980 107704
rect 253256 107664 264980 107692
rect 253256 107652 253262 107664
rect 264974 107652 264980 107664
rect 265032 107652 265038 107704
rect 231762 107584 231768 107636
rect 231820 107624 231826 107636
rect 264514 107624 264520 107636
rect 231820 107596 264520 107624
rect 231820 107584 231826 107596
rect 264514 107584 264520 107596
rect 264572 107584 264578 107636
rect 282822 107584 282828 107636
rect 282880 107624 282886 107636
rect 291194 107624 291200 107636
rect 282880 107596 291200 107624
rect 282880 107584 282886 107596
rect 291194 107584 291200 107596
rect 291252 107584 291258 107636
rect 231670 107516 231676 107568
rect 231728 107556 231734 107568
rect 263042 107556 263048 107568
rect 231728 107528 263048 107556
rect 231728 107516 231734 107528
rect 263042 107516 263048 107528
rect 263100 107516 263106 107568
rect 298094 106904 298100 106956
rect 298152 106944 298158 106956
rect 367830 106944 367836 106956
rect 298152 106916 367836 106944
rect 298152 106904 298158 106916
rect 367830 106904 367836 106916
rect 367888 106904 367894 106956
rect 185762 106360 185768 106412
rect 185820 106400 185826 106412
rect 213914 106400 213920 106412
rect 185820 106372 213920 106400
rect 185820 106360 185826 106372
rect 213914 106360 213920 106372
rect 213972 106360 213978 106412
rect 377398 106360 377404 106412
rect 377456 106400 377462 106412
rect 397454 106400 397460 106412
rect 377456 106372 397460 106400
rect 377456 106360 377462 106372
rect 397454 106360 397460 106372
rect 397512 106360 397518 106412
rect 166442 106292 166448 106344
rect 166500 106332 166506 106344
rect 214006 106332 214012 106344
rect 166500 106304 214012 106332
rect 166500 106292 166506 106304
rect 214006 106292 214012 106304
rect 214064 106292 214070 106344
rect 262950 106292 262956 106344
rect 263008 106332 263014 106344
rect 265250 106332 265256 106344
rect 263008 106304 265256 106332
rect 263008 106292 263014 106304
rect 265250 106292 265256 106304
rect 265308 106292 265314 106344
rect 370590 106292 370596 106344
rect 370648 106332 370654 106344
rect 397546 106332 397552 106344
rect 370648 106304 397552 106332
rect 370648 106292 370654 106304
rect 397546 106292 397552 106304
rect 397604 106292 397610 106344
rect 231302 106224 231308 106276
rect 231360 106264 231366 106276
rect 240962 106264 240968 106276
rect 231360 106236 240968 106264
rect 231360 106224 231366 106236
rect 240962 106224 240968 106236
rect 241020 106224 241026 106276
rect 294690 106224 294696 106276
rect 294748 106264 294754 106276
rect 397454 106264 397460 106276
rect 294748 106236 397460 106264
rect 294748 106224 294754 106236
rect 397454 106224 397460 106236
rect 397512 106224 397518 106276
rect 442718 106224 442724 106276
rect 442776 106264 442782 106276
rect 452654 106264 452660 106276
rect 442776 106236 452660 106264
rect 442776 106224 442782 106236
rect 452654 106224 452660 106236
rect 452712 106224 452718 106276
rect 231578 106156 231584 106208
rect 231636 106196 231642 106208
rect 234062 106196 234068 106208
rect 231636 106168 234068 106196
rect 231636 106156 231642 106168
rect 234062 106156 234068 106168
rect 234120 106156 234126 106208
rect 173434 105544 173440 105596
rect 173492 105584 173498 105596
rect 202598 105584 202604 105596
rect 173492 105556 202604 105584
rect 173492 105544 173498 105556
rect 202598 105544 202604 105556
rect 202656 105544 202662 105596
rect 236730 105544 236736 105596
rect 236788 105584 236794 105596
rect 246574 105584 246580 105596
rect 236788 105556 246580 105584
rect 236788 105544 236794 105556
rect 246574 105544 246580 105556
rect 246632 105544 246638 105596
rect 374638 105544 374644 105596
rect 374696 105584 374702 105596
rect 397914 105584 397920 105596
rect 374696 105556 397920 105584
rect 374696 105544 374702 105556
rect 397914 105544 397920 105556
rect 397972 105544 397978 105596
rect 231210 105068 231216 105120
rect 231268 105108 231274 105120
rect 231486 105108 231492 105120
rect 231268 105080 231492 105108
rect 231268 105068 231274 105080
rect 231486 105068 231492 105080
rect 231544 105068 231550 105120
rect 202322 104932 202328 104984
rect 202380 104972 202386 104984
rect 213914 104972 213920 104984
rect 202380 104944 213920 104972
rect 202380 104932 202386 104944
rect 213914 104932 213920 104944
rect 213972 104932 213978 104984
rect 263318 104932 263324 104984
rect 263376 104972 263382 104984
rect 265158 104972 265164 104984
rect 263376 104944 265164 104972
rect 263376 104932 263382 104944
rect 265158 104932 265164 104944
rect 265216 104932 265222 104984
rect 178678 104864 178684 104916
rect 178736 104904 178742 104916
rect 214006 104904 214012 104916
rect 178736 104876 214012 104904
rect 178736 104864 178742 104876
rect 214006 104864 214012 104876
rect 214064 104864 214070 104916
rect 245194 104864 245200 104916
rect 245252 104904 245258 104916
rect 264974 104904 264980 104916
rect 245252 104876 264980 104904
rect 245252 104864 245258 104876
rect 264974 104864 264980 104876
rect 265032 104864 265038 104916
rect 442350 104864 442356 104916
rect 442408 104904 442414 104916
rect 445846 104904 445852 104916
rect 442408 104876 445852 104904
rect 442408 104864 442414 104876
rect 445846 104864 445852 104876
rect 445904 104864 445910 104916
rect 231762 104796 231768 104848
rect 231820 104836 231826 104848
rect 247862 104836 247868 104848
rect 231820 104808 247868 104836
rect 231820 104796 231826 104808
rect 247862 104796 247868 104808
rect 247920 104796 247926 104848
rect 281534 104796 281540 104848
rect 281592 104836 281598 104848
rect 284386 104836 284392 104848
rect 281592 104808 284392 104836
rect 281592 104796 281598 104808
rect 284386 104796 284392 104808
rect 284444 104796 284450 104848
rect 347038 104796 347044 104848
rect 347096 104836 347102 104848
rect 397454 104836 397460 104848
rect 347096 104808 397460 104836
rect 347096 104796 347102 104808
rect 397454 104796 397460 104808
rect 397512 104796 397518 104848
rect 391198 104728 391204 104780
rect 391256 104768 391262 104780
rect 397546 104768 397552 104780
rect 391256 104740 397552 104768
rect 391256 104728 391262 104740
rect 397546 104728 397552 104740
rect 397604 104728 397610 104780
rect 231670 104660 231676 104712
rect 231728 104700 231734 104712
rect 236822 104700 236828 104712
rect 231728 104672 236828 104700
rect 231728 104660 231734 104672
rect 236822 104660 236828 104672
rect 236880 104660 236886 104712
rect 167730 104184 167736 104236
rect 167788 104224 167794 104236
rect 185670 104224 185676 104236
rect 167788 104196 185676 104224
rect 167788 104184 167794 104196
rect 185670 104184 185676 104196
rect 185728 104184 185734 104236
rect 171962 104116 171968 104168
rect 172020 104156 172026 104168
rect 195422 104156 195428 104168
rect 172020 104128 195428 104156
rect 172020 104116 172026 104128
rect 195422 104116 195428 104128
rect 195480 104116 195486 104168
rect 263042 104116 263048 104168
rect 263100 104156 263106 104168
rect 265066 104156 265072 104168
rect 263100 104128 265072 104156
rect 263100 104116 263106 104128
rect 265066 104116 265072 104128
rect 265124 104116 265130 104168
rect 238110 103504 238116 103556
rect 238168 103544 238174 103556
rect 264974 103544 264980 103556
rect 238168 103516 264980 103544
rect 238168 103504 238174 103516
rect 264974 103504 264980 103516
rect 265032 103504 265038 103556
rect 230750 103436 230756 103488
rect 230808 103476 230814 103488
rect 249150 103476 249156 103488
rect 230808 103448 249156 103476
rect 230808 103436 230814 103448
rect 249150 103436 249156 103448
rect 249208 103436 249214 103488
rect 359458 103436 359464 103488
rect 359516 103476 359522 103488
rect 397454 103476 397460 103488
rect 359516 103448 397460 103476
rect 359516 103436 359522 103448
rect 397454 103436 397460 103448
rect 397512 103436 397518 103488
rect 231302 102824 231308 102876
rect 231360 102864 231366 102876
rect 235350 102864 235356 102876
rect 231360 102836 235356 102864
rect 231360 102824 231366 102836
rect 235350 102824 235356 102836
rect 235408 102824 235414 102876
rect 256142 102756 256148 102808
rect 256200 102796 256206 102808
rect 263318 102796 263324 102808
rect 256200 102768 263324 102796
rect 256200 102756 256206 102768
rect 263318 102756 263324 102768
rect 263376 102756 263382 102808
rect 325050 102756 325056 102808
rect 325108 102796 325114 102808
rect 366910 102796 366916 102808
rect 325108 102768 366916 102796
rect 325108 102756 325114 102768
rect 366910 102756 366916 102768
rect 366968 102756 366974 102808
rect 198182 102144 198188 102196
rect 198240 102184 198246 102196
rect 213914 102184 213920 102196
rect 198240 102156 213920 102184
rect 198240 102144 198246 102156
rect 213914 102144 213920 102156
rect 213972 102144 213978 102196
rect 249242 102144 249248 102196
rect 249300 102184 249306 102196
rect 264974 102184 264980 102196
rect 249300 102156 264980 102184
rect 249300 102144 249306 102156
rect 264974 102144 264980 102156
rect 265032 102144 265038 102196
rect 449158 102076 449164 102128
rect 449216 102116 449222 102128
rect 583202 102116 583208 102128
rect 449216 102088 583208 102116
rect 449216 102076 449222 102088
rect 583202 102076 583208 102088
rect 583260 102076 583266 102128
rect 231578 102008 231584 102060
rect 231636 102048 231642 102060
rect 257614 102048 257620 102060
rect 231636 102020 257620 102048
rect 231636 102008 231642 102020
rect 257614 102008 257620 102020
rect 257672 102008 257678 102060
rect 230566 101872 230572 101924
rect 230624 101912 230630 101924
rect 232590 101912 232596 101924
rect 230624 101884 232596 101912
rect 230624 101872 230630 101884
rect 232590 101872 232596 101884
rect 232648 101872 232654 101924
rect 442166 101600 442172 101652
rect 442224 101640 442230 101652
rect 445938 101640 445944 101652
rect 442224 101612 445944 101640
rect 442224 101600 442230 101612
rect 445938 101600 445944 101612
rect 445996 101600 446002 101652
rect 363690 101532 363696 101584
rect 363748 101572 363754 101584
rect 439314 101572 439320 101584
rect 363748 101544 439320 101572
rect 363748 101532 363754 101544
rect 439314 101532 439320 101544
rect 439372 101532 439378 101584
rect 329098 101396 329104 101448
rect 329156 101436 329162 101448
rect 360838 101436 360844 101448
rect 329156 101408 360844 101436
rect 329156 101396 329162 101408
rect 360838 101396 360844 101408
rect 360896 101396 360902 101448
rect 176102 100784 176108 100836
rect 176160 100824 176166 100836
rect 214006 100824 214012 100836
rect 176160 100796 214012 100824
rect 176160 100784 176166 100796
rect 214006 100784 214012 100796
rect 214064 100784 214070 100836
rect 262766 100784 262772 100836
rect 262824 100824 262830 100836
rect 265158 100824 265164 100836
rect 262824 100796 265164 100824
rect 262824 100784 262830 100796
rect 265158 100784 265164 100796
rect 265216 100784 265222 100836
rect 169294 100716 169300 100768
rect 169352 100756 169358 100768
rect 213914 100756 213920 100768
rect 169352 100728 213920 100756
rect 169352 100716 169358 100728
rect 213914 100716 213920 100728
rect 213972 100716 213978 100768
rect 255958 100716 255964 100768
rect 256016 100756 256022 100768
rect 264974 100756 264980 100768
rect 256016 100728 264980 100756
rect 256016 100716 256022 100728
rect 264974 100716 264980 100728
rect 265032 100716 265038 100768
rect 392578 100716 392584 100768
rect 392636 100756 392642 100768
rect 397454 100756 397460 100768
rect 392636 100728 397460 100756
rect 392636 100716 392642 100728
rect 397454 100716 397460 100728
rect 397512 100716 397518 100768
rect 231670 100648 231676 100700
rect 231728 100688 231734 100700
rect 258810 100688 258816 100700
rect 231728 100660 258816 100688
rect 231728 100648 231734 100660
rect 258810 100648 258816 100660
rect 258868 100648 258874 100700
rect 442902 100648 442908 100700
rect 442960 100688 442966 100700
rect 449158 100688 449164 100700
rect 442960 100660 449164 100688
rect 442960 100648 442966 100660
rect 449158 100648 449164 100660
rect 449216 100648 449222 100700
rect 231762 100580 231768 100632
rect 231820 100620 231826 100632
rect 245286 100620 245292 100632
rect 231820 100592 245292 100620
rect 231820 100580 231826 100592
rect 245286 100580 245292 100592
rect 245344 100580 245350 100632
rect 164970 99968 164976 100020
rect 165028 100008 165034 100020
rect 196802 100008 196808 100020
rect 165028 99980 196808 100008
rect 165028 99968 165034 99980
rect 196802 99968 196808 99980
rect 196860 99968 196866 100020
rect 202874 99968 202880 100020
rect 202932 100008 202938 100020
rect 217226 100008 217232 100020
rect 202932 99980 217232 100008
rect 202932 99968 202938 99980
rect 217226 99968 217232 99980
rect 217284 99968 217290 100020
rect 281994 99968 282000 100020
rect 282052 100008 282058 100020
rect 309226 100008 309232 100020
rect 282052 99980 309232 100008
rect 282052 99968 282058 99980
rect 309226 99968 309232 99980
rect 309284 99968 309290 100020
rect 165062 99832 165068 99884
rect 165120 99872 165126 99884
rect 171870 99872 171876 99884
rect 165120 99844 171876 99872
rect 165120 99832 165126 99844
rect 171870 99832 171876 99844
rect 171928 99832 171934 99884
rect 371970 99424 371976 99476
rect 372028 99464 372034 99476
rect 408402 99464 408408 99476
rect 372028 99436 408408 99464
rect 372028 99424 372034 99436
rect 408402 99424 408408 99436
rect 408460 99424 408466 99476
rect 172054 99356 172060 99408
rect 172112 99396 172118 99408
rect 213914 99396 213920 99408
rect 172112 99368 213920 99396
rect 172112 99356 172118 99368
rect 213914 99356 213920 99368
rect 213972 99356 213978 99408
rect 254670 99356 254676 99408
rect 254728 99396 254734 99408
rect 264974 99396 264980 99408
rect 254728 99368 264980 99396
rect 254728 99356 254734 99368
rect 264974 99356 264980 99368
rect 265032 99356 265038 99408
rect 336090 99356 336096 99408
rect 336148 99396 336154 99408
rect 405826 99396 405832 99408
rect 336148 99368 405832 99396
rect 336148 99356 336154 99368
rect 405826 99356 405832 99368
rect 405884 99356 405890 99408
rect 580166 99396 580172 99408
rect 434640 99368 580172 99396
rect 231670 99288 231676 99340
rect 231728 99328 231734 99340
rect 250714 99328 250720 99340
rect 231728 99300 250720 99328
rect 231728 99288 231734 99300
rect 250714 99288 250720 99300
rect 250772 99288 250778 99340
rect 377490 99288 377496 99340
rect 377548 99328 377554 99340
rect 429010 99328 429016 99340
rect 377548 99300 429016 99328
rect 377548 99288 377554 99300
rect 429010 99288 429016 99300
rect 429068 99288 429074 99340
rect 231762 99220 231768 99272
rect 231820 99260 231826 99272
rect 239490 99260 239496 99272
rect 231820 99232 239496 99260
rect 231820 99220 231826 99232
rect 239490 99220 239496 99232
rect 239548 99220 239554 99272
rect 398650 99220 398656 99272
rect 398708 99260 398714 99272
rect 403250 99260 403256 99272
rect 398708 99232 403256 99260
rect 398708 99220 398714 99232
rect 403250 99220 403256 99232
rect 403308 99220 403314 99272
rect 405826 99220 405832 99272
rect 405884 99260 405890 99272
rect 434640 99260 434668 99368
rect 580166 99356 580172 99368
rect 580224 99356 580230 99408
rect 436830 99288 436836 99340
rect 436888 99328 436894 99340
rect 439498 99328 439504 99340
rect 436888 99300 439504 99328
rect 436888 99288 436894 99300
rect 439498 99288 439504 99300
rect 439556 99288 439562 99340
rect 445754 99328 445760 99340
rect 441586 99300 445760 99328
rect 405884 99232 434668 99260
rect 405884 99220 405890 99232
rect 434162 99152 434168 99204
rect 434220 99192 434226 99204
rect 441586 99192 441614 99300
rect 445754 99288 445760 99300
rect 445812 99288 445818 99340
rect 434220 99164 441614 99192
rect 434220 99152 434226 99164
rect 246298 98608 246304 98660
rect 246356 98648 246362 98660
rect 264514 98648 264520 98660
rect 246356 98620 264520 98648
rect 246356 98608 246362 98620
rect 264514 98608 264520 98620
rect 264572 98608 264578 98660
rect 205174 98064 205180 98116
rect 205232 98104 205238 98116
rect 213914 98104 213920 98116
rect 205232 98076 213920 98104
rect 205232 98064 205238 98076
rect 213914 98064 213920 98076
rect 213972 98064 213978 98116
rect 189810 97996 189816 98048
rect 189868 98036 189874 98048
rect 214006 98036 214012 98048
rect 189868 98008 214012 98036
rect 189868 97996 189874 98008
rect 214006 97996 214012 98008
rect 214064 97996 214070 98048
rect 261662 97996 261668 98048
rect 261720 98036 261726 98048
rect 264974 98036 264980 98048
rect 261720 98008 264980 98036
rect 261720 97996 261726 98008
rect 264974 97996 264980 98008
rect 265032 97996 265038 98048
rect 356698 97928 356704 97980
rect 356756 97968 356762 97980
rect 432874 97968 432880 97980
rect 356756 97940 432880 97968
rect 356756 97928 356762 97940
rect 432874 97928 432880 97940
rect 432932 97928 432938 97980
rect 438026 97928 438032 97980
rect 438084 97968 438090 97980
rect 447134 97968 447140 97980
rect 438084 97940 447140 97968
rect 438084 97928 438090 97940
rect 447134 97928 447140 97940
rect 447192 97928 447198 97980
rect 392762 97860 392768 97912
rect 392820 97900 392826 97912
rect 403894 97900 403900 97912
rect 392820 97872 403900 97900
rect 392820 97860 392826 97872
rect 403894 97860 403900 97872
rect 403952 97860 403958 97912
rect 167822 97248 167828 97300
rect 167880 97288 167886 97300
rect 202230 97288 202236 97300
rect 167880 97260 202236 97288
rect 167880 97248 167886 97260
rect 202230 97248 202236 97260
rect 202288 97248 202294 97300
rect 213454 97248 213460 97300
rect 213512 97288 213518 97300
rect 264974 97288 264980 97300
rect 213512 97260 264980 97288
rect 213512 97248 213518 97260
rect 264974 97248 264980 97260
rect 265032 97248 265038 97300
rect 432690 97180 432696 97232
rect 432748 97220 432754 97232
rect 440418 97220 440424 97232
rect 432748 97192 440424 97220
rect 432748 97180 432754 97192
rect 440418 97180 440424 97192
rect 440476 97180 440482 97232
rect 413278 96908 413284 96960
rect 413336 96948 413342 96960
rect 416130 96948 416136 96960
rect 413336 96920 416136 96948
rect 413336 96908 413342 96920
rect 416130 96908 416136 96920
rect 416188 96908 416194 96960
rect 409046 96840 409052 96892
rect 409104 96880 409110 96892
rect 409966 96880 409972 96892
rect 409104 96852 409972 96880
rect 409104 96840 409110 96852
rect 409966 96840 409972 96852
rect 410024 96840 410030 96892
rect 423214 96840 423220 96892
rect 423272 96880 423278 96892
rect 429286 96880 429292 96892
rect 423272 96852 429292 96880
rect 423272 96840 423278 96852
rect 429286 96840 429292 96852
rect 429344 96840 429350 96892
rect 210418 96704 210424 96756
rect 210476 96744 210482 96756
rect 210476 96716 219204 96744
rect 210476 96704 210482 96716
rect 196802 96636 196808 96688
rect 196860 96676 196866 96688
rect 213914 96676 213920 96688
rect 196860 96648 213920 96676
rect 196860 96636 196866 96648
rect 213914 96636 213920 96648
rect 213972 96636 213978 96688
rect 219176 96076 219204 96716
rect 231670 96636 231676 96688
rect 231728 96676 231734 96688
rect 246482 96676 246488 96688
rect 231728 96648 246488 96676
rect 231728 96636 231734 96648
rect 246482 96636 246488 96648
rect 246540 96636 246546 96688
rect 382918 96568 382924 96620
rect 382976 96608 382982 96620
rect 419994 96608 420000 96620
rect 382976 96580 420000 96608
rect 382976 96568 382982 96580
rect 419994 96568 420000 96580
rect 420052 96568 420058 96620
rect 412910 96364 412916 96416
rect 412968 96404 412974 96416
rect 413370 96404 413376 96416
rect 412968 96376 413376 96404
rect 412968 96364 412974 96376
rect 413370 96364 413376 96376
rect 413428 96364 413434 96416
rect 219158 96024 219164 96076
rect 219216 96024 219222 96076
rect 230474 96024 230480 96076
rect 230532 96064 230538 96076
rect 232590 96064 232596 96076
rect 230532 96036 232596 96064
rect 230532 96024 230538 96036
rect 232590 96024 232596 96036
rect 232648 96024 232654 96076
rect 213178 95956 213184 96008
rect 213236 95996 213242 96008
rect 225598 95996 225604 96008
rect 213236 95968 225604 95996
rect 213236 95956 213242 95968
rect 225598 95956 225604 95968
rect 225656 95956 225662 96008
rect 178862 95888 178868 95940
rect 178920 95928 178926 95940
rect 214650 95928 214656 95940
rect 178920 95900 214656 95928
rect 178920 95888 178926 95900
rect 214650 95888 214656 95900
rect 214708 95888 214714 95940
rect 227070 95888 227076 95940
rect 227128 95928 227134 95940
rect 262766 95928 262772 95940
rect 227128 95900 262772 95928
rect 227128 95888 227134 95900
rect 262766 95888 262772 95900
rect 262824 95888 262830 95940
rect 432598 95820 432604 95872
rect 432656 95860 432662 95872
rect 439130 95860 439136 95872
rect 432656 95832 439136 95860
rect 432656 95820 432662 95832
rect 439130 95820 439136 95832
rect 439188 95820 439194 95872
rect 401318 95208 401324 95260
rect 401376 95248 401382 95260
rect 402974 95248 402980 95260
rect 401376 95220 402980 95248
rect 401376 95208 401382 95220
rect 402974 95208 402980 95220
rect 403032 95208 403038 95260
rect 413370 95208 413376 95260
rect 413428 95248 413434 95260
rect 582742 95248 582748 95260
rect 413428 95220 582748 95248
rect 413428 95208 413434 95220
rect 582742 95208 582748 95220
rect 582800 95208 582806 95260
rect 259362 95140 259368 95192
rect 259420 95180 259426 95192
rect 279418 95180 279424 95192
rect 259420 95152 279424 95180
rect 259420 95140 259426 95152
rect 279418 95140 279424 95152
rect 279476 95140 279482 95192
rect 353938 95140 353944 95192
rect 353996 95180 354002 95192
rect 429654 95180 429660 95192
rect 353996 95152 429660 95180
rect 353996 95140 354002 95152
rect 429654 95140 429660 95152
rect 429712 95140 429718 95192
rect 267826 95072 267832 95124
rect 267884 95112 267890 95124
rect 269114 95112 269120 95124
rect 267884 95084 269120 95112
rect 267884 95072 267890 95084
rect 269114 95072 269120 95084
rect 269172 95072 269178 95124
rect 366910 95072 366916 95124
rect 366968 95112 366974 95124
rect 412266 95112 412272 95124
rect 366968 95084 412272 95112
rect 366968 95072 366974 95084
rect 412266 95072 412272 95084
rect 412324 95072 412330 95124
rect 216214 94528 216220 94580
rect 216272 94568 216278 94580
rect 232774 94568 232780 94580
rect 216272 94540 232780 94568
rect 216272 94528 216278 94540
rect 232774 94528 232780 94540
rect 232832 94528 232838 94580
rect 66070 94460 66076 94512
rect 66128 94500 66134 94512
rect 111150 94500 111156 94512
rect 66128 94472 111156 94500
rect 66128 94460 66134 94472
rect 111150 94460 111156 94472
rect 111208 94460 111214 94512
rect 176194 94460 176200 94512
rect 176252 94500 176258 94512
rect 202414 94500 202420 94512
rect 176252 94472 202420 94500
rect 176252 94460 176258 94472
rect 202414 94460 202420 94472
rect 202472 94460 202478 94512
rect 216674 94460 216680 94512
rect 216732 94500 216738 94512
rect 223482 94500 223488 94512
rect 216732 94472 223488 94500
rect 216732 94460 216738 94472
rect 223482 94460 223488 94472
rect 223540 94460 223546 94512
rect 226978 94460 226984 94512
rect 227036 94500 227042 94512
rect 247954 94500 247960 94512
rect 227036 94472 247960 94500
rect 227036 94460 227042 94472
rect 247954 94460 247960 94472
rect 248012 94460 248018 94512
rect 120626 93916 120632 93968
rect 120684 93956 120690 93968
rect 176010 93956 176016 93968
rect 120684 93928 176016 93956
rect 120684 93916 120690 93928
rect 176010 93916 176016 93928
rect 176068 93916 176074 93968
rect 100662 93848 100668 93900
rect 100720 93888 100726 93900
rect 166534 93888 166540 93900
rect 100720 93860 166540 93888
rect 100720 93848 100726 93860
rect 166534 93848 166540 93860
rect 166592 93848 166598 93900
rect 421282 93848 421288 93900
rect 421340 93888 421346 93900
rect 582834 93888 582840 93900
rect 421340 93860 582840 93888
rect 421340 93848 421346 93860
rect 582834 93848 582840 93860
rect 582892 93848 582898 93900
rect 267734 93780 267740 93832
rect 267792 93820 267798 93832
rect 273990 93820 273996 93832
rect 267792 93792 273996 93820
rect 267792 93780 267798 93792
rect 273990 93780 273996 93792
rect 274048 93780 274054 93832
rect 322198 93780 322204 93832
rect 322256 93820 322262 93832
rect 426434 93820 426440 93832
rect 322256 93792 426440 93820
rect 322256 93780 322262 93792
rect 426434 93780 426440 93792
rect 426492 93780 426498 93832
rect 381722 93712 381728 93764
rect 381780 93752 381786 93764
rect 424502 93752 424508 93764
rect 381780 93724 424508 93752
rect 381780 93712 381786 93724
rect 424502 93712 424508 93724
rect 424560 93712 424566 93764
rect 67358 93168 67364 93220
rect 67416 93208 67422 93220
rect 97258 93208 97264 93220
rect 67416 93180 97264 93208
rect 67416 93168 67422 93180
rect 97258 93168 97264 93180
rect 97316 93168 97322 93220
rect 124122 93168 124128 93220
rect 124180 93208 124186 93220
rect 166258 93208 166264 93220
rect 124180 93180 166264 93208
rect 124180 93168 124186 93180
rect 166258 93168 166264 93180
rect 166316 93168 166322 93220
rect 216030 93168 216036 93220
rect 216088 93208 216094 93220
rect 243446 93208 243452 93220
rect 216088 93180 243452 93208
rect 216088 93168 216094 93180
rect 243446 93168 243452 93180
rect 243504 93168 243510 93220
rect 262122 93168 262128 93220
rect 262180 93208 262186 93220
rect 270586 93208 270592 93220
rect 262180 93180 270592 93208
rect 262180 93168 262186 93180
rect 270586 93168 270592 93180
rect 270644 93168 270650 93220
rect 64782 93100 64788 93152
rect 64840 93140 64846 93152
rect 98638 93140 98644 93152
rect 64840 93112 98644 93140
rect 64840 93100 64846 93112
rect 98638 93100 98644 93112
rect 98696 93100 98702 93152
rect 118234 93100 118240 93152
rect 118292 93140 118298 93152
rect 180334 93140 180340 93152
rect 118292 93112 180340 93140
rect 118292 93100 118298 93112
rect 180334 93100 180340 93112
rect 180392 93100 180398 93152
rect 220078 93100 220084 93152
rect 220136 93140 220142 93152
rect 265894 93140 265900 93152
rect 220136 93112 265900 93140
rect 220136 93100 220142 93112
rect 265894 93100 265900 93112
rect 265952 93100 265958 93152
rect 108114 92488 108120 92540
rect 108172 92528 108178 92540
rect 122098 92528 122104 92540
rect 108172 92500 122104 92528
rect 108172 92488 108178 92500
rect 122098 92488 122104 92500
rect 122156 92488 122162 92540
rect 258810 92488 258816 92540
rect 258868 92528 258874 92540
rect 260374 92528 260380 92540
rect 258868 92500 260380 92528
rect 258868 92488 258874 92500
rect 260374 92488 260380 92500
rect 260432 92488 260438 92540
rect 125778 92420 125784 92472
rect 125836 92460 125842 92472
rect 173250 92460 173256 92472
rect 125836 92432 173256 92460
rect 125836 92420 125842 92432
rect 173250 92420 173256 92432
rect 173308 92420 173314 92472
rect 217226 92420 217232 92472
rect 217284 92460 217290 92472
rect 280430 92460 280436 92472
rect 217284 92432 280436 92460
rect 217284 92420 217290 92432
rect 280430 92420 280436 92432
rect 280488 92420 280494 92472
rect 373258 92420 373264 92472
rect 373316 92460 373322 92472
rect 432230 92460 432236 92472
rect 373316 92432 432236 92460
rect 373316 92420 373322 92432
rect 432230 92420 432236 92432
rect 432288 92420 432294 92472
rect 110138 92352 110144 92404
rect 110196 92392 110202 92404
rect 112438 92392 112444 92404
rect 110196 92364 112444 92392
rect 110196 92352 110202 92364
rect 112438 92352 112444 92364
rect 112496 92352 112502 92404
rect 133138 92352 133144 92404
rect 133196 92392 133202 92404
rect 169110 92392 169116 92404
rect 133196 92364 169116 92392
rect 133196 92352 133202 92364
rect 169110 92352 169116 92364
rect 169168 92352 169174 92404
rect 171870 91808 171876 91860
rect 171928 91848 171934 91860
rect 187142 91848 187148 91860
rect 171928 91820 187148 91848
rect 171928 91808 171934 91820
rect 187142 91808 187148 91820
rect 187200 91808 187206 91860
rect 213178 91808 213184 91860
rect 213236 91848 213242 91860
rect 236914 91848 236920 91860
rect 213236 91820 236920 91848
rect 213236 91808 213242 91820
rect 236914 91808 236920 91820
rect 236972 91808 236978 91860
rect 60642 91740 60648 91792
rect 60700 91780 60706 91792
rect 100018 91780 100024 91792
rect 60700 91752 100024 91780
rect 60700 91740 60706 91752
rect 100018 91740 100024 91752
rect 100076 91740 100082 91792
rect 178034 91740 178040 91792
rect 178092 91780 178098 91792
rect 213362 91780 213368 91792
rect 178092 91752 213368 91780
rect 178092 91740 178098 91752
rect 213362 91740 213368 91752
rect 213420 91740 213426 91792
rect 398742 91740 398748 91792
rect 398800 91780 398806 91792
rect 583018 91780 583024 91792
rect 398800 91752 583024 91780
rect 398800 91740 398806 91752
rect 583018 91740 583024 91752
rect 583076 91740 583082 91792
rect 103422 91128 103428 91180
rect 103480 91168 103486 91180
rect 108298 91168 108304 91180
rect 103480 91140 108304 91168
rect 103480 91128 103486 91140
rect 108298 91128 108304 91140
rect 108356 91128 108362 91180
rect 85114 91060 85120 91112
rect 85172 91100 85178 91112
rect 105538 91100 105544 91112
rect 85172 91072 105544 91100
rect 85172 91060 85178 91072
rect 105538 91060 105544 91072
rect 105596 91060 105602 91112
rect 111242 91060 111248 91112
rect 111300 91100 111306 91112
rect 115290 91100 115296 91112
rect 111300 91072 115296 91100
rect 111300 91060 111306 91072
rect 115290 91060 115296 91072
rect 115348 91060 115354 91112
rect 116762 91060 116768 91112
rect 116820 91100 116826 91112
rect 132862 91100 132868 91112
rect 116820 91072 132868 91100
rect 116820 91060 116826 91072
rect 132862 91060 132868 91072
rect 132920 91060 132926 91112
rect 115750 90992 115756 91044
rect 115808 91032 115814 91044
rect 174630 91032 174636 91044
rect 115808 91004 174636 91032
rect 115808 90992 115814 91004
rect 174630 90992 174636 91004
rect 174688 90992 174694 91044
rect 223482 90992 223488 91044
rect 223540 91032 223546 91044
rect 280338 91032 280344 91044
rect 223540 91004 280344 91032
rect 223540 90992 223546 91004
rect 280338 90992 280344 91004
rect 280396 90992 280402 91044
rect 243446 90924 243452 90976
rect 243504 90964 243510 90976
rect 281718 90964 281724 90976
rect 243504 90936 281724 90964
rect 243504 90924 243510 90936
rect 281718 90924 281724 90936
rect 281776 90924 281782 90976
rect 185578 90380 185584 90432
rect 185636 90420 185642 90432
rect 213454 90420 213460 90432
rect 185636 90392 213460 90420
rect 185636 90380 185642 90392
rect 213454 90380 213460 90392
rect 213512 90380 213518 90432
rect 218698 90380 218704 90432
rect 218756 90420 218762 90432
rect 239674 90420 239680 90432
rect 218756 90392 239680 90420
rect 218756 90380 218762 90392
rect 239674 90380 239680 90392
rect 239732 90380 239738 90432
rect 67542 90312 67548 90364
rect 67600 90352 67606 90364
rect 115198 90352 115204 90364
rect 67600 90324 115204 90352
rect 67600 90312 67606 90324
rect 115198 90312 115204 90324
rect 115256 90312 115262 90364
rect 193858 90312 193864 90364
rect 193916 90352 193922 90364
rect 223022 90352 223028 90364
rect 193916 90324 223028 90352
rect 193916 90312 193922 90324
rect 223022 90312 223028 90324
rect 223080 90312 223086 90364
rect 119890 89632 119896 89684
rect 119948 89672 119954 89684
rect 171778 89672 171784 89684
rect 119948 89644 171784 89672
rect 119948 89632 119954 89644
rect 171778 89632 171784 89644
rect 171836 89632 171842 89684
rect 360838 89632 360844 89684
rect 360896 89672 360902 89684
rect 430298 89672 430304 89684
rect 360896 89644 430304 89672
rect 360896 89632 360902 89644
rect 430298 89632 430304 89644
rect 430356 89632 430362 89684
rect 151630 89564 151636 89616
rect 151688 89604 151694 89616
rect 167822 89604 167828 89616
rect 151688 89576 167828 89604
rect 151688 89564 151694 89576
rect 167822 89564 167828 89576
rect 167880 89564 167886 89616
rect 168374 89564 168380 89616
rect 168432 89604 168438 89616
rect 206370 89604 206376 89616
rect 168432 89576 206376 89604
rect 168432 89564 168438 89576
rect 206370 89564 206376 89576
rect 206428 89564 206434 89616
rect 224218 89020 224224 89072
rect 224276 89060 224282 89072
rect 242434 89060 242440 89072
rect 224276 89032 242440 89060
rect 224276 89020 224282 89032
rect 242434 89020 242440 89032
rect 242492 89020 242498 89072
rect 64690 88952 64696 89004
rect 64748 88992 64754 89004
rect 111058 88992 111064 89004
rect 64748 88964 111064 88992
rect 64748 88952 64754 88964
rect 111058 88952 111064 88964
rect 111116 88952 111122 89004
rect 192662 88952 192668 89004
rect 192720 88992 192726 89004
rect 216122 88992 216128 89004
rect 192720 88964 216128 88992
rect 192720 88952 192726 88964
rect 216122 88952 216128 88964
rect 216180 88952 216186 89004
rect 221458 88952 221464 89004
rect 221516 88992 221522 89004
rect 250806 88992 250812 89004
rect 221516 88964 250812 88992
rect 221516 88952 221522 88964
rect 250806 88952 250812 88964
rect 250864 88952 250870 89004
rect 122282 88272 122288 88324
rect 122340 88312 122346 88324
rect 196710 88312 196716 88324
rect 122340 88284 196716 88312
rect 122340 88272 122346 88284
rect 196710 88272 196716 88284
rect 196768 88272 196774 88324
rect 276014 88272 276020 88324
rect 276072 88312 276078 88324
rect 443362 88312 443368 88324
rect 276072 88284 443368 88312
rect 276072 88272 276078 88284
rect 443362 88272 443368 88284
rect 443420 88272 443426 88324
rect 109218 88204 109224 88256
rect 109276 88244 109282 88256
rect 170582 88244 170588 88256
rect 109276 88216 170588 88244
rect 109276 88204 109282 88216
rect 170582 88204 170588 88216
rect 170640 88204 170646 88256
rect 216306 88204 216312 88256
rect 216364 88244 216370 88256
rect 280522 88244 280528 88256
rect 216364 88216 280528 88244
rect 216364 88204 216370 88216
rect 280522 88204 280528 88216
rect 280580 88204 280586 88256
rect 366358 88204 366364 88256
rect 366416 88244 366422 88256
rect 425146 88244 425152 88256
rect 366416 88216 425152 88244
rect 366416 88204 366422 88216
rect 425146 88204 425152 88216
rect 425204 88204 425210 88256
rect 178954 87660 178960 87712
rect 179012 87700 179018 87712
rect 214834 87700 214840 87712
rect 179012 87672 214840 87700
rect 179012 87660 179018 87672
rect 214834 87660 214840 87672
rect 214892 87660 214898 87712
rect 75270 87592 75276 87644
rect 75328 87632 75334 87644
rect 112530 87632 112536 87644
rect 75328 87604 112536 87632
rect 75328 87592 75334 87604
rect 112530 87592 112536 87604
rect 112588 87592 112594 87644
rect 204898 87592 204904 87644
rect 204956 87632 204962 87644
rect 253474 87632 253480 87644
rect 204956 87604 253480 87632
rect 204956 87592 204962 87604
rect 253474 87592 253480 87604
rect 253532 87592 253538 87644
rect 88058 86912 88064 86964
rect 88116 86952 88122 86964
rect 172054 86952 172060 86964
rect 88116 86924 172060 86952
rect 88116 86912 88122 86924
rect 172054 86912 172060 86924
rect 172112 86912 172118 86964
rect 246482 86912 246488 86964
rect 246540 86952 246546 86964
rect 305638 86952 305644 86964
rect 246540 86924 305644 86952
rect 246540 86912 246546 86924
rect 305638 86912 305644 86924
rect 305696 86952 305702 86964
rect 432690 86952 432696 86964
rect 305696 86924 432696 86952
rect 305696 86912 305702 86924
rect 432690 86912 432696 86924
rect 432748 86912 432754 86964
rect 114370 86844 114376 86896
rect 114428 86884 114434 86896
rect 192570 86884 192576 86896
rect 114428 86856 192576 86884
rect 114428 86844 114434 86856
rect 192570 86844 192576 86856
rect 192628 86844 192634 86896
rect 225598 86844 225604 86896
rect 225656 86884 225662 86896
rect 281626 86884 281632 86896
rect 225656 86856 281632 86884
rect 225656 86844 225662 86856
rect 281626 86844 281632 86856
rect 281684 86844 281690 86896
rect 195238 86232 195244 86284
rect 195296 86272 195302 86284
rect 222838 86272 222844 86284
rect 195296 86244 222844 86272
rect 195296 86232 195302 86244
rect 222838 86232 222844 86244
rect 222896 86232 222902 86284
rect 299658 86232 299664 86284
rect 299716 86272 299722 86284
rect 444466 86272 444472 86284
rect 299716 86244 444472 86272
rect 299716 86232 299722 86244
rect 444466 86232 444472 86244
rect 444524 86232 444530 86284
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 17218 85524 17224 85536
rect 3568 85496 17224 85524
rect 3568 85484 3574 85496
rect 17218 85484 17224 85496
rect 17276 85484 17282 85536
rect 108666 85484 108672 85536
rect 108724 85524 108730 85536
rect 188430 85524 188436 85536
rect 108724 85496 188436 85524
rect 108724 85484 108730 85496
rect 188430 85484 188436 85496
rect 188488 85484 188494 85536
rect 214558 85484 214564 85536
rect 214616 85524 214622 85536
rect 413370 85524 413376 85536
rect 214616 85496 413376 85524
rect 214616 85484 214622 85496
rect 413370 85484 413376 85496
rect 413428 85484 413434 85536
rect 151722 85416 151728 85468
rect 151780 85456 151786 85468
rect 171962 85456 171968 85468
rect 151780 85428 171968 85456
rect 151780 85416 151786 85428
rect 171962 85416 171968 85428
rect 172020 85416 172026 85468
rect 177390 84804 177396 84856
rect 177448 84844 177454 84856
rect 243722 84844 243728 84856
rect 177448 84816 243728 84844
rect 177448 84804 177454 84816
rect 243722 84804 243728 84816
rect 243780 84804 243786 84856
rect 97902 84124 97908 84176
rect 97960 84164 97966 84176
rect 177666 84164 177672 84176
rect 97960 84136 177672 84164
rect 97960 84124 97966 84136
rect 177666 84124 177672 84136
rect 177724 84124 177730 84176
rect 126790 84056 126796 84108
rect 126848 84096 126854 84108
rect 164878 84096 164884 84108
rect 126848 84068 164884 84096
rect 126848 84056 126854 84068
rect 164878 84056 164884 84068
rect 164936 84056 164942 84108
rect 207658 83444 207664 83496
rect 207716 83484 207722 83496
rect 220170 83484 220176 83496
rect 207716 83456 220176 83484
rect 207716 83444 207722 83456
rect 220170 83444 220176 83456
rect 220228 83444 220234 83496
rect 222930 83444 222936 83496
rect 222988 83484 222994 83496
rect 238202 83484 238208 83496
rect 222988 83456 238208 83484
rect 222988 83444 222994 83456
rect 238202 83444 238208 83456
rect 238260 83444 238266 83496
rect 324958 83444 324964 83496
rect 325016 83484 325022 83496
rect 440326 83484 440332 83496
rect 325016 83456 440332 83484
rect 325016 83444 325022 83456
rect 440326 83444 440332 83456
rect 440384 83444 440390 83496
rect 86770 82764 86776 82816
rect 86828 82804 86834 82816
rect 189810 82804 189816 82816
rect 86828 82776 189816 82804
rect 86828 82764 86834 82776
rect 189810 82764 189816 82776
rect 189868 82764 189874 82816
rect 294598 82764 294604 82816
rect 294656 82804 294662 82816
rect 432598 82804 432604 82816
rect 294656 82776 432604 82804
rect 294656 82764 294662 82776
rect 432598 82764 432604 82776
rect 432656 82764 432662 82816
rect 153102 82696 153108 82748
rect 153160 82736 153166 82748
rect 178770 82736 178776 82748
rect 153160 82708 178776 82736
rect 153160 82696 153166 82708
rect 178770 82696 178776 82708
rect 178828 82696 178834 82748
rect 217318 82152 217324 82204
rect 217376 82192 217382 82204
rect 239582 82192 239588 82204
rect 217376 82164 239588 82192
rect 217376 82152 217382 82164
rect 239582 82152 239588 82164
rect 239640 82152 239646 82204
rect 67450 82084 67456 82136
rect 67508 82124 67514 82136
rect 123478 82124 123484 82136
rect 67508 82096 123484 82124
rect 67508 82084 67514 82096
rect 123478 82084 123484 82096
rect 123536 82084 123542 82136
rect 206278 82084 206284 82136
rect 206336 82124 206342 82136
rect 258810 82124 258816 82136
rect 206336 82096 258816 82124
rect 206336 82084 206342 82096
rect 258810 82084 258816 82096
rect 258868 82084 258874 82136
rect 343542 82084 343548 82136
rect 343600 82124 343606 82136
rect 404354 82124 404360 82136
rect 343600 82096 404360 82124
rect 343600 82084 343606 82096
rect 404354 82084 404360 82096
rect 404412 82084 404418 82136
rect 113082 81336 113088 81388
rect 113140 81376 113146 81388
rect 184382 81376 184388 81388
rect 113140 81348 184388 81376
rect 113140 81336 113146 81348
rect 184382 81336 184388 81348
rect 184440 81336 184446 81388
rect 135162 81268 135168 81320
rect 135220 81308 135226 81320
rect 160738 81308 160744 81320
rect 135220 81280 160744 81308
rect 135220 81268 135226 81280
rect 160738 81268 160744 81280
rect 160796 81268 160802 81320
rect 214650 80724 214656 80776
rect 214708 80764 214714 80776
rect 247770 80764 247776 80776
rect 214708 80736 247776 80764
rect 214708 80724 214714 80736
rect 247770 80724 247776 80736
rect 247828 80724 247834 80776
rect 195238 80656 195244 80708
rect 195296 80696 195302 80708
rect 235534 80696 235540 80708
rect 195296 80668 235540 80696
rect 195296 80656 195302 80668
rect 235534 80656 235540 80668
rect 235592 80656 235598 80708
rect 304258 80656 304264 80708
rect 304316 80696 304322 80708
rect 360930 80696 360936 80708
rect 304316 80668 360936 80696
rect 304316 80656 304322 80668
rect 360930 80656 360936 80668
rect 360988 80656 360994 80708
rect 111150 79976 111156 80028
rect 111208 80016 111214 80028
rect 176102 80016 176108 80028
rect 111208 79988 176108 80016
rect 111208 79976 111214 79988
rect 176102 79976 176108 79988
rect 176160 79976 176166 80028
rect 331214 79976 331220 80028
rect 331272 80016 331278 80028
rect 331858 80016 331864 80028
rect 331272 79988 331864 80016
rect 331272 79976 331278 79988
rect 331858 79976 331864 79988
rect 331916 80016 331922 80028
rect 436738 80016 436744 80028
rect 331916 79988 436744 80016
rect 331916 79976 331922 79988
rect 436738 79976 436744 79988
rect 436796 79976 436802 80028
rect 107562 79908 107568 79960
rect 107620 79948 107626 79960
rect 169202 79948 169208 79960
rect 107620 79920 169208 79948
rect 107620 79908 107626 79920
rect 169202 79908 169208 79920
rect 169260 79908 169266 79960
rect 214558 79296 214564 79348
rect 214616 79336 214622 79348
rect 254762 79336 254768 79348
rect 214616 79308 254768 79336
rect 214616 79296 214622 79308
rect 254762 79296 254768 79308
rect 254820 79296 254826 79348
rect 101950 78616 101956 78668
rect 102008 78656 102014 78668
rect 173434 78656 173440 78668
rect 102008 78628 173440 78656
rect 102008 78616 102014 78628
rect 173434 78616 173440 78628
rect 173492 78616 173498 78668
rect 108942 77936 108948 77988
rect 109000 77976 109006 77988
rect 238294 77976 238300 77988
rect 109000 77948 238300 77976
rect 109000 77936 109006 77948
rect 238294 77936 238300 77948
rect 238352 77936 238358 77988
rect 125410 77188 125416 77240
rect 125468 77228 125474 77240
rect 176194 77228 176200 77240
rect 125468 77200 176200 77228
rect 125468 77188 125474 77200
rect 176194 77188 176200 77200
rect 176252 77188 176258 77240
rect 122098 77120 122104 77172
rect 122156 77160 122162 77172
rect 164970 77160 164976 77172
rect 122156 77132 164976 77160
rect 122156 77120 122162 77132
rect 164970 77120 164976 77132
rect 165028 77120 165034 77172
rect 332594 76508 332600 76560
rect 332652 76548 332658 76560
rect 393406 76548 393412 76560
rect 332652 76520 393412 76548
rect 332652 76508 332658 76520
rect 393406 76508 393412 76520
rect 393464 76508 393470 76560
rect 98638 75828 98644 75880
rect 98696 75868 98702 75880
rect 214742 75868 214748 75880
rect 98696 75840 214748 75868
rect 98696 75828 98702 75840
rect 214742 75828 214748 75840
rect 214800 75828 214806 75880
rect 244918 75828 244924 75880
rect 244976 75868 244982 75880
rect 247034 75868 247040 75880
rect 244976 75840 247040 75868
rect 244976 75828 244982 75840
rect 247034 75828 247040 75840
rect 247092 75868 247098 75880
rect 439222 75868 439228 75880
rect 247092 75840 439228 75868
rect 247092 75828 247098 75840
rect 439222 75828 439228 75840
rect 439280 75828 439286 75880
rect 115290 75760 115296 75812
rect 115348 75800 115354 75812
rect 177574 75800 177580 75812
rect 115348 75772 177580 75800
rect 115348 75760 115354 75772
rect 177574 75760 177580 75772
rect 177632 75760 177638 75812
rect 67634 74468 67640 74520
rect 67692 74508 67698 74520
rect 174722 74508 174728 74520
rect 67692 74480 174728 74508
rect 67692 74468 67698 74480
rect 174722 74468 174728 74480
rect 174780 74468 174786 74520
rect 100662 74400 100668 74452
rect 100720 74440 100726 74452
rect 170490 74440 170496 74452
rect 100720 74412 170496 74440
rect 100720 74400 100726 74412
rect 170490 74400 170496 74412
rect 170548 74400 170554 74452
rect 335354 73788 335360 73840
rect 335412 73828 335418 73840
rect 441706 73828 441712 73840
rect 335412 73800 441712 73828
rect 335412 73788 335418 73800
rect 441706 73788 441712 73800
rect 441764 73788 441770 73840
rect 107562 72496 107568 72548
rect 107620 72536 107626 72548
rect 229738 72536 229744 72548
rect 107620 72508 229744 72536
rect 107620 72496 107626 72508
rect 229738 72496 229744 72508
rect 229796 72496 229802 72548
rect 122742 72428 122748 72480
rect 122800 72468 122806 72480
rect 261570 72468 261576 72480
rect 122800 72440 261576 72468
rect 122800 72428 122806 72440
rect 261570 72428 261576 72440
rect 261628 72428 261634 72480
rect 344278 72428 344284 72480
rect 344336 72468 344342 72480
rect 414198 72468 414204 72480
rect 344336 72440 414204 72468
rect 344336 72428 344342 72440
rect 414198 72428 414204 72440
rect 414256 72428 414262 72480
rect 100018 71680 100024 71732
rect 100076 71720 100082 71732
rect 202322 71720 202328 71732
rect 100076 71692 202328 71720
rect 100076 71680 100082 71692
rect 202322 71680 202328 71692
rect 202380 71680 202386 71732
rect 126882 71612 126888 71664
rect 126940 71652 126946 71664
rect 173158 71652 173164 71664
rect 126940 71624 173164 71652
rect 126940 71612 126946 71624
rect 173158 71612 173164 71624
rect 173216 71612 173222 71664
rect 99190 70320 99196 70372
rect 99248 70360 99254 70372
rect 171870 70360 171876 70372
rect 99248 70332 171876 70360
rect 99248 70320 99254 70332
rect 171870 70320 171876 70332
rect 171928 70320 171934 70372
rect 48130 69640 48136 69692
rect 48188 69680 48194 69692
rect 249242 69680 249248 69692
rect 48188 69652 249248 69680
rect 48188 69640 48194 69652
rect 249242 69640 249248 69652
rect 249300 69640 249306 69692
rect 336734 69640 336740 69692
rect 336792 69680 336798 69692
rect 440234 69680 440240 69692
rect 336792 69652 440240 69680
rect 336792 69640 336798 69652
rect 440234 69640 440240 69652
rect 440292 69640 440298 69692
rect 115198 68960 115204 69012
rect 115256 69000 115262 69012
rect 196802 69000 196808 69012
rect 115256 68972 196808 69000
rect 115256 68960 115262 68972
rect 196802 68960 196808 68972
rect 196860 68960 196866 69012
rect 106090 68892 106096 68944
rect 106148 68932 106154 68944
rect 180242 68932 180248 68944
rect 106148 68904 180248 68932
rect 106148 68892 106154 68904
rect 180242 68892 180248 68904
rect 180300 68892 180306 68944
rect 330478 67668 330484 67720
rect 330536 67708 330542 67720
rect 335354 67708 335360 67720
rect 330536 67680 335360 67708
rect 330536 67668 330542 67680
rect 335354 67668 335360 67680
rect 335412 67668 335418 67720
rect 334618 67600 334624 67652
rect 334676 67640 334682 67652
rect 336734 67640 336740 67652
rect 334676 67612 336740 67640
rect 334676 67600 334682 67612
rect 336734 67600 336740 67612
rect 336792 67600 336798 67652
rect 103330 67532 103336 67584
rect 103388 67572 103394 67584
rect 199378 67572 199384 67584
rect 103388 67544 199384 67572
rect 103388 67532 103394 67544
rect 199378 67532 199384 67544
rect 199436 67532 199442 67584
rect 337470 67532 337476 67584
rect 337528 67572 337534 67584
rect 401962 67572 401968 67584
rect 337528 67544 401968 67572
rect 337528 67532 337534 67544
rect 401962 67532 401968 67544
rect 402020 67532 402026 67584
rect 124030 67464 124036 67516
rect 124088 67504 124094 67516
rect 178862 67504 178868 67516
rect 124088 67476 178868 67504
rect 124088 67464 124094 67476
rect 178862 67464 178868 67476
rect 178920 67464 178926 67516
rect 323670 66852 323676 66904
rect 323728 66892 323734 66904
rect 337470 66892 337476 66904
rect 323728 66864 337476 66892
rect 323728 66852 323734 66864
rect 337470 66852 337476 66864
rect 337528 66852 337534 66904
rect 110138 66172 110144 66224
rect 110196 66212 110202 66224
rect 192662 66212 192668 66224
rect 110196 66184 192668 66212
rect 110196 66172 110202 66184
rect 192662 66172 192668 66184
rect 192720 66172 192726 66224
rect 151538 66104 151544 66156
rect 151596 66144 151602 66156
rect 169018 66144 169024 66156
rect 151596 66116 169024 66144
rect 151596 66104 151602 66116
rect 169018 66104 169024 66116
rect 169076 66104 169082 66156
rect 292482 65492 292488 65544
rect 292540 65532 292546 65544
rect 428366 65532 428372 65544
rect 292540 65504 428372 65532
rect 292540 65492 292546 65504
rect 428366 65492 428372 65504
rect 428424 65492 428430 65544
rect 102042 64812 102048 64864
rect 102100 64852 102106 64864
rect 205082 64852 205088 64864
rect 102100 64824 205088 64852
rect 102100 64812 102106 64824
rect 205082 64812 205088 64824
rect 205140 64812 205146 64864
rect 112530 64744 112536 64796
rect 112588 64784 112594 64796
rect 178954 64784 178960 64796
rect 112588 64756 178960 64784
rect 112588 64744 112594 64756
rect 178954 64744 178960 64756
rect 179012 64744 179018 64796
rect 284938 64132 284944 64184
rect 284996 64172 285002 64184
rect 352742 64172 352748 64184
rect 284996 64144 352748 64172
rect 284996 64132 285002 64144
rect 352742 64132 352748 64144
rect 352800 64132 352806 64184
rect 89622 63452 89628 63504
rect 89680 63492 89686 63504
rect 162118 63492 162124 63504
rect 89680 63464 162124 63492
rect 89680 63452 89686 63464
rect 162118 63452 162124 63464
rect 162176 63452 162182 63504
rect 292666 63452 292672 63504
rect 292724 63492 292730 63504
rect 425698 63492 425704 63504
rect 292724 63464 425704 63492
rect 292724 63452 292730 63464
rect 425698 63452 425704 63464
rect 425756 63452 425762 63504
rect 124122 63384 124128 63436
rect 124180 63424 124186 63436
rect 193950 63424 193956 63436
rect 124180 63396 193956 63424
rect 124180 63384 124186 63396
rect 193950 63384 193956 63396
rect 194008 63384 194014 63436
rect 266354 62772 266360 62824
rect 266412 62812 266418 62824
rect 292666 62812 292672 62824
rect 266412 62784 292672 62812
rect 266412 62772 266418 62784
rect 292666 62772 292672 62784
rect 292724 62772 292730 62824
rect 104158 62024 104164 62076
rect 104216 62064 104222 62076
rect 203518 62064 203524 62076
rect 104216 62036 203524 62064
rect 104216 62024 104222 62036
rect 203518 62024 203524 62036
rect 203576 62024 203582 62076
rect 262950 61412 262956 61464
rect 263008 61452 263014 61464
rect 399478 61452 399484 61464
rect 263008 61424 399484 61452
rect 263008 61412 263014 61424
rect 399478 61412 399484 61424
rect 399536 61412 399542 61464
rect 59262 61344 59268 61396
rect 59320 61384 59326 61396
rect 263042 61384 263048 61396
rect 59320 61356 263048 61384
rect 59320 61344 59326 61356
rect 263042 61344 263048 61356
rect 263100 61344 263106 61396
rect 116578 60664 116584 60716
rect 116636 60704 116642 60716
rect 210510 60704 210516 60716
rect 116636 60676 210516 60704
rect 116636 60664 116642 60676
rect 210510 60664 210516 60676
rect 210568 60664 210574 60716
rect 84102 59984 84108 60036
rect 84160 60024 84166 60036
rect 242250 60024 242256 60036
rect 84160 59996 242256 60024
rect 84160 59984 84166 59996
rect 242250 59984 242256 59996
rect 242308 59984 242314 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 40678 59344 40684 59356
rect 3108 59316 40684 59344
rect 3108 59304 3114 59316
rect 40678 59304 40684 59316
rect 40736 59304 40742 59356
rect 108298 59304 108304 59356
rect 108356 59344 108362 59356
rect 209130 59344 209136 59356
rect 108356 59316 209136 59344
rect 108356 59304 108362 59316
rect 209130 59304 209136 59316
rect 209188 59304 209194 59356
rect 311894 59304 311900 59356
rect 311952 59344 311958 59356
rect 407114 59344 407120 59356
rect 311952 59316 407120 59344
rect 311952 59304 311958 59316
rect 407114 59304 407120 59316
rect 407172 59304 407178 59356
rect 115842 58624 115848 58676
rect 115900 58664 115906 58676
rect 247678 58664 247684 58676
rect 115900 58636 247684 58664
rect 115900 58624 115906 58636
rect 247678 58624 247684 58636
rect 247736 58624 247742 58676
rect 248322 58624 248328 58676
rect 248380 58664 248386 58676
rect 311894 58664 311900 58676
rect 248380 58636 311900 58664
rect 248380 58624 248386 58636
rect 311894 58624 311900 58636
rect 311952 58624 311958 58676
rect 107470 57876 107476 57928
rect 107528 57916 107534 57928
rect 211798 57916 211804 57928
rect 107528 57888 211804 57916
rect 107528 57876 107534 57888
rect 211798 57876 211804 57888
rect 211856 57876 211862 57928
rect 220170 57264 220176 57316
rect 220228 57304 220234 57316
rect 259454 57304 259460 57316
rect 220228 57276 259460 57304
rect 220228 57264 220234 57276
rect 259454 57264 259460 57276
rect 259512 57304 259518 57316
rect 342990 57304 342996 57316
rect 259512 57276 342996 57304
rect 259512 57264 259518 57276
rect 342990 57264 342996 57276
rect 343048 57264 343054 57316
rect 104802 57196 104808 57248
rect 104860 57236 104866 57248
rect 260282 57236 260288 57248
rect 104860 57208 260288 57236
rect 104860 57196 104866 57208
rect 260282 57196 260288 57208
rect 260340 57196 260346 57248
rect 346394 57196 346400 57248
rect 346452 57236 346458 57248
rect 446030 57236 446036 57248
rect 346452 57208 446036 57236
rect 346452 57196 346458 57208
rect 446030 57196 446036 57208
rect 446088 57196 446094 57248
rect 123478 56516 123484 56568
rect 123536 56556 123542 56568
rect 213270 56556 213276 56568
rect 123536 56528 213276 56556
rect 123536 56516 123542 56528
rect 213270 56516 213276 56528
rect 213328 56516 213334 56568
rect 91002 55836 91008 55888
rect 91060 55876 91066 55888
rect 264422 55876 264428 55888
rect 91060 55848 264428 55876
rect 91060 55836 91066 55848
rect 264422 55836 264428 55848
rect 264480 55836 264486 55888
rect 112438 55156 112444 55208
rect 112496 55196 112502 55208
rect 198090 55196 198096 55208
rect 112496 55168 198096 55196
rect 112496 55156 112502 55168
rect 198090 55156 198096 55168
rect 198148 55156 198154 55208
rect 382918 54544 382924 54596
rect 382976 54584 382982 54596
rect 422570 54584 422576 54596
rect 382976 54556 422576 54584
rect 382976 54544 382982 54556
rect 422570 54544 422576 54556
rect 422628 54544 422634 54596
rect 89622 54476 89628 54528
rect 89680 54516 89686 54528
rect 243538 54516 243544 54528
rect 89680 54488 243544 54516
rect 89680 54476 89686 54488
rect 243538 54476 243544 54488
rect 243596 54476 243602 54528
rect 335354 54476 335360 54528
rect 335412 54516 335418 54528
rect 383010 54516 383016 54528
rect 335412 54488 383016 54516
rect 335412 54476 335418 54488
rect 383010 54476 383016 54488
rect 383068 54476 383074 54528
rect 340782 53728 340788 53780
rect 340840 53768 340846 53780
rect 435450 53768 435456 53780
rect 340840 53740 435456 53768
rect 340840 53728 340846 53740
rect 435450 53728 435456 53740
rect 435508 53728 435514 53780
rect 340138 53252 340144 53304
rect 340196 53292 340202 53304
rect 340782 53292 340788 53304
rect 340196 53264 340788 53292
rect 340196 53252 340202 53264
rect 340782 53252 340788 53264
rect 340840 53252 340846 53304
rect 146938 53116 146944 53168
rect 146996 53156 147002 53168
rect 227070 53156 227076 53168
rect 146996 53128 227076 53156
rect 146996 53116 147002 53128
rect 227070 53116 227076 53128
rect 227128 53116 227134 53168
rect 41322 53048 41328 53100
rect 41380 53088 41386 53100
rect 231118 53088 231124 53100
rect 41380 53060 231124 53088
rect 41380 53048 41386 53060
rect 231118 53048 231124 53060
rect 231176 53048 231182 53100
rect 117130 52368 117136 52420
rect 117188 52408 117194 52420
rect 191190 52408 191196 52420
rect 117188 52380 191196 52408
rect 117188 52368 117194 52380
rect 191190 52368 191196 52380
rect 191248 52368 191254 52420
rect 250530 51756 250536 51808
rect 250588 51796 250594 51808
rect 416774 51796 416780 51808
rect 250588 51768 416780 51796
rect 250588 51756 250594 51768
rect 416774 51756 416780 51768
rect 416832 51756 416838 51808
rect 17862 51688 17868 51740
rect 17920 51728 17926 51740
rect 254670 51728 254676 51740
rect 17920 51700 254676 51728
rect 17920 51688 17926 51700
rect 254670 51688 254676 51700
rect 254728 51688 254734 51740
rect 106182 51008 106188 51060
rect 106240 51048 106246 51060
rect 195330 51048 195336 51060
rect 106240 51020 195336 51048
rect 106240 51008 106246 51020
rect 195330 51008 195336 51020
rect 195388 51008 195394 51060
rect 136542 50940 136548 50992
rect 136600 50980 136606 50992
rect 180150 50980 180156 50992
rect 136600 50952 180156 50980
rect 136600 50940 136606 50952
rect 180150 50940 180156 50952
rect 180208 50940 180214 50992
rect 52362 50328 52368 50380
rect 52420 50368 52426 50380
rect 135254 50368 135260 50380
rect 52420 50340 135260 50368
rect 52420 50328 52426 50340
rect 135254 50328 135260 50340
rect 135312 50328 135318 50380
rect 186958 50328 186964 50380
rect 187016 50368 187022 50380
rect 302970 50368 302976 50380
rect 187016 50340 302976 50368
rect 187016 50328 187022 50340
rect 302970 50328 302976 50340
rect 303028 50328 303034 50380
rect 321554 50328 321560 50380
rect 321612 50368 321618 50380
rect 408494 50368 408500 50380
rect 321612 50340 408500 50368
rect 321612 50328 321618 50340
rect 408494 50328 408500 50340
rect 408552 50328 408558 50380
rect 86862 49648 86868 49700
rect 86920 49688 86926 49700
rect 205174 49688 205180 49700
rect 86920 49660 205180 49688
rect 86920 49648 86926 49660
rect 205174 49648 205180 49660
rect 205232 49648 205238 49700
rect 114462 48968 114468 49020
rect 114520 49008 114526 49020
rect 236638 49008 236644 49020
rect 114520 48980 236644 49008
rect 114520 48968 114526 48980
rect 236638 48968 236644 48980
rect 236696 48968 236702 49020
rect 297358 48968 297364 49020
rect 297416 49008 297422 49020
rect 444374 49008 444380 49020
rect 297416 48980 444380 49008
rect 297416 48968 297422 48980
rect 444374 48968 444380 48980
rect 444432 48968 444438 49020
rect 129642 48220 129648 48272
rect 129700 48260 129706 48272
rect 192478 48260 192484 48272
rect 129700 48232 192484 48260
rect 129700 48220 129706 48232
rect 192478 48220 192484 48232
rect 192536 48220 192542 48272
rect 227070 47608 227076 47660
rect 227128 47648 227134 47660
rect 269114 47648 269120 47660
rect 227128 47620 269120 47648
rect 227128 47608 227134 47620
rect 269114 47608 269120 47620
rect 269172 47608 269178 47660
rect 133138 47540 133144 47592
rect 133196 47580 133202 47592
rect 217318 47580 217324 47592
rect 133196 47552 217324 47580
rect 133196 47540 133202 47552
rect 217318 47540 217324 47552
rect 217376 47540 217382 47592
rect 268378 47540 268384 47592
rect 268436 47580 268442 47592
rect 454126 47580 454132 47592
rect 268436 47552 454132 47580
rect 268436 47540 268442 47552
rect 454126 47540 454132 47552
rect 454184 47540 454190 47592
rect 300762 46860 300768 46912
rect 300820 46900 300826 46912
rect 400674 46900 400680 46912
rect 300820 46872 400680 46900
rect 300820 46860 300826 46872
rect 400674 46860 400680 46872
rect 400732 46860 400738 46912
rect 85482 46248 85488 46300
rect 85540 46288 85546 46300
rect 266998 46288 267004 46300
rect 85540 46260 267004 46288
rect 85540 46248 85546 46260
rect 266998 46248 267004 46260
rect 267056 46248 267062 46300
rect 71038 46180 71044 46232
rect 71096 46220 71102 46232
rect 258718 46220 258724 46232
rect 71096 46192 258724 46220
rect 71096 46180 71102 46192
rect 258718 46180 258724 46192
rect 258776 46180 258782 46232
rect 269758 46180 269764 46232
rect 269816 46220 269822 46232
rect 299474 46220 299480 46232
rect 269816 46192 299480 46220
rect 269816 46180 269822 46192
rect 299474 46180 299480 46192
rect 299532 46220 299538 46232
rect 300762 46220 300768 46232
rect 299532 46192 300768 46220
rect 299532 46180 299538 46192
rect 300762 46180 300768 46192
rect 300820 46180 300826 46232
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 43438 45540 43444 45552
rect 3568 45512 43444 45540
rect 3568 45500 3574 45512
rect 43438 45500 43444 45512
rect 43496 45500 43502 45552
rect 95050 44820 95056 44872
rect 95108 44860 95114 44872
rect 253198 44860 253204 44872
rect 95108 44832 253204 44860
rect 95108 44820 95114 44832
rect 253198 44820 253204 44832
rect 253256 44820 253262 44872
rect 257338 44820 257344 44872
rect 257396 44860 257402 44872
rect 400858 44860 400864 44872
rect 257396 44832 400864 44860
rect 257396 44820 257402 44832
rect 400858 44820 400864 44832
rect 400916 44820 400922 44872
rect 12250 43392 12256 43444
rect 12308 43432 12314 43444
rect 245010 43432 245016 43444
rect 12308 43404 245016 43432
rect 12308 43392 12314 43404
rect 245010 43392 245016 43404
rect 245068 43392 245074 43444
rect 246390 43392 246396 43444
rect 246448 43432 246454 43444
rect 405734 43432 405740 43444
rect 246448 43404 405740 43432
rect 246448 43392 246454 43404
rect 405734 43392 405740 43404
rect 405792 43392 405798 43444
rect 283558 42712 283564 42764
rect 283616 42752 283622 42764
rect 452746 42752 452752 42764
rect 283616 42724 452752 42752
rect 283616 42712 283622 42724
rect 452746 42712 452752 42724
rect 452804 42712 452810 42764
rect 37182 42100 37188 42152
rect 37240 42140 37246 42152
rect 147030 42140 147036 42152
rect 37240 42112 147036 42140
rect 37240 42100 37246 42112
rect 147030 42100 147036 42112
rect 147088 42100 147094 42152
rect 147122 42100 147128 42152
rect 147180 42140 147186 42152
rect 230474 42140 230480 42152
rect 147180 42112 230480 42140
rect 147180 42100 147186 42112
rect 230474 42100 230480 42112
rect 230532 42100 230538 42152
rect 105538 42032 105544 42084
rect 105596 42072 105602 42084
rect 250438 42072 250444 42084
rect 105596 42044 250444 42072
rect 105596 42032 105602 42044
rect 250438 42032 250444 42044
rect 250496 42032 250502 42084
rect 99282 40740 99288 40792
rect 99340 40780 99346 40792
rect 239398 40780 239404 40792
rect 99340 40752 239404 40780
rect 99340 40740 99346 40752
rect 239398 40740 239404 40752
rect 239456 40740 239462 40792
rect 46842 40672 46848 40724
rect 46900 40712 46906 40724
rect 240870 40712 240876 40724
rect 46900 40684 240876 40712
rect 46900 40672 46906 40684
rect 240870 40672 240876 40684
rect 240928 40672 240934 40724
rect 228358 39312 228364 39364
rect 228416 39352 228422 39364
rect 258074 39352 258080 39364
rect 228416 39324 258080 39352
rect 228416 39312 228422 39324
rect 258074 39312 258080 39324
rect 258132 39352 258138 39364
rect 436094 39352 436100 39364
rect 258132 39324 436100 39352
rect 258132 39312 258138 39324
rect 436094 39312 436100 39324
rect 436152 39312 436158 39364
rect 39942 37884 39948 37936
rect 40000 37924 40006 37936
rect 222930 37924 222936 37936
rect 40000 37896 222936 37924
rect 40000 37884 40006 37896
rect 222930 37884 222936 37896
rect 222988 37884 222994 37936
rect 314654 37884 314660 37936
rect 314712 37924 314718 37936
rect 456886 37924 456892 37936
rect 314712 37896 456892 37924
rect 314712 37884 314718 37896
rect 456886 37884 456892 37896
rect 456944 37884 456950 37936
rect 320818 37204 320824 37256
rect 320876 37244 320882 37256
rect 392578 37244 392584 37256
rect 320876 37216 392584 37244
rect 320876 37204 320882 37216
rect 392578 37204 392584 37216
rect 392636 37204 392642 37256
rect 320174 36864 320180 36916
rect 320232 36904 320238 36916
rect 320818 36904 320824 36916
rect 320232 36876 320824 36904
rect 320232 36864 320238 36876
rect 320818 36864 320824 36876
rect 320876 36864 320882 36916
rect 247034 36660 247040 36712
rect 247092 36700 247098 36712
rect 248322 36700 248328 36712
rect 247092 36672 248328 36700
rect 247092 36660 247098 36672
rect 248322 36660 248328 36672
rect 248380 36660 248386 36712
rect 54478 36524 54484 36576
rect 54536 36564 54542 36576
rect 265710 36564 265716 36576
rect 54536 36536 265716 36564
rect 54536 36524 54542 36536
rect 265710 36524 265716 36536
rect 265768 36524 265774 36576
rect 316770 35844 316776 35896
rect 316828 35884 316834 35896
rect 442994 35884 443000 35896
rect 316828 35856 443000 35884
rect 316828 35844 316834 35856
rect 442994 35844 443000 35856
rect 443052 35844 443058 35896
rect 186958 35232 186964 35284
rect 187016 35272 187022 35284
rect 221458 35272 221464 35284
rect 187016 35244 221464 35272
rect 187016 35232 187022 35244
rect 221458 35232 221464 35244
rect 221516 35232 221522 35284
rect 61930 35164 61936 35216
rect 61988 35204 61994 35216
rect 224310 35204 224316 35216
rect 61988 35176 224316 35204
rect 61988 35164 61994 35176
rect 224310 35164 224316 35176
rect 224368 35164 224374 35216
rect 316034 34484 316040 34536
rect 316092 34524 316098 34536
rect 316770 34524 316776 34536
rect 316092 34496 316776 34524
rect 316092 34484 316098 34496
rect 316770 34484 316776 34496
rect 316828 34484 316834 34536
rect 86862 33804 86868 33856
rect 86920 33844 86926 33856
rect 226978 33844 226984 33856
rect 86920 33816 226984 33844
rect 86920 33804 86926 33816
rect 226978 33804 226984 33816
rect 227036 33804 227042 33856
rect 61378 33736 61384 33788
rect 61436 33776 61442 33788
rect 279418 33776 279424 33788
rect 61436 33748 279424 33776
rect 61436 33736 61442 33748
rect 279418 33736 279424 33748
rect 279476 33736 279482 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 15838 33096 15844 33108
rect 3568 33068 15844 33096
rect 3568 33056 3574 33068
rect 15838 33056 15844 33068
rect 15896 33056 15902 33108
rect 74442 32444 74448 32496
rect 74500 32484 74506 32496
rect 260098 32484 260104 32496
rect 74500 32456 260104 32484
rect 74500 32444 74506 32456
rect 260098 32444 260104 32456
rect 260156 32444 260162 32496
rect 62022 32376 62028 32428
rect 62080 32416 62086 32428
rect 274634 32416 274640 32428
rect 62080 32388 274640 32416
rect 62080 32376 62086 32388
rect 274634 32376 274640 32388
rect 274692 32376 274698 32428
rect 309870 32376 309876 32428
rect 309928 32416 309934 32428
rect 393958 32416 393964 32428
rect 309928 32388 393964 32416
rect 309928 32376 309934 32388
rect 393958 32376 393964 32388
rect 394016 32376 394022 32428
rect 78582 31084 78588 31136
rect 78640 31124 78646 31136
rect 262858 31124 262864 31136
rect 78640 31096 262864 31124
rect 78640 31084 78646 31096
rect 262858 31084 262864 31096
rect 262916 31084 262922 31136
rect 59998 31016 60004 31068
rect 60056 31056 60062 31068
rect 246298 31056 246304 31068
rect 60056 31028 246304 31056
rect 60056 31016 60062 31028
rect 246298 31016 246304 31028
rect 246356 31016 246362 31068
rect 252554 31016 252560 31068
rect 252612 31056 252618 31068
rect 304258 31056 304264 31068
rect 252612 31028 304264 31056
rect 252612 31016 252618 31028
rect 304258 31016 304264 31028
rect 304316 31016 304322 31068
rect 112438 29656 112444 29708
rect 112496 29696 112502 29708
rect 204898 29696 204904 29708
rect 112496 29668 204904 29696
rect 112496 29656 112502 29668
rect 204898 29656 204904 29668
rect 204956 29656 204962 29708
rect 56502 29588 56508 29640
rect 56560 29628 56566 29640
rect 264330 29628 264336 29640
rect 56560 29600 264336 29628
rect 56560 29588 56566 29600
rect 264330 29588 264336 29600
rect 264388 29588 264394 29640
rect 282270 29588 282276 29640
rect 282328 29628 282334 29640
rect 389910 29628 389916 29640
rect 282328 29600 389916 29628
rect 282328 29588 282334 29600
rect 389910 29588 389916 29600
rect 389968 29588 389974 29640
rect 160738 28364 160744 28416
rect 160796 28404 160802 28416
rect 214650 28404 214656 28416
rect 160796 28376 214656 28404
rect 160796 28364 160802 28376
rect 214650 28364 214656 28376
rect 214708 28364 214714 28416
rect 37090 28296 37096 28348
rect 37148 28336 37154 28348
rect 178678 28336 178684 28348
rect 37148 28308 178684 28336
rect 37148 28296 37154 28308
rect 178678 28296 178684 28308
rect 178736 28296 178742 28348
rect 106 28228 112 28280
rect 164 28268 170 28280
rect 147122 28268 147128 28280
rect 164 28240 147128 28268
rect 164 28228 170 28240
rect 147122 28228 147128 28240
rect 147180 28228 147186 28280
rect 188338 28228 188344 28280
rect 188396 28268 188402 28280
rect 270494 28268 270500 28280
rect 188396 28240 270500 28268
rect 188396 28228 188402 28240
rect 270494 28228 270500 28240
rect 270552 28228 270558 28280
rect 277394 28228 277400 28280
rect 277452 28268 277458 28280
rect 294598 28268 294604 28280
rect 277452 28240 294604 28268
rect 277452 28228 277458 28240
rect 294598 28228 294604 28240
rect 294656 28228 294662 28280
rect 303614 28228 303620 28280
rect 303672 28268 303678 28280
rect 327074 28268 327080 28280
rect 303672 28240 327080 28268
rect 303672 28228 303678 28240
rect 327074 28228 327080 28240
rect 327132 28228 327138 28280
rect 274634 27548 274640 27600
rect 274692 27588 274698 27600
rect 417418 27588 417424 27600
rect 274692 27560 417424 27588
rect 274692 27548 274698 27560
rect 417418 27548 417424 27560
rect 417476 27548 417482 27600
rect 81342 26936 81348 26988
rect 81400 26976 81406 26988
rect 232498 26976 232504 26988
rect 81400 26948 232504 26976
rect 81400 26936 81406 26948
rect 232498 26936 232504 26948
rect 232556 26936 232562 26988
rect 16482 26868 16488 26920
rect 16540 26908 16546 26920
rect 185578 26908 185584 26920
rect 16540 26880 185584 26908
rect 16540 26868 16546 26880
rect 185578 26868 185584 26880
rect 185636 26868 185642 26920
rect 270494 26188 270500 26240
rect 270552 26228 270558 26240
rect 371878 26228 371884 26240
rect 270552 26200 371884 26228
rect 270552 26188 270558 26200
rect 371878 26188 371884 26200
rect 371936 26188 371942 26240
rect 200758 25576 200764 25628
rect 200816 25616 200822 25628
rect 268470 25616 268476 25628
rect 200816 25588 268476 25616
rect 200816 25576 200822 25588
rect 268470 25576 268476 25588
rect 268528 25576 268534 25628
rect 125502 25508 125508 25560
rect 125560 25548 125566 25560
rect 216030 25548 216036 25560
rect 125560 25520 216036 25548
rect 125560 25508 125566 25520
rect 216030 25508 216036 25520
rect 216088 25508 216094 25560
rect 327074 24148 327080 24200
rect 327132 24188 327138 24200
rect 419350 24188 419356 24200
rect 327132 24160 419356 24188
rect 327132 24148 327138 24160
rect 419350 24148 419356 24160
rect 419408 24148 419414 24200
rect 100662 24080 100668 24132
rect 100720 24120 100726 24132
rect 235258 24120 235264 24132
rect 100720 24092 235264 24120
rect 100720 24080 100726 24092
rect 235258 24080 235264 24092
rect 235316 24080 235322 24132
rect 264330 24080 264336 24132
rect 264388 24120 264394 24132
rect 374730 24120 374736 24132
rect 264388 24092 374736 24120
rect 264388 24080 264394 24092
rect 374730 24080 374736 24092
rect 374788 24080 374794 24132
rect 67174 22788 67180 22840
rect 67232 22828 67238 22840
rect 255958 22828 255964 22840
rect 67232 22800 255964 22828
rect 67232 22788 67238 22800
rect 255958 22788 255964 22800
rect 256016 22788 256022 22840
rect 259546 22788 259552 22840
rect 259604 22828 259610 22840
rect 395338 22828 395344 22840
rect 259604 22800 395344 22828
rect 259604 22788 259610 22800
rect 395338 22788 395344 22800
rect 395396 22788 395402 22840
rect 20622 22720 20628 22772
rect 20680 22760 20686 22772
rect 261478 22760 261484 22772
rect 20680 22732 261484 22760
rect 20680 22720 20686 22732
rect 261478 22720 261484 22732
rect 261536 22720 261542 22772
rect 111610 21428 111616 21480
rect 111668 21468 111674 21480
rect 238018 21468 238024 21480
rect 111668 21440 238024 21468
rect 111668 21428 111674 21440
rect 238018 21428 238024 21440
rect 238076 21428 238082 21480
rect 57882 21360 57888 21412
rect 57940 21400 57946 21412
rect 251910 21400 251916 21412
rect 57940 21372 251916 21400
rect 57940 21360 57946 21372
rect 251910 21360 251916 21372
rect 251968 21360 251974 21412
rect 257430 21360 257436 21412
rect 257488 21400 257494 21412
rect 447226 21400 447232 21412
rect 257488 21372 447232 21400
rect 257488 21360 257494 21372
rect 447226 21360 447232 21372
rect 447284 21360 447290 21412
rect 334710 20612 334716 20664
rect 334768 20652 334774 20664
rect 335262 20652 335268 20664
rect 334768 20624 335268 20652
rect 334768 20612 334774 20624
rect 335262 20612 335268 20624
rect 335320 20652 335326 20664
rect 429286 20652 429292 20664
rect 335320 20624 429292 20652
rect 335320 20612 335326 20624
rect 429286 20612 429292 20624
rect 429344 20612 429350 20664
rect 45462 20000 45468 20052
rect 45520 20040 45526 20052
rect 133138 20040 133144 20052
rect 45520 20012 133144 20040
rect 45520 20000 45526 20012
rect 133138 20000 133144 20012
rect 133196 20000 133202 20052
rect 189718 20000 189724 20052
rect 189776 20040 189782 20052
rect 215938 20040 215944 20052
rect 189776 20012 215944 20040
rect 189776 20000 189782 20012
rect 215938 20000 215944 20012
rect 215996 20000 216002 20052
rect 88242 19932 88248 19984
rect 88300 19972 88306 19984
rect 249058 19972 249064 19984
rect 88300 19944 249064 19972
rect 88300 19932 88306 19944
rect 249058 19932 249064 19944
rect 249116 19932 249122 19984
rect 250438 19932 250444 19984
rect 250496 19972 250502 19984
rect 385034 19972 385040 19984
rect 250496 19944 385040 19972
rect 250496 19932 250502 19944
rect 385034 19932 385040 19944
rect 385092 19932 385098 19984
rect 323578 19320 323584 19372
rect 323636 19360 323642 19372
rect 327074 19360 327080 19372
rect 323636 19332 327080 19360
rect 323636 19320 323642 19332
rect 327074 19320 327080 19332
rect 327132 19320 327138 19372
rect 222838 18640 222844 18692
rect 222896 18680 222902 18692
rect 245654 18680 245660 18692
rect 222896 18652 245660 18680
rect 222896 18640 222902 18652
rect 245654 18640 245660 18652
rect 245712 18680 245718 18692
rect 245712 18652 248414 18680
rect 245712 18640 245718 18652
rect 103422 18572 103428 18624
rect 103480 18612 103486 18624
rect 236730 18612 236736 18624
rect 103480 18584 236736 18612
rect 103480 18572 103486 18584
rect 236730 18572 236736 18584
rect 236788 18572 236794 18624
rect 248386 18612 248414 18652
rect 409966 18612 409972 18624
rect 248386 18584 409972 18612
rect 409966 18572 409972 18584
rect 410024 18572 410030 18624
rect 50982 17892 50988 17944
rect 51040 17932 51046 17944
rect 296714 17932 296720 17944
rect 51040 17904 296720 17932
rect 51040 17892 51046 17904
rect 296714 17892 296720 17904
rect 296772 17932 296778 17944
rect 297358 17932 297364 17944
rect 296772 17904 297364 17932
rect 296772 17892 296778 17904
rect 297358 17892 297364 17904
rect 297416 17892 297422 17944
rect 28810 17212 28816 17264
rect 28868 17252 28874 17264
rect 242158 17252 242164 17264
rect 28868 17224 242164 17252
rect 28868 17212 28874 17224
rect 242158 17212 242164 17224
rect 242216 17212 242222 17264
rect 243538 17212 243544 17264
rect 243596 17252 243602 17264
rect 413278 17252 413284 17264
rect 243596 17224 413284 17252
rect 243596 17212 243602 17224
rect 413278 17212 413284 17224
rect 413336 17212 413342 17264
rect 249150 16532 249156 16584
rect 249208 16572 249214 16584
rect 370590 16572 370596 16584
rect 249208 16544 370596 16572
rect 249208 16532 249214 16544
rect 370590 16532 370596 16544
rect 370648 16532 370654 16584
rect 126238 15920 126244 15972
rect 126296 15960 126302 15972
rect 214558 15960 214564 15972
rect 126296 15932 214564 15960
rect 126296 15920 126302 15932
rect 214558 15920 214564 15932
rect 214616 15920 214622 15972
rect 9582 15852 9588 15904
rect 9640 15892 9646 15904
rect 197998 15892 198004 15904
rect 9640 15864 198004 15892
rect 9640 15852 9646 15864
rect 197998 15852 198004 15864
rect 198056 15852 198062 15904
rect 341518 15852 341524 15904
rect 341576 15892 341582 15904
rect 342346 15892 342352 15904
rect 341576 15864 342352 15892
rect 341576 15852 341582 15864
rect 342346 15852 342352 15864
rect 342404 15892 342410 15904
rect 407758 15892 407764 15904
rect 342404 15864 407764 15892
rect 342404 15852 342410 15864
rect 407758 15852 407764 15864
rect 407816 15852 407822 15904
rect 248414 15172 248420 15224
rect 248472 15212 248478 15224
rect 249150 15212 249156 15224
rect 248472 15184 249156 15212
rect 248472 15172 248478 15184
rect 249150 15172 249156 15184
rect 249208 15172 249214 15224
rect 255866 15104 255872 15156
rect 255924 15144 255930 15156
rect 311158 15144 311164 15156
rect 255924 15116 311164 15144
rect 255924 15104 255930 15116
rect 311158 15104 311164 15116
rect 311216 15104 311222 15156
rect 96246 14424 96252 14476
rect 96304 14464 96310 14476
rect 218698 14464 218704 14476
rect 96304 14436 218704 14464
rect 96304 14424 96310 14436
rect 218698 14424 218704 14436
rect 218756 14424 218762 14476
rect 196618 13744 196624 13796
rect 196676 13784 196682 13796
rect 264330 13784 264336 13796
rect 196676 13756 264336 13784
rect 196676 13744 196682 13756
rect 264330 13744 264336 13756
rect 264388 13744 264394 13796
rect 280890 13744 280896 13796
rect 280948 13784 280954 13796
rect 367738 13784 367744 13796
rect 280948 13756 367744 13784
rect 280948 13744 280954 13756
rect 367738 13744 367744 13756
rect 367796 13744 367802 13796
rect 112806 13132 112812 13184
rect 112864 13172 112870 13184
rect 160738 13172 160744 13184
rect 112864 13144 160744 13172
rect 112864 13132 112870 13144
rect 160738 13132 160744 13144
rect 160796 13132 160802 13184
rect 45278 13064 45284 13116
rect 45336 13104 45342 13116
rect 224218 13104 224224 13116
rect 45336 13076 224224 13104
rect 45336 13064 45342 13076
rect 224218 13064 224224 13076
rect 224276 13064 224282 13116
rect 288342 13064 288348 13116
rect 288400 13104 288406 13116
rect 414658 13104 414664 13116
rect 288400 13076 414664 13104
rect 288400 13064 288406 13076
rect 414658 13064 414664 13076
rect 414716 13064 414722 13116
rect 280706 12452 280712 12504
rect 280764 12492 280770 12504
rect 280890 12492 280896 12504
rect 280764 12464 280896 12492
rect 280764 12452 280770 12464
rect 280890 12452 280896 12464
rect 280948 12452 280954 12504
rect 348050 12384 348056 12436
rect 348108 12424 348114 12436
rect 448514 12424 448520 12436
rect 348108 12396 448520 12424
rect 348108 12384 348114 12396
rect 448514 12384 448520 12396
rect 448572 12384 448578 12436
rect 268470 12316 268476 12368
rect 268528 12356 268534 12368
rect 349798 12356 349804 12368
rect 268528 12328 349804 12356
rect 268528 12316 268534 12328
rect 349798 12316 349804 12328
rect 349856 12316 349862 12368
rect 267734 11908 267740 11960
rect 267792 11948 267798 11960
rect 268470 11948 268476 11960
rect 267792 11920 268476 11948
rect 267792 11908 267798 11920
rect 268470 11908 268476 11920
rect 268528 11908 268534 11960
rect 135254 11772 135260 11824
rect 135312 11812 135318 11824
rect 136450 11812 136456 11824
rect 135312 11784 136456 11812
rect 135312 11772 135318 11784
rect 136450 11772 136456 11784
rect 136508 11772 136514 11824
rect 106826 11704 106832 11756
rect 106884 11744 106890 11756
rect 227070 11744 227076 11756
rect 106884 11716 227076 11744
rect 106884 11704 106890 11716
rect 227070 11704 227076 11716
rect 227128 11704 227134 11756
rect 242158 11704 242164 11756
rect 242216 11744 242222 11756
rect 264238 11744 264244 11756
rect 242216 11716 264244 11744
rect 242216 11704 242222 11716
rect 264238 11704 264244 11716
rect 264296 11704 264302 11756
rect 71498 10344 71504 10396
rect 71556 10384 71562 10396
rect 195238 10384 195244 10396
rect 71556 10356 195244 10384
rect 71556 10344 71562 10356
rect 195238 10344 195244 10356
rect 195296 10344 195302 10396
rect 311434 10344 311440 10396
rect 311492 10384 311498 10396
rect 378778 10384 378784 10396
rect 311492 10356 378784 10384
rect 311492 10344 311498 10356
rect 378778 10344 378784 10356
rect 378836 10344 378842 10396
rect 54938 10276 54944 10328
rect 54996 10316 55002 10328
rect 238110 10316 238116 10328
rect 54996 10288 238116 10316
rect 54996 10276 55002 10288
rect 238110 10276 238116 10288
rect 238168 10276 238174 10328
rect 261754 10276 261760 10328
rect 261812 10316 261818 10328
rect 449894 10316 449900 10328
rect 261812 10288 449900 10316
rect 261812 10276 261818 10288
rect 449894 10276 449900 10288
rect 449952 10276 449958 10328
rect 180426 9596 180432 9648
rect 180484 9636 180490 9648
rect 242894 9636 242900 9648
rect 180484 9608 242900 9636
rect 180484 9596 180490 9608
rect 242894 9596 242900 9608
rect 242952 9636 242958 9648
rect 243538 9636 243544 9648
rect 242952 9608 243544 9636
rect 242952 9596 242958 9608
rect 243538 9596 243544 9608
rect 243596 9596 243602 9648
rect 257338 9596 257344 9648
rect 257396 9636 257402 9648
rect 258718 9636 258724 9648
rect 257396 9608 258724 9636
rect 257396 9596 257402 9608
rect 258718 9596 258724 9608
rect 258776 9596 258782 9648
rect 334618 9596 334624 9648
rect 334676 9636 334682 9648
rect 337470 9636 337476 9648
rect 334676 9608 337476 9636
rect 334676 9596 334682 9608
rect 337470 9596 337476 9608
rect 337528 9596 337534 9648
rect 349982 9596 349988 9648
rect 350040 9636 350046 9648
rect 350442 9636 350448 9648
rect 350040 9608 350448 9636
rect 350040 9596 350046 9608
rect 350442 9596 350448 9608
rect 350500 9636 350506 9648
rect 439406 9636 439412 9648
rect 350500 9608 439412 9636
rect 350500 9596 350506 9608
rect 439406 9596 439412 9608
rect 439464 9596 439470 9648
rect 91554 8984 91560 9036
rect 91612 9024 91618 9036
rect 202230 9024 202236 9036
rect 91612 8996 202236 9024
rect 91612 8984 91618 8996
rect 202230 8984 202236 8996
rect 202288 8984 202294 9036
rect 332686 8984 332692 9036
rect 332744 9024 332750 9036
rect 349982 9024 349988 9036
rect 332744 8996 349988 9024
rect 332744 8984 332750 8996
rect 349982 8984 349988 8996
rect 350040 8984 350046 9036
rect 26510 8916 26516 8968
rect 26568 8956 26574 8968
rect 146938 8956 146944 8968
rect 26568 8928 146944 8956
rect 26568 8916 26574 8928
rect 146938 8916 146944 8928
rect 146996 8916 147002 8968
rect 327994 8916 328000 8968
rect 328052 8956 328058 8968
rect 358814 8956 358820 8968
rect 328052 8928 358820 8956
rect 328052 8916 328058 8928
rect 358814 8916 358820 8928
rect 358872 8916 358878 8968
rect 59630 7624 59636 7676
rect 59688 7664 59694 7676
rect 112438 7664 112444 7676
rect 59688 7636 112444 7664
rect 59688 7624 59694 7636
rect 112438 7624 112444 7636
rect 112496 7624 112502 7676
rect 117590 7624 117596 7676
rect 117648 7664 117654 7676
rect 206278 7664 206284 7676
rect 117648 7636 206284 7664
rect 117648 7624 117654 7636
rect 206278 7624 206284 7636
rect 206336 7624 206342 7676
rect 329190 7624 329196 7676
rect 329248 7664 329254 7676
rect 381630 7664 381636 7676
rect 329248 7636 381636 7664
rect 329248 7624 329254 7636
rect 381630 7624 381636 7636
rect 381688 7624 381694 7676
rect 66714 7556 66720 7608
rect 66772 7596 66778 7608
rect 240778 7596 240784 7608
rect 66772 7568 240784 7596
rect 66772 7556 66778 7568
rect 240778 7556 240784 7568
rect 240836 7556 240842 7608
rect 288986 7556 288992 7608
rect 289044 7596 289050 7608
rect 354030 7596 354036 7608
rect 289044 7568 354036 7596
rect 289044 7556 289050 7568
rect 354030 7556 354036 7568
rect 354088 7556 354094 7608
rect 308398 6808 308404 6860
rect 308456 6848 308462 6860
rect 309778 6848 309784 6860
rect 308456 6820 309784 6848
rect 308456 6808 308462 6820
rect 309778 6808 309784 6820
rect 309836 6808 309842 6860
rect 325050 6808 325056 6860
rect 325108 6848 325114 6860
rect 411622 6848 411628 6860
rect 325108 6820 411628 6848
rect 325108 6808 325114 6820
rect 411622 6808 411628 6820
rect 411680 6808 411686 6860
rect 24210 6196 24216 6248
rect 24268 6236 24274 6248
rect 191098 6236 191104 6248
rect 24268 6208 191104 6236
rect 24268 6196 24274 6208
rect 191098 6196 191104 6208
rect 191156 6196 191162 6248
rect 62022 6128 62028 6180
rect 62080 6168 62086 6180
rect 233878 6168 233884 6180
rect 62080 6140 233884 6168
rect 62080 6128 62086 6140
rect 233878 6128 233884 6140
rect 233936 6128 233942 6180
rect 278038 6128 278044 6180
rect 278096 6168 278102 6180
rect 285398 6168 285404 6180
rect 278096 6140 285404 6168
rect 278096 6128 278102 6140
rect 285398 6128 285404 6140
rect 285456 6168 285462 6180
rect 427906 6168 427912 6180
rect 285456 6140 427912 6168
rect 285456 6128 285462 6140
rect 427906 6128 427912 6140
rect 427964 6128 427970 6180
rect 282822 5516 282828 5568
rect 282880 5556 282886 5568
rect 283558 5556 283564 5568
rect 282880 5528 283564 5556
rect 282880 5516 282886 5528
rect 283558 5516 283564 5528
rect 283616 5516 283622 5568
rect 324498 5516 324504 5568
rect 324556 5556 324562 5568
rect 325050 5556 325056 5568
rect 324556 5528 325056 5556
rect 324556 5516 324562 5528
rect 325050 5516 325056 5528
rect 325108 5516 325114 5568
rect 306742 5448 306748 5500
rect 306800 5488 306806 5500
rect 307018 5488 307024 5500
rect 306800 5460 307024 5488
rect 306800 5448 306806 5460
rect 307018 5448 307024 5460
rect 307076 5488 307082 5500
rect 396718 5488 396724 5500
rect 307076 5460 396724 5488
rect 307076 5448 307082 5460
rect 396718 5448 396724 5460
rect 396776 5448 396782 5500
rect 105722 4768 105728 4820
rect 105780 4808 105786 4820
rect 186958 4808 186964 4820
rect 105780 4780 186964 4808
rect 105780 4768 105786 4780
rect 186958 4768 186964 4780
rect 187016 4768 187022 4820
rect 232590 4156 232596 4208
rect 232648 4196 232654 4208
rect 235810 4196 235816 4208
rect 232648 4168 235816 4196
rect 232648 4156 232654 4168
rect 235810 4156 235816 4168
rect 235868 4156 235874 4208
rect 247770 4088 247776 4140
rect 247828 4128 247834 4140
rect 250530 4128 250536 4140
rect 247828 4100 250536 4128
rect 247828 4088 247834 4100
rect 250530 4088 250536 4100
rect 250588 4088 250594 4140
rect 265342 4088 265348 4140
rect 265400 4128 265406 4140
rect 269758 4128 269764 4140
rect 265400 4100 269764 4128
rect 265400 4088 265406 4100
rect 269758 4088 269764 4100
rect 269816 4088 269822 4140
rect 279418 4088 279424 4140
rect 279476 4128 279482 4140
rect 286318 4128 286324 4140
rect 279476 4100 286324 4128
rect 279476 4088 279482 4100
rect 286318 4088 286324 4100
rect 286376 4088 286382 4140
rect 305546 4088 305552 4140
rect 305604 4128 305610 4140
rect 307110 4128 307116 4140
rect 305604 4100 307116 4128
rect 305604 4088 305610 4100
rect 307110 4088 307116 4100
rect 307168 4088 307174 4140
rect 315298 4088 315304 4140
rect 315356 4128 315362 4140
rect 319714 4128 319720 4140
rect 315356 4100 319720 4128
rect 315356 4088 315362 4100
rect 319714 4088 319720 4100
rect 319772 4088 319778 4140
rect 326338 4088 326344 4140
rect 326396 4128 326402 4140
rect 326798 4128 326804 4140
rect 326396 4100 326804 4128
rect 326396 4088 326402 4100
rect 326798 4088 326804 4100
rect 326856 4128 326862 4140
rect 329098 4128 329104 4140
rect 326856 4100 329104 4128
rect 326856 4088 326862 4100
rect 329098 4088 329104 4100
rect 329156 4088 329162 4140
rect 268378 4020 268384 4072
rect 268436 4060 268442 4072
rect 268838 4060 268844 4072
rect 268436 4032 268844 4060
rect 268436 4020 268442 4032
rect 268838 4020 268844 4032
rect 268896 4020 268902 4072
rect 302878 4020 302884 4072
rect 302936 4060 302942 4072
rect 309870 4060 309876 4072
rect 302936 4032 309876 4060
rect 302936 4020 302942 4032
rect 309870 4020 309876 4032
rect 309928 4020 309934 4072
rect 345750 4020 345756 4072
rect 345808 4060 345814 4072
rect 402974 4060 402980 4072
rect 345808 4032 402980 4060
rect 345808 4020 345814 4032
rect 402974 4020 402980 4032
rect 403032 4020 403038 4072
rect 254670 3748 254676 3800
rect 254728 3788 254734 3800
rect 258074 3788 258080 3800
rect 254728 3760 258080 3788
rect 254728 3748 254734 3760
rect 258074 3748 258080 3760
rect 258132 3748 258138 3800
rect 351178 3612 351184 3664
rect 351236 3652 351242 3664
rect 351638 3652 351644 3664
rect 351236 3624 351644 3652
rect 351236 3612 351242 3624
rect 351638 3612 351644 3624
rect 351696 3612 351702 3664
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 12250 3584 12256 3596
rect 11204 3556 12256 3584
rect 11204 3544 11210 3556
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 20530 3544 20536 3596
rect 20588 3584 20594 3596
rect 20588 3556 20760 3584
rect 20588 3544 20594 3556
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 4062 3516 4068 3528
rect 2924 3488 4068 3516
rect 2924 3476 2930 3488
rect 4062 3476 4068 3488
rect 4120 3476 4126 3528
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 9582 3516 9588 3528
rect 8812 3488 9588 3516
rect 8812 3476 8818 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 16482 3516 16488 3528
rect 15988 3488 16488 3516
rect 15988 3476 15994 3488
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 17862 3516 17868 3528
rect 17092 3488 17868 3516
rect 17092 3476 17098 3488
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 19242 3516 19248 3528
rect 18288 3488 19248 3516
rect 18288 3476 18294 3488
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 20622 3516 20628 3528
rect 19484 3488 20628 3516
rect 19484 3476 19490 3488
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 20732 3516 20760 3556
rect 25314 3544 25320 3596
rect 25372 3584 25378 3596
rect 26142 3584 26148 3596
rect 25372 3556 26148 3584
rect 25372 3544 25378 3556
rect 26142 3544 26148 3556
rect 26200 3544 26206 3596
rect 27706 3544 27712 3596
rect 27764 3584 27770 3596
rect 28810 3584 28816 3596
rect 27764 3556 28816 3584
rect 27764 3544 27770 3556
rect 28810 3544 28816 3556
rect 28868 3544 28874 3596
rect 32398 3544 32404 3596
rect 32456 3584 32462 3596
rect 33042 3584 33048 3596
rect 32456 3556 33048 3584
rect 32456 3544 32462 3556
rect 33042 3544 33048 3556
rect 33100 3544 33106 3596
rect 33594 3544 33600 3596
rect 33652 3584 33658 3596
rect 34422 3584 34428 3596
rect 33652 3556 34428 3584
rect 33652 3544 33658 3556
rect 34422 3544 34428 3556
rect 34480 3544 34486 3596
rect 34790 3544 34796 3596
rect 34848 3584 34854 3596
rect 35802 3584 35808 3596
rect 34848 3556 35808 3584
rect 34848 3544 34854 3556
rect 35802 3544 35808 3556
rect 35860 3544 35866 3596
rect 35986 3544 35992 3596
rect 36044 3584 36050 3596
rect 37090 3584 37096 3596
rect 36044 3556 37096 3584
rect 36044 3544 36050 3556
rect 37090 3544 37096 3556
rect 37148 3544 37154 3596
rect 40678 3544 40684 3596
rect 40736 3584 40742 3596
rect 41322 3584 41328 3596
rect 40736 3556 41328 3584
rect 40736 3544 40742 3556
rect 41322 3544 41328 3556
rect 41380 3544 41386 3596
rect 41874 3544 41880 3596
rect 41932 3584 41938 3596
rect 42702 3584 42708 3596
rect 41932 3556 42708 3584
rect 41932 3544 41938 3556
rect 42702 3544 42708 3556
rect 42760 3544 42766 3596
rect 43070 3544 43076 3596
rect 43128 3584 43134 3596
rect 44082 3584 44088 3596
rect 43128 3556 44088 3584
rect 43128 3544 43134 3556
rect 44082 3544 44088 3556
rect 44140 3544 44146 3596
rect 44266 3544 44272 3596
rect 44324 3584 44330 3596
rect 45370 3584 45376 3596
rect 44324 3556 45376 3584
rect 44324 3544 44330 3556
rect 45370 3544 45376 3556
rect 45428 3544 45434 3596
rect 54478 3584 54484 3596
rect 45526 3556 54484 3584
rect 45526 3516 45554 3556
rect 54478 3544 54484 3556
rect 54536 3544 54542 3596
rect 64322 3544 64328 3596
rect 64380 3584 64386 3596
rect 64782 3584 64788 3596
rect 64380 3556 64788 3584
rect 64380 3544 64386 3556
rect 64782 3544 64788 3556
rect 64840 3544 64846 3596
rect 71038 3584 71044 3596
rect 65444 3556 71044 3584
rect 20732 3488 45554 3516
rect 48958 3476 48964 3528
rect 49016 3516 49022 3528
rect 49602 3516 49608 3528
rect 49016 3488 49608 3516
rect 49016 3476 49022 3488
rect 49602 3476 49608 3488
rect 49660 3476 49666 3528
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50890 3516 50896 3528
rect 50212 3488 50896 3516
rect 50212 3476 50218 3488
rect 50890 3476 50896 3488
rect 50948 3476 50954 3528
rect 52546 3476 52552 3528
rect 52604 3516 52610 3528
rect 53650 3516 53656 3528
rect 52604 3488 53656 3516
rect 52604 3476 52610 3488
rect 53650 3476 53656 3488
rect 53708 3476 53714 3528
rect 56042 3476 56048 3528
rect 56100 3516 56106 3528
rect 56502 3516 56508 3528
rect 56100 3488 56508 3516
rect 56100 3476 56106 3488
rect 56502 3476 56508 3488
rect 56560 3476 56566 3528
rect 57238 3476 57244 3528
rect 57296 3516 57302 3528
rect 57790 3516 57796 3528
rect 57296 3488 57796 3516
rect 57296 3476 57302 3488
rect 57790 3476 57796 3488
rect 57848 3476 57854 3528
rect 58434 3476 58440 3528
rect 58492 3516 58498 3528
rect 59262 3516 59268 3528
rect 58492 3488 59268 3516
rect 58492 3476 58498 3488
rect 59262 3476 59268 3488
rect 59320 3476 59326 3528
rect 60826 3476 60832 3528
rect 60884 3516 60890 3528
rect 61930 3516 61936 3528
rect 60884 3488 61936 3516
rect 60884 3476 60890 3488
rect 61930 3476 61936 3488
rect 61988 3476 61994 3528
rect 63218 3476 63224 3528
rect 63276 3516 63282 3528
rect 65444 3516 65472 3556
rect 71038 3544 71044 3556
rect 71096 3544 71102 3596
rect 78490 3544 78496 3596
rect 78548 3584 78554 3596
rect 78548 3556 78720 3584
rect 78548 3544 78554 3556
rect 63276 3488 65472 3516
rect 63276 3476 63282 3488
rect 65518 3476 65524 3528
rect 65576 3516 65582 3528
rect 66162 3516 66168 3528
rect 65576 3488 66168 3516
rect 65576 3476 65582 3488
rect 66162 3476 66168 3488
rect 66220 3476 66226 3528
rect 67910 3476 67916 3528
rect 67968 3516 67974 3528
rect 68922 3516 68928 3528
rect 67968 3488 68928 3516
rect 67968 3476 67974 3488
rect 68922 3476 68928 3488
rect 68980 3476 68986 3528
rect 69106 3476 69112 3528
rect 69164 3516 69170 3528
rect 70210 3516 70216 3528
rect 69164 3488 70216 3516
rect 69164 3476 69170 3488
rect 70210 3476 70216 3488
rect 70268 3476 70274 3528
rect 72602 3476 72608 3528
rect 72660 3516 72666 3528
rect 73062 3516 73068 3528
rect 72660 3488 73068 3516
rect 72660 3476 72666 3488
rect 73062 3476 73068 3488
rect 73120 3476 73126 3528
rect 73798 3476 73804 3528
rect 73856 3516 73862 3528
rect 74442 3516 74448 3528
rect 73856 3488 74448 3516
rect 73856 3476 73862 3488
rect 74442 3476 74448 3488
rect 74500 3476 74506 3528
rect 74994 3476 75000 3528
rect 75052 3516 75058 3528
rect 75822 3516 75828 3528
rect 75052 3488 75828 3516
rect 75052 3476 75058 3488
rect 75822 3476 75828 3488
rect 75880 3476 75886 3528
rect 76190 3476 76196 3528
rect 76248 3516 76254 3528
rect 77202 3516 77208 3528
rect 76248 3488 77208 3516
rect 76248 3476 76254 3488
rect 77202 3476 77208 3488
rect 77260 3476 77266 3528
rect 77386 3476 77392 3528
rect 77444 3516 77450 3528
rect 78582 3516 78588 3528
rect 77444 3488 78588 3516
rect 77444 3476 77450 3488
rect 78582 3476 78588 3488
rect 78640 3476 78646 3528
rect 78692 3516 78720 3556
rect 80882 3544 80888 3596
rect 80940 3584 80946 3596
rect 81342 3584 81348 3596
rect 80940 3556 81348 3584
rect 80940 3544 80946 3556
rect 81342 3544 81348 3556
rect 81400 3544 81406 3596
rect 83274 3544 83280 3596
rect 83332 3584 83338 3596
rect 84102 3584 84108 3596
rect 83332 3556 84108 3584
rect 83332 3544 83338 3556
rect 84102 3544 84108 3556
rect 84160 3544 84166 3596
rect 87598 3584 87604 3596
rect 84396 3556 87604 3584
rect 84396 3516 84424 3556
rect 87598 3544 87604 3556
rect 87656 3544 87662 3596
rect 126238 3584 126244 3596
rect 122806 3556 126244 3584
rect 78692 3488 84424 3516
rect 84470 3476 84476 3528
rect 84528 3516 84534 3528
rect 85482 3516 85488 3528
rect 84528 3488 85488 3516
rect 84528 3476 84534 3488
rect 85482 3476 85488 3488
rect 85540 3476 85546 3528
rect 89162 3476 89168 3528
rect 89220 3516 89226 3528
rect 89622 3516 89628 3528
rect 89220 3488 89628 3516
rect 89220 3476 89226 3488
rect 89622 3476 89628 3488
rect 89680 3476 89686 3528
rect 90358 3476 90364 3528
rect 90416 3516 90422 3528
rect 91002 3516 91008 3528
rect 90416 3488 91008 3516
rect 90416 3476 90422 3488
rect 91002 3476 91008 3488
rect 91060 3476 91066 3528
rect 92750 3476 92756 3528
rect 92808 3516 92814 3528
rect 93762 3516 93768 3528
rect 92808 3488 93768 3516
rect 92808 3476 92814 3488
rect 93762 3476 93768 3488
rect 93820 3476 93826 3528
rect 93946 3476 93952 3528
rect 94004 3516 94010 3528
rect 95050 3516 95056 3528
rect 94004 3488 95056 3516
rect 94004 3476 94010 3488
rect 95050 3476 95056 3488
rect 95108 3476 95114 3528
rect 97442 3476 97448 3528
rect 97500 3516 97506 3528
rect 97902 3516 97908 3528
rect 97500 3488 97908 3516
rect 97500 3476 97506 3488
rect 97902 3476 97908 3488
rect 97960 3476 97966 3528
rect 98638 3476 98644 3528
rect 98696 3516 98702 3528
rect 99282 3516 99288 3528
rect 98696 3488 99288 3516
rect 98696 3476 98702 3488
rect 99282 3476 99288 3488
rect 99340 3476 99346 3528
rect 99834 3476 99840 3528
rect 99892 3516 99898 3528
rect 100662 3516 100668 3528
rect 99892 3488 100668 3516
rect 99892 3476 99898 3488
rect 100662 3476 100668 3488
rect 100720 3476 100726 3528
rect 101030 3476 101036 3528
rect 101088 3516 101094 3528
rect 102042 3516 102048 3528
rect 101088 3488 102048 3516
rect 101088 3476 101094 3488
rect 102042 3476 102048 3488
rect 102100 3476 102106 3528
rect 106918 3476 106924 3528
rect 106976 3516 106982 3528
rect 107562 3516 107568 3528
rect 106976 3488 107568 3516
rect 106976 3476 106982 3488
rect 107562 3476 107568 3488
rect 107620 3476 107626 3528
rect 108114 3476 108120 3528
rect 108172 3516 108178 3528
rect 108942 3516 108948 3528
rect 108172 3488 108948 3516
rect 108172 3476 108178 3488
rect 108942 3476 108948 3488
rect 109000 3476 109006 3528
rect 109310 3476 109316 3528
rect 109368 3516 109374 3528
rect 122806 3516 122834 3556
rect 126238 3544 126244 3556
rect 126296 3544 126302 3596
rect 109368 3488 122834 3516
rect 109368 3476 109374 3488
rect 124674 3476 124680 3528
rect 124732 3516 124738 3528
rect 125502 3516 125508 3528
rect 124732 3488 125508 3516
rect 124732 3476 124738 3488
rect 125502 3476 125508 3488
rect 125560 3476 125566 3528
rect 125870 3476 125876 3528
rect 125928 3516 125934 3528
rect 126882 3516 126888 3528
rect 125928 3488 126888 3516
rect 125928 3476 125934 3488
rect 126882 3476 126888 3488
rect 126940 3476 126946 3528
rect 129366 3476 129372 3528
rect 129424 3516 129430 3528
rect 130378 3516 130384 3528
rect 129424 3488 130384 3516
rect 129424 3476 129430 3488
rect 130378 3476 130384 3488
rect 130436 3476 130442 3528
rect 140038 3476 140044 3528
rect 140096 3516 140102 3528
rect 141418 3516 141424 3528
rect 140096 3488 141424 3516
rect 140096 3476 140102 3488
rect 141418 3476 141424 3488
rect 141476 3476 141482 3528
rect 143534 3476 143540 3528
rect 143592 3516 143598 3528
rect 144822 3516 144828 3528
rect 143592 3488 144828 3516
rect 143592 3476 143598 3488
rect 144822 3476 144828 3488
rect 144880 3476 144886 3528
rect 251174 3476 251180 3528
rect 251232 3516 251238 3528
rect 251910 3516 251916 3528
rect 251232 3488 251916 3516
rect 251232 3476 251238 3488
rect 251910 3476 251916 3488
rect 251968 3476 251974 3528
rect 258258 3476 258264 3528
rect 258316 3516 258322 3528
rect 258718 3516 258724 3528
rect 258316 3488 258724 3516
rect 258316 3476 258322 3488
rect 258718 3476 258724 3488
rect 258776 3476 258782 3528
rect 272426 3476 272432 3528
rect 272484 3516 272490 3528
rect 273254 3516 273260 3528
rect 272484 3488 273260 3516
rect 272484 3476 272490 3488
rect 273254 3476 273260 3488
rect 273312 3476 273318 3528
rect 273622 3476 273628 3528
rect 273680 3516 273686 3528
rect 274542 3516 274548 3528
rect 273680 3488 274548 3516
rect 273680 3476 273686 3488
rect 274542 3476 274548 3488
rect 274600 3476 274606 3528
rect 292482 3476 292488 3528
rect 292540 3516 292546 3528
rect 294874 3516 294880 3528
rect 292540 3488 294880 3516
rect 292540 3476 292546 3488
rect 294874 3476 294880 3488
rect 294932 3476 294938 3528
rect 296714 3476 296720 3528
rect 296772 3516 296778 3528
rect 297266 3516 297272 3528
rect 296772 3488 297272 3516
rect 296772 3476 296778 3488
rect 297266 3476 297272 3488
rect 297324 3476 297330 3528
rect 307938 3476 307944 3528
rect 307996 3516 308002 3528
rect 309134 3516 309140 3528
rect 307996 3488 309140 3516
rect 307996 3476 308002 3488
rect 309134 3476 309140 3488
rect 309192 3476 309198 3528
rect 313826 3476 313832 3528
rect 313884 3516 313890 3528
rect 314562 3516 314568 3528
rect 313884 3488 314568 3516
rect 313884 3476 313890 3488
rect 314562 3476 314568 3488
rect 314620 3476 314626 3528
rect 316034 3476 316040 3528
rect 316092 3516 316098 3528
rect 317322 3516 317328 3528
rect 316092 3488 317328 3516
rect 316092 3476 316098 3488
rect 317322 3476 317328 3488
rect 317380 3476 317386 3528
rect 324406 3476 324412 3528
rect 324464 3516 324470 3528
rect 325602 3516 325608 3528
rect 324464 3488 325608 3516
rect 324464 3476 324470 3488
rect 325602 3476 325608 3488
rect 325660 3476 325666 3528
rect 332594 3476 332600 3528
rect 332652 3516 332658 3528
rect 333882 3516 333888 3528
rect 332652 3488 333888 3516
rect 332652 3476 332658 3488
rect 333882 3476 333888 3488
rect 333940 3476 333946 3528
rect 339862 3476 339868 3528
rect 339920 3516 339926 3528
rect 340782 3516 340788 3528
rect 339920 3488 340788 3516
rect 339920 3476 339926 3488
rect 340782 3476 340788 3488
rect 340840 3476 340846 3528
rect 340966 3476 340972 3528
rect 341024 3516 341030 3528
rect 342346 3516 342352 3528
rect 341024 3488 342352 3516
rect 341024 3476 341030 3488
rect 342346 3476 342352 3488
rect 342404 3476 342410 3528
rect 582190 3476 582196 3528
rect 582248 3516 582254 3528
rect 583570 3516 583576 3528
rect 582248 3488 583576 3516
rect 582248 3476 582254 3488
rect 583570 3476 583576 3488
rect 583628 3476 583634 3528
rect 106826 3448 106832 3460
rect 4080 3420 106832 3448
rect 4080 3392 4108 3420
rect 106826 3408 106832 3420
rect 106884 3408 106890 3460
rect 114002 3408 114008 3460
rect 114060 3448 114066 3460
rect 114462 3448 114468 3460
rect 114060 3420 114468 3448
rect 114060 3408 114066 3420
rect 114462 3408 114468 3420
rect 114520 3408 114526 3460
rect 115198 3408 115204 3460
rect 115256 3448 115262 3460
rect 115842 3448 115848 3460
rect 115256 3420 115848 3448
rect 115256 3408 115262 3420
rect 115842 3408 115848 3420
rect 115900 3408 115906 3460
rect 116394 3408 116400 3460
rect 116452 3448 116458 3460
rect 117222 3448 117228 3460
rect 116452 3420 117228 3448
rect 116452 3408 116458 3420
rect 117222 3408 117228 3420
rect 117280 3408 117286 3460
rect 122282 3408 122288 3460
rect 122340 3448 122346 3460
rect 122742 3448 122748 3460
rect 122340 3420 122748 3448
rect 122340 3408 122346 3420
rect 122742 3408 122748 3420
rect 122800 3408 122806 3460
rect 123478 3408 123484 3460
rect 123536 3448 123542 3460
rect 220078 3448 220084 3460
rect 123536 3420 220084 3448
rect 123536 3408 123542 3420
rect 220078 3408 220084 3420
rect 220136 3408 220142 3460
rect 245654 3408 245660 3460
rect 245712 3448 245718 3460
rect 257062 3448 257068 3460
rect 245712 3420 257068 3448
rect 245712 3408 245718 3420
rect 257062 3408 257068 3420
rect 257120 3408 257126 3460
rect 276106 3408 276112 3460
rect 276164 3448 276170 3460
rect 277118 3448 277124 3460
rect 276164 3420 277124 3448
rect 276164 3408 276170 3420
rect 277118 3408 277124 3420
rect 277176 3448 277182 3460
rect 282178 3448 282184 3460
rect 277176 3420 282184 3448
rect 277176 3408 277182 3420
rect 282178 3408 282184 3420
rect 282236 3408 282242 3460
rect 312630 3408 312636 3460
rect 312688 3448 312694 3460
rect 323670 3448 323676 3460
rect 312688 3420 323676 3448
rect 312688 3408 312694 3420
rect 323670 3408 323676 3420
rect 323728 3408 323734 3460
rect 349246 3408 349252 3460
rect 349304 3448 349310 3460
rect 360838 3448 360844 3460
rect 349304 3420 360844 3448
rect 349304 3408 349310 3420
rect 360838 3408 360844 3420
rect 360896 3408 360902 3460
rect 4062 3340 4068 3392
rect 4120 3340 4126 3392
rect 240502 3340 240508 3392
rect 240560 3380 240566 3392
rect 246390 3380 246396 3392
rect 240560 3352 246396 3380
rect 240560 3340 240566 3352
rect 246390 3340 246396 3352
rect 246448 3340 246454 3392
rect 241698 3272 241704 3324
rect 241756 3312 241762 3324
rect 244918 3312 244924 3324
rect 241756 3284 244924 3312
rect 241756 3272 241762 3284
rect 244918 3272 244924 3284
rect 244976 3272 244982 3324
rect 110506 3068 110512 3120
rect 110564 3108 110570 3120
rect 111518 3108 111524 3120
rect 110564 3080 111524 3108
rect 110564 3068 110570 3080
rect 111518 3068 111524 3080
rect 111576 3068 111582 3120
rect 580994 3068 581000 3120
rect 581052 3108 581058 3120
rect 583754 3108 583760 3120
rect 581052 3080 583760 3108
rect 581052 3068 581058 3080
rect 583754 3068 583760 3080
rect 583812 3068 583818 3120
rect 245194 2932 245200 2984
rect 245252 2972 245258 2984
rect 247034 2972 247040 2984
rect 245252 2944 247040 2972
rect 245252 2932 245258 2944
rect 247034 2932 247040 2944
rect 247092 2932 247098 2984
rect 271782 2728 271788 2780
rect 271840 2768 271846 2780
rect 445846 2768 445852 2780
rect 271840 2740 445852 2768
rect 271840 2728 271846 2740
rect 445846 2728 445852 2740
rect 445904 2728 445910 2780
rect 51350 2116 51356 2168
rect 51408 2156 51414 2168
rect 59998 2156 60004 2168
rect 51408 2128 60004 2156
rect 51408 2116 51414 2128
rect 59998 2116 60004 2128
rect 60056 2116 60062 2168
rect 102226 2116 102232 2168
rect 102284 2156 102290 2168
rect 213178 2156 213184 2168
rect 102284 2128 213184 2156
rect 102284 2116 102290 2128
rect 213178 2116 213184 2128
rect 213236 2116 213242 2168
rect 239306 2116 239312 2168
rect 239364 2156 239370 2168
rect 270586 2156 270592 2168
rect 239364 2128 270592 2156
rect 239364 2116 239370 2128
rect 270586 2116 270592 2128
rect 270644 2156 270650 2168
rect 271782 2156 271788 2168
rect 270644 2128 271788 2156
rect 270644 2116 270650 2128
rect 271782 2116 271788 2128
rect 271840 2116 271846 2168
rect 7650 2048 7656 2100
rect 7708 2088 7714 2100
rect 105538 2088 105544 2100
rect 7708 2060 105544 2088
rect 7708 2048 7714 2060
rect 105538 2048 105544 2060
rect 105596 2048 105602 2100
rect 118786 2048 118792 2100
rect 118844 2088 118850 2100
rect 242158 2088 242164 2100
rect 118844 2060 242164 2088
rect 118844 2048 118850 2060
rect 242158 2048 242164 2060
rect 242216 2048 242222 2100
<< via1 >>
rect 62028 702992 62080 703044
rect 267648 702992 267700 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 169760 702924 169812 702976
rect 170312 702924 170364 702976
rect 281540 702924 281592 702976
rect 283840 702924 283892 702976
rect 351920 702924 351972 702976
rect 202788 702856 202840 702908
rect 273260 702856 273312 702908
rect 276020 702856 276072 702908
rect 478512 702856 478564 702908
rect 130384 702788 130436 702840
rect 218980 702788 219032 702840
rect 349804 702788 349856 702840
rect 494796 702788 494848 702840
rect 233884 702720 233936 702772
rect 397368 702720 397420 702772
rect 67640 702652 67692 702704
rect 169760 702652 169812 702704
rect 197268 702652 197320 702704
rect 364984 702652 365036 702704
rect 381544 702652 381596 702704
rect 462320 702652 462372 702704
rect 24308 702584 24360 702636
rect 79324 702584 79376 702636
rect 95148 702584 95200 702636
rect 300124 702584 300176 702636
rect 356152 702584 356204 702636
rect 360844 702584 360896 702636
rect 543464 702584 543516 702636
rect 88248 702516 88300 702568
rect 235172 702516 235224 702568
rect 264244 702516 264296 702568
rect 559656 702516 559708 702568
rect 8116 702448 8168 702500
rect 88800 702448 88852 702500
rect 93768 702448 93820 702500
rect 527180 702448 527232 702500
rect 75184 700272 75236 700324
rect 105452 700272 105504 700324
rect 124864 700272 124916 700324
rect 137836 700272 137888 700324
rect 327724 700272 327776 700324
rect 348792 700272 348844 700324
rect 376116 700272 376168 700324
rect 429844 700272 429896 700324
rect 66168 699660 66220 699712
rect 72976 699660 73028 699712
rect 86868 699660 86920 699712
rect 89168 699660 89220 699712
rect 3516 670692 3568 670744
rect 14464 670692 14516 670744
rect 2780 656956 2832 657008
rect 4804 656956 4856 657008
rect 3516 632068 3568 632120
rect 21364 632068 21416 632120
rect 3516 618264 3568 618316
rect 22744 618264 22796 618316
rect 3516 605820 3568 605872
rect 90364 605820 90416 605872
rect 67456 598952 67508 599004
rect 259460 598952 259512 599004
rect 82820 597524 82872 597576
rect 111156 597524 111208 597576
rect 79968 596776 80020 596828
rect 86868 596776 86920 596828
rect 92480 596776 92532 596828
rect 70308 596164 70360 596216
rect 349804 596164 349856 596216
rect 85948 594804 86000 594856
rect 155224 594804 155276 594856
rect 40040 594056 40092 594108
rect 89812 594056 89864 594108
rect 90364 593784 90416 593836
rect 91192 593784 91244 593836
rect 88248 593376 88300 593428
rect 113180 593376 113232 593428
rect 67364 592628 67416 592680
rect 75184 592628 75236 592680
rect 75644 592084 75696 592136
rect 96620 592084 96672 592136
rect 84108 592016 84160 592068
rect 111800 592016 111852 592068
rect 79324 591472 79376 591524
rect 80704 591472 80756 591524
rect 4804 591268 4856 591320
rect 69112 591268 69164 591320
rect 72148 590792 72200 590844
rect 79968 590792 80020 590844
rect 69112 590724 69164 590776
rect 71688 590724 71740 590776
rect 78588 590724 78640 590776
rect 93124 590724 93176 590776
rect 70124 590656 70176 590708
rect 74448 590656 74500 590708
rect 85028 590656 85080 590708
rect 88248 590656 88300 590708
rect 71688 589976 71740 590028
rect 89076 589976 89128 590028
rect 74908 589908 74960 589960
rect 75644 589908 75696 589960
rect 80704 589908 80756 589960
rect 106924 589908 106976 589960
rect 7564 589296 7616 589348
rect 74908 589296 74960 589348
rect 81900 588548 81952 588600
rect 94504 588548 94556 588600
rect 76104 588412 76156 588464
rect 88984 588140 89036 588192
rect 55128 587868 55180 587920
rect 66812 587868 66864 587920
rect 67548 587868 67600 587920
rect 351920 587868 351972 587920
rect 88800 587120 88852 587172
rect 115204 587120 115256 587172
rect 88984 586576 89036 586628
rect 98736 586576 98788 586628
rect 59084 586508 59136 586560
rect 66260 586508 66312 586560
rect 57888 585148 57940 585200
rect 66904 585148 66956 585200
rect 91284 584400 91336 584452
rect 95148 584400 95200 584452
rect 128360 584400 128412 584452
rect 93768 583720 93820 583772
rect 116584 583720 116636 583772
rect 91836 583652 91888 583704
rect 50896 582360 50948 582412
rect 66812 582360 66864 582412
rect 64696 581000 64748 581052
rect 66536 581000 66588 581052
rect 91284 581000 91336 581052
rect 108304 581000 108356 581052
rect 3056 580728 3108 580780
rect 7564 580728 7616 580780
rect 61936 579640 61988 579692
rect 66812 579640 66864 579692
rect 91284 576852 91336 576904
rect 111064 576852 111116 576904
rect 21364 576104 21416 576156
rect 39948 576104 40000 576156
rect 91192 576104 91244 576156
rect 122840 576104 122892 576156
rect 39948 575492 40000 575544
rect 66812 575492 66864 575544
rect 93124 574744 93176 574796
rect 103520 574744 103572 574796
rect 104164 574132 104216 574184
rect 109684 574132 109736 574184
rect 61844 574064 61896 574116
rect 67364 574064 67416 574116
rect 91744 574064 91796 574116
rect 136640 574064 136692 574116
rect 91744 572704 91796 572756
rect 112444 572704 112496 572756
rect 91192 571412 91244 571464
rect 94596 571412 94648 571464
rect 63316 571344 63368 571396
rect 66812 571344 66864 571396
rect 91744 571344 91796 571396
rect 122196 571344 122248 571396
rect 174544 569916 174596 569968
rect 341524 569916 341576 569968
rect 48136 569168 48188 569220
rect 67088 569168 67140 569220
rect 177948 568556 178000 568608
rect 320180 568556 320232 568608
rect 64788 567196 64840 567248
rect 66812 567196 66864 567248
rect 89812 567196 89864 567248
rect 133144 567196 133196 567248
rect 155868 567196 155920 567248
rect 311900 567196 311952 567248
rect 94596 566448 94648 566500
rect 138020 566448 138072 566500
rect 3240 565836 3292 565888
rect 43444 565836 43496 565888
rect 53656 565836 53708 565888
rect 67640 565836 67692 565888
rect 91560 565836 91612 565888
rect 116676 565836 116728 565888
rect 138020 565836 138072 565888
rect 213920 565836 213972 565888
rect 93124 565088 93176 565140
rect 133880 565088 133932 565140
rect 135168 565088 135220 565140
rect 55864 564408 55916 564460
rect 66812 564408 66864 564460
rect 91560 564408 91612 564460
rect 107016 564408 107068 564460
rect 135168 564408 135220 564460
rect 291200 564408 291252 564460
rect 52276 563048 52328 563100
rect 66812 563048 66864 563100
rect 91560 563048 91612 563100
rect 106188 563048 106240 563100
rect 191104 563048 191156 563100
rect 357440 563048 357492 563100
rect 106188 562300 106240 562352
rect 197360 562300 197412 562352
rect 197360 561756 197412 561808
rect 241520 561756 241572 561808
rect 37188 561688 37240 561740
rect 66812 561688 66864 561740
rect 186964 561688 187016 561740
rect 267740 561688 267792 561740
rect 263600 561620 263652 561672
rect 264244 561620 264296 561672
rect 178684 560328 178736 560380
rect 263600 560328 263652 560380
rect 41328 560260 41380 560312
rect 66812 560260 66864 560312
rect 111156 560260 111208 560312
rect 111708 560260 111760 560312
rect 359004 560260 359056 560312
rect 133144 560192 133196 560244
rect 133788 560192 133840 560244
rect 133788 558968 133840 559020
rect 209780 558968 209832 559020
rect 89628 558900 89680 558952
rect 129740 558900 129792 558952
rect 195888 558900 195940 558952
rect 288440 558900 288492 558952
rect 59176 558288 59228 558340
rect 62028 558288 62080 558340
rect 97264 558152 97316 558204
rect 118516 558152 118568 558204
rect 198648 558152 198700 558204
rect 582472 558152 582524 558204
rect 62028 557540 62080 557592
rect 66812 557540 66864 557592
rect 188344 557540 188396 557592
rect 268384 557540 268436 557592
rect 91100 557472 91152 557524
rect 91284 557472 91336 557524
rect 92296 556792 92348 556844
rect 148416 556792 148468 556844
rect 180156 556248 180208 556300
rect 248512 556248 248564 556300
rect 91100 556180 91152 556232
rect 122104 556180 122156 556232
rect 155316 556180 155368 556232
rect 207020 556180 207072 556232
rect 582472 556180 582524 556232
rect 190368 554820 190420 554872
rect 235264 554820 235316 554872
rect 43996 554752 44048 554804
rect 66812 554752 66864 554804
rect 91100 554752 91152 554804
rect 106188 554752 106240 554804
rect 247040 554752 247092 554804
rect 580356 554752 580408 554804
rect 57796 554004 57848 554056
rect 66628 554004 66680 554056
rect 2780 553800 2832 553852
rect 4804 553800 4856 553852
rect 197176 553460 197228 553512
rect 287060 553460 287112 553512
rect 118516 553392 118568 553444
rect 212540 553392 212592 553444
rect 91100 552100 91152 552152
rect 101404 552100 101456 552152
rect 184296 552100 184348 552152
rect 226984 552100 227036 552152
rect 91376 552032 91428 552084
rect 108396 552032 108448 552084
rect 192484 552032 192536 552084
rect 270500 552032 270552 552084
rect 198832 551284 198884 551336
rect 331220 551284 331272 551336
rect 182916 550672 182968 550724
rect 238760 550672 238812 550724
rect 91100 550604 91152 550656
rect 124220 550604 124272 550656
rect 187148 550604 187200 550656
rect 199844 549312 199896 549364
rect 251824 549312 251876 549364
rect 60648 549244 60700 549296
rect 66812 549244 66864 549296
rect 91100 549244 91152 549296
rect 97908 549244 97960 549296
rect 278044 549244 278096 549296
rect 90456 549176 90508 549228
rect 91284 549176 91336 549228
rect 193864 547952 193916 548004
rect 237380 547952 237432 548004
rect 59268 547884 59320 547936
rect 66812 547884 66864 547936
rect 91284 547884 91336 547936
rect 95240 547884 95292 547936
rect 177856 547884 177908 547936
rect 284300 547884 284352 547936
rect 95240 547136 95292 547188
rect 245660 547136 245712 547188
rect 52368 546456 52420 546508
rect 66812 546456 66864 546508
rect 185584 546456 185636 546508
rect 229100 546456 229152 546508
rect 324320 545572 324372 545624
rect 324872 545572 324924 545624
rect 327724 545572 327776 545624
rect 188436 545164 188488 545216
rect 324320 545164 324372 545216
rect 327080 545164 327132 545216
rect 367100 545164 367152 545216
rect 50988 545096 51040 545148
rect 66812 545096 66864 545148
rect 91560 545096 91612 545148
rect 97264 545096 97316 545148
rect 137928 545096 137980 545148
rect 300032 545096 300084 545148
rect 309968 545096 310020 545148
rect 360292 545096 360344 545148
rect 194508 543804 194560 543856
rect 223672 543804 223724 543856
rect 55036 543736 55088 543788
rect 66812 543736 66864 543788
rect 89628 543736 89680 543788
rect 270684 543736 270736 543788
rect 316592 543736 316644 543788
rect 363052 543736 363104 543788
rect 357348 543668 357400 543720
rect 582932 543668 582984 543720
rect 3424 542988 3476 543040
rect 34520 542988 34572 543040
rect 195336 542444 195388 542496
rect 218704 542444 218756 542496
rect 255964 542444 256016 542496
rect 257344 542444 257396 542496
rect 356060 542444 356112 542496
rect 357348 542444 357400 542496
rect 34520 542376 34572 542428
rect 35808 542376 35860 542428
rect 66812 542376 66864 542428
rect 91560 542376 91612 542428
rect 95976 542376 96028 542428
rect 129648 542376 129700 542428
rect 266728 542376 266780 542428
rect 67364 541832 67416 541884
rect 67548 541832 67600 541884
rect 14464 541628 14516 541680
rect 66996 541628 67048 541680
rect 67272 541628 67324 541680
rect 261760 541628 261812 541680
rect 360200 541628 360252 541680
rect 189724 541016 189776 541068
rect 230480 541016 230532 541068
rect 91928 540948 91980 541000
rect 92388 540948 92440 541000
rect 124864 540948 124916 541000
rect 258448 540948 258500 541000
rect 338304 540948 338356 541000
rect 367376 540948 367428 541000
rect 4804 540200 4856 540252
rect 65892 539656 65944 539708
rect 70400 539588 70452 539640
rect 81348 539588 81400 539640
rect 88800 539656 88852 539708
rect 195152 539656 195204 539708
rect 215852 539656 215904 539708
rect 315396 539656 315448 539708
rect 361580 539656 361632 539708
rect 250628 539588 250680 539640
rect 323584 539588 323636 539640
rect 379428 539588 379480 539640
rect 69848 539520 69900 539572
rect 85580 539520 85632 539572
rect 268384 539520 268436 539572
rect 272340 539520 272392 539572
rect 273260 539520 273312 539572
rect 275652 539520 275704 539572
rect 278044 539520 278096 539572
rect 278964 539520 279016 539572
rect 341524 539520 341576 539572
rect 343732 539520 343784 539572
rect 345388 539520 345440 539572
rect 349988 539520 350040 539572
rect 66168 538976 66220 539028
rect 72424 538976 72476 539028
rect 76748 538908 76800 538960
rect 171784 538908 171836 538960
rect 195152 538908 195204 538960
rect 7564 538840 7616 538892
rect 91100 538840 91152 538892
rect 169024 538840 169076 538892
rect 195244 538840 195296 538892
rect 195244 538296 195296 538348
rect 223212 538296 223264 538348
rect 347044 538296 347096 538348
rect 358820 538296 358872 538348
rect 226248 538228 226300 538280
rect 297180 538228 297232 538280
rect 350356 538228 350408 538280
rect 369860 538228 369912 538280
rect 88616 538160 88668 538212
rect 89628 538160 89680 538212
rect 379428 538160 379480 538212
rect 580172 538160 580224 538212
rect 12348 537548 12400 537600
rect 91192 537548 91244 537600
rect 67548 537480 67600 537532
rect 154764 537480 154816 537532
rect 197544 536868 197596 536920
rect 220820 536868 220872 536920
rect 330484 536868 330536 536920
rect 364432 536868 364484 536920
rect 178776 536800 178828 536852
rect 233884 536800 233936 536852
rect 234068 536800 234120 536852
rect 342076 536800 342128 536852
rect 378140 536800 378192 536852
rect 43444 536732 43496 536784
rect 69572 536732 69624 536784
rect 86868 536732 86920 536784
rect 130384 536732 130436 536784
rect 68652 536664 68704 536716
rect 81348 536664 81400 536716
rect 75184 536596 75236 536648
rect 85580 536596 85632 536648
rect 84292 536460 84344 536512
rect 89076 536460 89128 536512
rect 81532 535576 81584 535628
rect 83464 535576 83516 535628
rect 170496 535508 170548 535560
rect 313372 535508 313424 535560
rect 332416 535508 332468 535560
rect 358912 535508 358964 535560
rect 89628 535440 89680 535492
rect 90548 535440 90600 535492
rect 146944 535440 146996 535492
rect 293500 535440 293552 535492
rect 302332 535440 302384 535492
rect 582748 535440 582800 535492
rect 199660 535372 199712 535424
rect 202052 535372 202104 535424
rect 196624 534760 196676 534812
rect 226248 535236 226300 535288
rect 355600 535236 355652 535288
rect 425060 534760 425112 534812
rect 78312 534692 78364 534744
rect 135260 534692 135312 534744
rect 136180 534692 136232 534744
rect 151084 534692 151136 534744
rect 198740 534692 198792 534744
rect 136180 534080 136232 534132
rect 143448 534080 143500 534132
rect 41328 534012 41380 534064
rect 191104 534012 191156 534064
rect 78680 533332 78732 533384
rect 79508 533332 79560 533384
rect 143448 532652 143500 532704
rect 197452 532652 197504 532704
rect 81072 532040 81124 532092
rect 132500 532040 132552 532092
rect 133696 532040 133748 532092
rect 3424 531972 3476 532024
rect 89720 531972 89772 532024
rect 358728 531972 358780 532024
rect 359004 531972 359056 532024
rect 582932 531972 582984 532024
rect 133696 531292 133748 531344
rect 144184 531292 144236 531344
rect 79324 531224 79376 531276
rect 79968 531224 80020 531276
rect 180064 530612 180116 530664
rect 197544 530612 197596 530664
rect 64696 530544 64748 530596
rect 79324 530544 79376 530596
rect 153108 530544 153160 530596
rect 199660 530544 199712 530596
rect 50988 529864 51040 529916
rect 178684 529864 178736 529916
rect 154764 529796 154816 529848
rect 197452 529796 197504 529848
rect 358728 528572 358780 528624
rect 367284 528572 367336 528624
rect 187148 528504 187200 528556
rect 197452 528504 197504 528556
rect 358728 527144 358780 527196
rect 398840 527144 398892 527196
rect 70492 526532 70544 526584
rect 71044 526532 71096 526584
rect 71044 525784 71096 525836
rect 162216 525784 162268 525836
rect 61936 525104 61988 525156
rect 77944 525104 77996 525156
rect 50896 525036 50948 525088
rect 191104 525036 191156 525088
rect 358728 524424 358780 524476
rect 371240 524424 371292 524476
rect 34428 523676 34480 523728
rect 195336 523676 195388 523728
rect 60648 522928 60700 522980
rect 185676 522928 185728 522980
rect 155224 521636 155276 521688
rect 197452 521636 197504 521688
rect 167644 520956 167696 521008
rect 197544 520956 197596 521008
rect 63408 520888 63460 520940
rect 187056 520888 187108 520940
rect 358728 520888 358780 520940
rect 395988 520888 396040 520940
rect 395988 520276 396040 520328
rect 582380 520276 582432 520328
rect 53748 519528 53800 519580
rect 196716 519528 196768 519580
rect 358636 518916 358688 518968
rect 445760 518916 445812 518968
rect 52368 518848 52420 518900
rect 188436 518848 188488 518900
rect 52184 517488 52236 517540
rect 52368 517488 52420 517540
rect 162124 516128 162176 516180
rect 197452 516128 197504 516180
rect 358728 516128 358780 516180
rect 363604 516128 363656 516180
rect 3516 514768 3568 514820
rect 14464 514768 14516 514820
rect 162216 510552 162268 510604
rect 197452 510552 197504 510604
rect 49608 508512 49660 508564
rect 189724 508512 189776 508564
rect 134524 507084 134576 507136
rect 193956 507084 194008 507136
rect 358728 506472 358780 506524
rect 382280 506472 382332 506524
rect 358728 505112 358780 505164
rect 434720 505112 434772 505164
rect 61936 504364 61988 504416
rect 180156 504364 180208 504416
rect 173164 502936 173216 502988
rect 197452 502936 197504 502988
rect 358728 502392 358780 502444
rect 364340 502392 364392 502444
rect 187148 502324 187200 502376
rect 197452 502324 197504 502376
rect 2780 501848 2832 501900
rect 4804 501848 4856 501900
rect 144184 500896 144236 500948
rect 197452 500896 197504 500948
rect 363604 497428 363656 497480
rect 405740 497428 405792 497480
rect 358636 496748 358688 496800
rect 360200 496748 360252 496800
rect 583024 496748 583076 496800
rect 178684 495456 178736 495508
rect 197452 495456 197504 495508
rect 358728 494708 358780 494760
rect 385040 494708 385092 494760
rect 398932 494708 398984 494760
rect 412640 494708 412692 494760
rect 392216 493280 392268 493332
rect 398932 493280 398984 493332
rect 148324 492668 148376 492720
rect 197452 492668 197504 492720
rect 358728 492668 358780 492720
rect 392216 492668 392268 492720
rect 392584 492668 392636 492720
rect 187056 489880 187108 489932
rect 197452 489880 197504 489932
rect 148416 487772 148468 487824
rect 185400 487772 185452 487824
rect 184940 487160 184992 487212
rect 185400 487160 185452 487212
rect 197452 487160 197504 487212
rect 358728 487160 358780 487212
rect 380900 487160 380952 487212
rect 358176 484372 358228 484424
rect 410524 484372 410576 484424
rect 180156 483624 180208 483676
rect 197452 483624 197504 483676
rect 357900 481652 357952 481704
rect 367192 481652 367244 481704
rect 132408 480224 132460 480276
rect 197452 480224 197504 480276
rect 127624 477504 127676 477556
rect 182088 477504 182140 477556
rect 197452 477504 197504 477556
rect 357900 477504 357952 477556
rect 365720 477504 365772 477556
rect 145564 474716 145616 474768
rect 197452 474716 197504 474768
rect 358728 474716 358780 474768
rect 368572 474716 368624 474768
rect 3516 473968 3568 474020
rect 7564 473968 7616 474020
rect 15844 473968 15896 474020
rect 142804 473356 142856 473408
rect 197452 473356 197504 473408
rect 358084 473288 358136 473340
rect 360200 473288 360252 473340
rect 358728 471996 358780 472048
rect 374092 471996 374144 472048
rect 358728 470568 358780 470620
rect 371424 470568 371476 470620
rect 59084 468460 59136 468512
rect 85580 468460 85632 468512
rect 165528 467848 165580 467900
rect 197452 467848 197504 467900
rect 67824 467780 67876 467832
rect 74540 467780 74592 467832
rect 156604 465672 156656 465724
rect 197452 465672 197504 465724
rect 130568 465060 130620 465112
rect 156604 465060 156656 465112
rect 358728 465060 358780 465112
rect 379520 465060 379572 465112
rect 583300 465060 583352 465112
rect 106188 464312 106240 464364
rect 120816 464312 120868 464364
rect 65984 462952 66036 463004
rect 91560 462952 91612 463004
rect 107016 462952 107068 463004
rect 122932 462952 122984 463004
rect 2780 462544 2832 462596
rect 4804 462544 4856 462596
rect 187240 462340 187292 462392
rect 197452 462340 197504 462392
rect 358636 462340 358688 462392
rect 360384 462340 360436 462392
rect 63224 461592 63276 461644
rect 78772 461592 78824 461644
rect 76012 461456 76064 461508
rect 76564 461456 76616 461508
rect 76564 460912 76616 460964
rect 179420 460912 179472 460964
rect 191748 460844 191800 460896
rect 197452 460844 197504 460896
rect 52368 460164 52420 460216
rect 90456 460164 90508 460216
rect 166264 460164 166316 460216
rect 191748 460164 191800 460216
rect 372988 460164 373040 460216
rect 582564 460164 582616 460216
rect 56508 459552 56560 459604
rect 67732 459552 67784 459604
rect 91100 459552 91152 459604
rect 91560 459552 91612 459604
rect 159364 459552 159416 459604
rect 358728 459552 358780 459604
rect 372712 459552 372764 459604
rect 372988 459552 373040 459604
rect 67732 458804 67784 458856
rect 81440 458804 81492 458856
rect 91744 458804 91796 458856
rect 120632 458804 120684 458856
rect 55128 457444 55180 457496
rect 87604 457444 87656 457496
rect 115204 457444 115256 457496
rect 126980 457444 127032 457496
rect 69020 456764 69072 456816
rect 69848 456764 69900 456816
rect 157984 456764 158036 456816
rect 62028 456016 62080 456068
rect 78680 456016 78732 456068
rect 108304 456016 108356 456068
rect 127716 456016 127768 456068
rect 88340 455404 88392 455456
rect 88984 455404 89036 455456
rect 125600 455404 125652 455456
rect 191288 455404 191340 455456
rect 197452 455404 197504 455456
rect 358728 455404 358780 455456
rect 376760 455404 376812 455456
rect 582380 455404 582432 455456
rect 14464 455336 14516 455388
rect 111800 455336 111852 455388
rect 77300 455268 77352 455320
rect 77944 455268 77996 455320
rect 63316 454656 63368 454708
rect 67640 454656 67692 454708
rect 111800 454656 111852 454708
rect 183560 454656 183612 454708
rect 184296 454656 184348 454708
rect 77300 454112 77352 454164
rect 132592 454044 132644 454096
rect 193956 453500 194008 453552
rect 197360 453500 197412 453552
rect 61752 453364 61804 453416
rect 75920 453364 75972 453416
rect 57704 453296 57756 453348
rect 72424 453296 72476 453348
rect 112444 453296 112496 453348
rect 123024 453296 123076 453348
rect 125508 453296 125560 453348
rect 151084 453296 151136 453348
rect 72700 452616 72752 452668
rect 125508 452616 125560 452668
rect 358728 452616 358780 452668
rect 377404 452616 377456 452668
rect 66168 451936 66220 451988
rect 75184 451936 75236 451988
rect 116676 451936 116728 451988
rect 124312 451936 124364 451988
rect 3424 451868 3476 451920
rect 121460 451868 121512 451920
rect 95884 451188 95936 451240
rect 127624 451188 127676 451240
rect 4804 450508 4856 450560
rect 68100 450508 68152 450560
rect 50804 449964 50856 450016
rect 74540 449964 74592 450016
rect 74816 449964 74868 450016
rect 68100 449896 68152 449948
rect 68560 449896 68612 449948
rect 103520 449896 103572 449948
rect 103704 449896 103756 449948
rect 358728 449896 358780 449948
rect 374000 449896 374052 449948
rect 39948 449828 40000 449880
rect 72700 449828 72752 449880
rect 106924 449828 106976 449880
rect 129004 449828 129056 449880
rect 50896 449148 50948 449200
rect 80888 449148 80940 449200
rect 100668 449148 100720 449200
rect 108304 449148 108356 449200
rect 371516 449148 371568 449200
rect 582656 449148 582708 449200
rect 116584 448604 116636 448656
rect 120724 448604 120776 448656
rect 3148 448536 3200 448588
rect 25504 448536 25556 448588
rect 72700 448536 72752 448588
rect 73160 448536 73212 448588
rect 190276 448536 190328 448588
rect 197360 448536 197412 448588
rect 358728 448536 358780 448588
rect 371332 448536 371384 448588
rect 371516 448536 371568 448588
rect 94504 448468 94556 448520
rect 187240 448468 187292 448520
rect 64604 447788 64656 447840
rect 71044 447788 71096 447840
rect 11704 447108 11756 447160
rect 12348 447108 12400 447160
rect 125692 447108 125744 447160
rect 109684 447040 109736 447092
rect 146944 447040 146996 447092
rect 65984 446360 66036 446412
rect 73252 446360 73304 446412
rect 98644 445816 98696 445868
rect 100484 445816 100536 445868
rect 102232 445816 102284 445868
rect 7564 445748 7616 445800
rect 118700 445748 118752 445800
rect 174636 445748 174688 445800
rect 197360 445748 197412 445800
rect 358728 445748 358780 445800
rect 369952 445748 370004 445800
rect 67640 445680 67692 445732
rect 68744 445680 68796 445732
rect 119344 444524 119396 444576
rect 120908 444524 120960 444576
rect 53564 444456 53616 444508
rect 85580 444456 85632 444508
rect 100760 444456 100812 444508
rect 127624 444456 127676 444508
rect 68928 444388 68980 444440
rect 146944 444388 146996 444440
rect 166908 443708 166960 443760
rect 197360 443708 197412 443760
rect 124128 443640 124180 443692
rect 126980 443640 127032 443692
rect 169760 443640 169812 443692
rect 192576 443640 192628 443692
rect 358728 442960 358780 443012
rect 361672 442960 361724 443012
rect 48136 442892 48188 442944
rect 67732 442892 67784 442944
rect 124128 441600 124180 441652
rect 140044 441600 140096 441652
rect 192668 441396 192720 441448
rect 197728 441396 197780 441448
rect 60464 440240 60516 440292
rect 66904 440240 66956 440292
rect 121460 440172 121512 440224
rect 130568 440172 130620 440224
rect 358728 438880 358780 438932
rect 376024 438880 376076 438932
rect 63316 437520 63368 437572
rect 64788 437520 64840 437572
rect 66904 437520 66956 437572
rect 124128 437452 124180 437504
rect 128360 437452 128412 437504
rect 129004 437452 129056 437504
rect 155776 437384 155828 437436
rect 162124 437384 162176 437436
rect 162768 436092 162820 436144
rect 197360 436092 197412 436144
rect 358728 436092 358780 436144
rect 363144 436092 363196 436144
rect 53656 436024 53708 436076
rect 57888 436024 57940 436076
rect 155316 436024 155368 436076
rect 156604 436024 156656 436076
rect 57888 434732 57940 434784
rect 66904 434732 66956 434784
rect 120724 434732 120776 434784
rect 128360 434732 128412 434784
rect 165620 434664 165672 434716
rect 166264 434664 166316 434716
rect 127716 433984 127768 434036
rect 165620 433984 165672 434036
rect 46848 433304 46900 433356
rect 179328 433304 179380 433356
rect 197360 433304 197412 433356
rect 358728 433304 358780 433356
rect 365812 433304 365864 433356
rect 55864 433236 55916 433288
rect 66812 433236 66864 433288
rect 124128 433236 124180 433288
rect 127716 433236 127768 433288
rect 52276 431196 52328 431248
rect 65892 431196 65944 431248
rect 66536 431196 66588 431248
rect 124128 430584 124180 430636
rect 172428 430584 172480 430636
rect 173256 430584 173308 430636
rect 36728 429088 36780 429140
rect 37188 429088 37240 429140
rect 66720 429088 66772 429140
rect 121460 429088 121512 429140
rect 177304 429088 177356 429140
rect 14464 428408 14516 428460
rect 36728 428408 36780 428460
rect 192576 427796 192628 427848
rect 197360 427796 197412 427848
rect 358728 427796 358780 427848
rect 363236 427796 363288 427848
rect 137284 426436 137336 426488
rect 197360 426436 197412 426488
rect 358728 426436 358780 426488
rect 372620 426436 372672 426488
rect 41328 425688 41380 425740
rect 59084 425688 59136 425740
rect 59084 425076 59136 425128
rect 66260 425076 66312 425128
rect 61844 423648 61896 423700
rect 66076 423648 66128 423700
rect 167736 423648 167788 423700
rect 197360 423648 197412 423700
rect 3424 423580 3476 423632
rect 11704 423580 11756 423632
rect 124128 422220 124180 422272
rect 136640 422220 136692 422272
rect 52276 421540 52328 421592
rect 59176 421540 59228 421592
rect 66260 421540 66312 421592
rect 136640 421540 136692 421592
rect 162676 421540 162728 421592
rect 178776 421540 178828 421592
rect 123024 420860 123076 420912
rect 170496 420860 170548 420912
rect 43996 418752 44048 418804
rect 59176 418752 59228 418804
rect 176200 418140 176252 418192
rect 197360 418140 197412 418192
rect 358728 418140 358780 418192
rect 361764 418140 361816 418192
rect 59176 416780 59228 416832
rect 66904 416780 66956 416832
rect 358728 416780 358780 416832
rect 368480 416780 368532 416832
rect 57796 416032 57848 416084
rect 66260 416032 66312 416084
rect 57796 414672 57848 414724
rect 66260 414672 66312 414724
rect 124128 414672 124180 414724
rect 138020 414672 138072 414724
rect 181444 413992 181496 414044
rect 197360 413992 197412 414044
rect 358728 413992 358780 414044
rect 370044 413992 370096 414044
rect 122840 413244 122892 413296
rect 133880 413244 133932 413296
rect 161388 411272 161440 411324
rect 197360 411272 197412 411324
rect 358728 411272 358780 411324
rect 378232 411272 378284 411324
rect 121184 409844 121236 409896
rect 151084 409844 151136 409896
rect 130384 409776 130436 409828
rect 197360 409776 197412 409828
rect 124128 408416 124180 408468
rect 133788 408416 133840 408468
rect 134616 408416 134668 408468
rect 60648 407124 60700 407176
rect 66352 407124 66404 407176
rect 124312 405968 124364 406020
rect 124864 405968 124916 406020
rect 59268 405764 59320 405816
rect 63132 405764 63184 405816
rect 66812 405764 66864 405816
rect 133144 405696 133196 405748
rect 197360 405696 197412 405748
rect 358728 405696 358780 405748
rect 364524 405696 364576 405748
rect 189816 404336 189868 404388
rect 197360 404336 197412 404388
rect 122932 403520 122984 403572
rect 125048 403520 125100 403572
rect 48136 402908 48188 402960
rect 52184 402908 52236 402960
rect 52184 402228 52236 402280
rect 66628 403112 66680 403164
rect 358728 402976 358780 403028
rect 365904 402976 365956 403028
rect 122104 401616 122156 401668
rect 122932 401616 122984 401668
rect 358728 401616 358780 401668
rect 416780 401616 416832 401668
rect 166908 400936 166960 400988
rect 178040 400936 178092 400988
rect 50896 400868 50948 400920
rect 66812 400868 66864 400920
rect 123944 400868 123996 400920
rect 193956 400868 194008 400920
rect 55036 399440 55088 399492
rect 66812 399440 66864 399492
rect 124128 399440 124180 399492
rect 125692 399440 125744 399492
rect 192668 399440 192720 399492
rect 194048 398828 194100 398880
rect 197360 398828 197412 398880
rect 358636 398828 358688 398880
rect 361856 398828 361908 398880
rect 3516 397536 3568 397588
rect 7564 397536 7616 397588
rect 124128 396924 124180 396976
rect 129740 396924 129792 396976
rect 35808 396720 35860 396772
rect 66996 396720 67048 396772
rect 140044 396720 140096 396772
rect 164884 396720 164936 396772
rect 59176 395972 59228 396024
rect 66076 395972 66128 396024
rect 125508 395292 125560 395344
rect 148416 395292 148468 395344
rect 171048 394680 171100 394732
rect 197360 394680 197412 394732
rect 120724 393932 120776 393984
rect 120908 393932 120960 393984
rect 129740 393932 129792 393984
rect 177396 393932 177448 393984
rect 356336 393320 356388 393372
rect 393320 393320 393372 393372
rect 48228 393252 48280 393304
rect 65800 393252 65852 393304
rect 123760 392368 123812 392420
rect 131764 392368 131816 392420
rect 130384 391960 130436 392012
rect 180156 391960 180208 392012
rect 73068 391008 73120 391060
rect 145564 391212 145616 391264
rect 72056 390532 72108 390584
rect 73068 390532 73120 390584
rect 131120 390532 131172 390584
rect 132408 390532 132460 390584
rect 168380 390532 168432 390584
rect 66076 390464 66128 390516
rect 197360 390464 197412 390516
rect 65984 389172 66036 389224
rect 77852 389172 77904 389224
rect 131120 389172 131172 389224
rect 64604 389104 64656 389156
rect 73160 389104 73212 389156
rect 115204 389104 115256 389156
rect 120448 389104 120500 389156
rect 96252 388492 96304 388544
rect 188804 388492 188856 388544
rect 194048 388492 194100 388544
rect 15844 388424 15896 388476
rect 110328 388424 110380 388476
rect 88524 387812 88576 387864
rect 90364 387812 90416 387864
rect 110328 387812 110380 387864
rect 111432 387812 111484 387864
rect 123484 387812 123536 387864
rect 162124 387812 162176 387864
rect 64788 387064 64840 387116
rect 68744 387064 68796 387116
rect 113088 387064 113140 387116
rect 120908 387064 120960 387116
rect 7564 386384 7616 386436
rect 117320 386384 117372 386436
rect 117964 386384 118016 386436
rect 191196 386384 191248 386436
rect 197360 386384 197412 386436
rect 62028 386316 62080 386368
rect 86960 386316 87012 386368
rect 117596 385636 117648 385688
rect 191380 385636 191432 385688
rect 97264 385024 97316 385076
rect 197360 385024 197412 385076
rect 57704 384956 57756 385008
rect 82084 384956 82136 385008
rect 86868 384344 86920 384396
rect 100484 384344 100536 384396
rect 184388 384344 184440 384396
rect 63316 384276 63368 384328
rect 173808 384276 173860 384328
rect 193128 383664 193180 383716
rect 196716 383664 196768 383716
rect 357900 383664 357952 383716
rect 400864 383664 400916 383716
rect 77944 382916 77996 382968
rect 148324 382916 148376 382968
rect 157984 382916 158036 382968
rect 177304 382916 177356 382968
rect 147680 382304 147732 382356
rect 157340 382304 157392 382356
rect 119988 382236 120040 382288
rect 185584 382236 185636 382288
rect 3608 381488 3660 381540
rect 105544 381488 105596 381540
rect 110328 381488 110380 381540
rect 157984 381488 158036 381540
rect 157340 380944 157392 380996
rect 163412 380944 163464 380996
rect 67548 380876 67600 380928
rect 195520 380876 195572 380928
rect 44088 380808 44140 380860
rect 75920 380808 75972 380860
rect 76564 380808 76616 380860
rect 75184 380196 75236 380248
rect 113180 380196 113232 380248
rect 103336 380128 103388 380180
rect 152464 380128 152516 380180
rect 177396 380128 177448 380180
rect 194416 380128 194468 380180
rect 197360 380128 197412 380180
rect 129832 379584 129884 379636
rect 195336 379584 195388 379636
rect 357900 379516 357952 379568
rect 360476 379516 360528 379568
rect 117964 378768 118016 378820
rect 159456 378768 159508 378820
rect 60556 378156 60608 378208
rect 190460 378156 190512 378208
rect 191288 378156 191340 378208
rect 70308 377476 70360 377528
rect 167000 377476 167052 377528
rect 11704 377408 11756 377460
rect 122840 377408 122892 377460
rect 190276 377408 190328 377460
rect 203616 377408 203668 377460
rect 354128 377408 354180 377460
rect 360292 377408 360344 377460
rect 153844 376728 153896 376780
rect 185676 376728 185728 376780
rect 66904 376660 66956 376712
rect 67364 376660 67416 376712
rect 345756 376048 345808 376100
rect 357716 376048 357768 376100
rect 60648 375980 60700 376032
rect 71688 375980 71740 376032
rect 172428 375980 172480 376032
rect 184296 375980 184348 376032
rect 198924 375980 198976 376032
rect 204352 375980 204404 376032
rect 248052 375980 248104 376032
rect 376116 375980 376168 376032
rect 197084 375640 197136 375692
rect 200304 375640 200356 375692
rect 66904 375368 66956 375420
rect 195888 375368 195940 375420
rect 191380 375300 191432 375352
rect 205824 375300 205876 375352
rect 206652 375300 206704 375352
rect 207020 375300 207072 375352
rect 208308 375300 208360 375352
rect 258724 375300 258776 375352
rect 261484 375300 261536 375352
rect 269856 375300 269908 375352
rect 274732 375300 274784 375352
rect 279516 375300 279568 375352
rect 280160 375300 280212 375352
rect 311900 375300 311952 375352
rect 312820 375300 312872 375352
rect 317972 375300 318024 375352
rect 320180 375300 320232 375352
rect 351184 375300 351236 375352
rect 354404 375300 354456 375352
rect 199384 375232 199436 375284
rect 199936 375232 199988 375284
rect 278228 375096 278280 375148
rect 279700 375096 279752 375148
rect 112444 374688 112496 374740
rect 130384 374688 130436 374740
rect 233884 374688 233936 374740
rect 244740 374756 244792 374808
rect 242164 374688 242216 374740
rect 243084 374688 243136 374740
rect 250444 374688 250496 374740
rect 251364 374688 251416 374740
rect 338764 374688 338816 374740
rect 347780 374688 347832 374740
rect 59084 374620 59136 374672
rect 162860 374620 162912 374672
rect 163412 374620 163464 374672
rect 186412 374620 186464 374672
rect 199844 374620 199896 374672
rect 207112 374620 207164 374672
rect 209044 374620 209096 374672
rect 213276 374620 213328 374672
rect 217324 374620 217376 374672
rect 239772 374620 239824 374672
rect 298744 374620 298796 374672
rect 316132 374620 316184 374672
rect 342168 374620 342220 374672
rect 352748 374620 352800 374672
rect 267648 374076 267700 374128
rect 269764 374076 269816 374128
rect 131764 374008 131816 374060
rect 189724 374008 189776 374060
rect 213276 374008 213328 374060
rect 219900 374008 219952 374060
rect 267004 374008 267056 374060
rect 268108 374008 268160 374060
rect 271144 374008 271196 374060
rect 278044 374008 278096 374060
rect 290464 374008 290516 374060
rect 297916 374008 297968 374060
rect 308404 374008 308456 374060
rect 309876 374008 309928 374060
rect 325608 374008 325660 374060
rect 327908 374008 327960 374060
rect 197176 373328 197228 373380
rect 205640 373328 205692 373380
rect 349804 373328 349856 373380
rect 360476 373328 360528 373380
rect 84108 373260 84160 373312
rect 115204 373260 115256 373312
rect 188804 373260 188856 373312
rect 215944 373260 215996 373312
rect 352656 373260 352708 373312
rect 365904 373260 365956 373312
rect 124956 372648 125008 372700
rect 172060 372648 172112 372700
rect 53564 372580 53616 372632
rect 196808 372580 196860 372632
rect 52092 372512 52144 372564
rect 370044 372512 370096 372564
rect 89628 371832 89680 371884
rect 356336 371832 356388 371884
rect 2964 371356 3016 371408
rect 4804 371356 4856 371408
rect 125048 371152 125100 371204
rect 129740 371152 129792 371204
rect 146208 370540 146260 370592
rect 207020 370540 207072 370592
rect 347044 370540 347096 370592
rect 365812 370540 365864 370592
rect 185584 370472 185636 370524
rect 253940 370472 253992 370524
rect 262864 370472 262916 370524
rect 357624 370472 357676 370524
rect 207020 370268 207072 370320
rect 208308 370268 208360 370320
rect 129188 369860 129240 369912
rect 173256 369860 173308 369912
rect 252560 369860 252612 369912
rect 253296 369860 253348 369912
rect 302884 369860 302936 369912
rect 25504 369792 25556 369844
rect 26148 369792 26200 369844
rect 131764 369792 131816 369844
rect 182088 369180 182140 369232
rect 191288 369180 191340 369232
rect 195244 369180 195296 369232
rect 256056 369180 256108 369232
rect 71596 369112 71648 369164
rect 73160 369112 73212 369164
rect 76564 369112 76616 369164
rect 155224 369112 155276 369164
rect 166908 369112 166960 369164
rect 241428 369112 241480 369164
rect 253204 369112 253256 369164
rect 255964 369112 256016 369164
rect 309784 369112 309836 369164
rect 311900 369112 311952 369164
rect 318064 369112 318116 369164
rect 359096 369112 359148 369164
rect 144828 368500 144880 368552
rect 181628 368500 181680 368552
rect 186412 368432 186464 368484
rect 189908 368432 189960 368484
rect 147772 368296 147824 368348
rect 148416 368296 148468 368348
rect 67732 367820 67784 367872
rect 126244 367820 126296 367872
rect 73804 367752 73856 367804
rect 153844 367752 153896 367804
rect 190368 367752 190420 367804
rect 213184 367752 213236 367804
rect 147772 367072 147824 367124
rect 194600 367072 194652 367124
rect 234620 366800 234672 366852
rect 235356 366800 235408 366852
rect 331864 366392 331916 366444
rect 356244 366392 356296 366444
rect 56508 366324 56560 366376
rect 85488 366324 85540 366376
rect 316684 366324 316736 366376
rect 336740 366324 336792 366376
rect 340880 366324 340932 366376
rect 412640 366324 412692 366376
rect 114652 365780 114704 365832
rect 182916 365780 182968 365832
rect 203524 365780 203576 365832
rect 209780 365780 209832 365832
rect 118516 365712 118568 365764
rect 120264 365712 120316 365764
rect 235356 365712 235408 365764
rect 61660 364964 61712 365016
rect 74540 364964 74592 365016
rect 266360 364964 266412 365016
rect 274640 364964 274692 365016
rect 297364 364964 297416 365016
rect 331220 364964 331272 365016
rect 340236 364964 340288 365016
rect 367376 364964 367428 365016
rect 201592 364692 201644 364744
rect 202144 364692 202196 364744
rect 72424 364420 72476 364472
rect 201592 364420 201644 364472
rect 124128 364352 124180 364404
rect 265624 364352 265676 364404
rect 177948 363740 178000 363792
rect 204904 363740 204956 363792
rect 189908 363672 189960 363724
rect 195428 363672 195480 363724
rect 133880 363604 133932 363656
rect 177948 363604 178000 363656
rect 202236 363604 202288 363656
rect 235264 363604 235316 363656
rect 317328 363604 317380 363656
rect 360384 363604 360436 363656
rect 77208 362924 77260 362976
rect 171784 362924 171836 362976
rect 171968 362924 172020 362976
rect 195520 362244 195572 362296
rect 202236 362244 202288 362296
rect 61844 362176 61896 362228
rect 131028 362176 131080 362228
rect 162676 362176 162728 362228
rect 164240 362176 164292 362228
rect 136548 361564 136600 361616
rect 231860 361564 231912 361616
rect 232596 361564 232648 361616
rect 167000 361496 167052 361548
rect 309140 361496 309192 361548
rect 91008 360884 91060 360936
rect 114652 360884 114704 360936
rect 322204 360884 322256 360936
rect 361764 360884 361816 360936
rect 54944 360816 54996 360868
rect 112444 360816 112496 360868
rect 345020 360816 345072 360868
rect 418804 360816 418856 360868
rect 166356 360272 166408 360324
rect 167000 360272 167052 360324
rect 111800 360204 111852 360256
rect 113088 360204 113140 360256
rect 264336 360204 264388 360256
rect 195336 359524 195388 359576
rect 234528 359524 234580 359576
rect 126980 359456 127032 359508
rect 127624 359456 127676 359508
rect 259552 359456 259604 359508
rect 282184 359456 282236 359508
rect 368572 359456 368624 359508
rect 104900 358776 104952 358828
rect 186964 358776 187016 358828
rect 3424 358572 3476 358624
rect 7564 358572 7616 358624
rect 207112 358504 207164 358556
rect 207664 358504 207716 358556
rect 270408 358028 270460 358080
rect 319444 358028 319496 358080
rect 358176 358028 358228 358080
rect 374092 358028 374144 358080
rect 90364 357484 90416 357536
rect 207664 357484 207716 357536
rect 130384 357416 130436 357468
rect 131120 357416 131172 357468
rect 269764 357416 269816 357468
rect 270408 357416 270460 357468
rect 234528 357348 234580 357400
rect 354128 357348 354180 357400
rect 63132 356736 63184 356788
rect 108304 356736 108356 356788
rect 81624 356668 81676 356720
rect 82084 356668 82136 356720
rect 258724 356668 258776 356720
rect 141516 356056 141568 356108
rect 170496 356056 170548 356108
rect 170588 356056 170640 356108
rect 171048 356056 171100 356108
rect 226984 356056 227036 356108
rect 3424 355376 3476 355428
rect 92480 355376 92532 355428
rect 196808 355376 196860 355428
rect 215392 355376 215444 355428
rect 87604 355308 87656 355360
rect 122288 355308 122340 355360
rect 174820 355308 174872 355360
rect 181536 355308 181588 355360
rect 211160 355308 211212 355360
rect 356704 355308 356756 355360
rect 382280 355308 382332 355360
rect 192484 354968 192536 355020
rect 192760 354968 192812 355020
rect 93768 354696 93820 354748
rect 192484 354696 192536 354748
rect 265624 354628 265676 354680
rect 353944 354628 353996 354680
rect 171784 353948 171836 354000
rect 222200 353948 222252 354000
rect 101864 353336 101916 353388
rect 170588 353336 170640 353388
rect 124864 353268 124916 353320
rect 127072 353268 127124 353320
rect 128176 353268 128228 353320
rect 133144 353268 133196 353320
rect 205732 353268 205784 353320
rect 206284 353268 206336 353320
rect 125600 353200 125652 353252
rect 233884 353200 233936 353252
rect 77392 352588 77444 352640
rect 94504 352588 94556 352640
rect 81348 352520 81400 352572
rect 125600 352520 125652 352572
rect 270408 352520 270460 352572
rect 363052 352520 363104 352572
rect 110328 351908 110380 351960
rect 196624 351908 196676 351960
rect 158076 351840 158128 351892
rect 158628 351840 158680 351892
rect 364524 351840 364576 351892
rect 85488 351160 85540 351212
rect 94044 351160 94096 351212
rect 111156 351160 111208 351212
rect 138020 351160 138072 351212
rect 146944 351092 146996 351144
rect 147588 351092 147640 351144
rect 167828 351160 167880 351212
rect 84384 350548 84436 350600
rect 85396 350548 85448 350600
rect 157340 350548 157392 350600
rect 97908 349800 97960 349852
rect 132592 349800 132644 349852
rect 188528 349800 188580 349852
rect 197268 349800 197320 349852
rect 358084 349800 358136 349852
rect 89536 349120 89588 349172
rect 193864 349120 193916 349172
rect 110420 349052 110472 349104
rect 137284 349052 137336 349104
rect 223580 348984 223632 349036
rect 224224 348984 224276 349036
rect 235356 348440 235408 348492
rect 251824 348440 251876 348492
rect 79968 348372 80020 348424
rect 110972 348372 111024 348424
rect 140688 348372 140740 348424
rect 199016 348372 199068 348424
rect 242164 348372 242216 348424
rect 272524 348372 272576 348424
rect 358912 348372 358964 348424
rect 106924 347760 106976 347812
rect 121460 347760 121512 347812
rect 151084 347760 151136 347812
rect 224224 347760 224276 347812
rect 205640 347692 205692 347744
rect 206376 347692 206428 347744
rect 169576 347012 169628 347064
rect 322204 347012 322256 347064
rect 338856 347012 338908 347064
rect 356796 347012 356848 347064
rect 66076 346468 66128 346520
rect 150440 346468 150492 346520
rect 64604 346400 64656 346452
rect 66904 346400 66956 346452
rect 67272 346400 67324 346452
rect 99104 346400 99156 346452
rect 206376 346400 206428 346452
rect 157340 346332 157392 346384
rect 181536 346332 181588 346384
rect 350448 346332 350500 346384
rect 352564 346332 352616 346384
rect 99288 345652 99340 345704
rect 158076 345652 158128 345704
rect 189724 345652 189776 345704
rect 209780 345652 209832 345704
rect 249064 345652 249116 345704
rect 269856 345652 269908 345704
rect 122840 345040 122892 345092
rect 123484 345040 123536 345092
rect 249064 345040 249116 345092
rect 150440 344972 150492 345024
rect 198004 344972 198056 345024
rect 286232 344292 286284 344344
rect 420920 344292 420972 344344
rect 115848 343612 115900 343664
rect 125048 343612 125100 343664
rect 137284 343612 137336 343664
rect 156788 343612 156840 343664
rect 157984 343612 158036 343664
rect 159548 343612 159600 343664
rect 186228 343612 186280 343664
rect 190460 343612 190512 343664
rect 264336 343544 264388 343596
rect 343640 343544 343692 343596
rect 71688 342932 71740 342984
rect 87144 342932 87196 342984
rect 96436 342932 96488 342984
rect 111156 342932 111208 342984
rect 60372 342864 60424 342916
rect 97264 342864 97316 342916
rect 195520 342864 195572 342916
rect 261484 342864 261536 342916
rect 264336 342796 264388 342848
rect 264888 342796 264940 342848
rect 115756 342320 115808 342372
rect 183192 342320 183244 342372
rect 111708 342252 111760 342304
rect 115848 342252 115900 342304
rect 144184 342252 144236 342304
rect 220084 342252 220136 342304
rect 69756 341504 69808 341556
rect 141516 341504 141568 341556
rect 153844 341504 153896 341556
rect 163596 341504 163648 341556
rect 188436 341504 188488 341556
rect 211804 341504 211856 341556
rect 142344 340960 142396 341012
rect 154028 340960 154080 341012
rect 85580 340892 85632 340944
rect 252560 340892 252612 340944
rect 251916 340824 251968 340876
rect 259092 340824 259144 340876
rect 53656 340144 53708 340196
rect 86960 340144 87012 340196
rect 107476 340144 107528 340196
rect 133144 340144 133196 340196
rect 224224 340144 224276 340196
rect 243544 340144 243596 340196
rect 258816 340144 258868 340196
rect 259092 340144 259144 340196
rect 349160 340144 349212 340196
rect 134248 339532 134300 339584
rect 213276 339532 213328 339584
rect 67824 339464 67876 339516
rect 229744 339464 229796 339516
rect 237932 339396 237984 339448
rect 240140 339396 240192 339448
rect 84108 338716 84160 338768
rect 104164 338716 104216 338768
rect 283564 338716 283616 338768
rect 379520 338716 379572 338768
rect 100576 338172 100628 338224
rect 154488 338172 154540 338224
rect 155316 338172 155368 338224
rect 237932 338172 237984 338224
rect 238668 338172 238720 338224
rect 103704 338104 103756 338156
rect 252652 338104 252704 338156
rect 151084 338036 151136 338088
rect 152648 338036 152700 338088
rect 176108 337560 176160 337612
rect 183008 337560 183060 337612
rect 209136 337424 209188 337476
rect 264980 337424 265032 337476
rect 183100 337356 183152 337408
rect 202880 337356 202932 337408
rect 245016 337356 245068 337408
rect 367284 337356 367336 337408
rect 114468 336812 114520 336864
rect 174544 336812 174596 336864
rect 64696 336744 64748 336796
rect 224224 336744 224276 336796
rect 67732 336676 67784 336728
rect 71780 336676 71832 336728
rect 76656 336064 76708 336116
rect 87604 336064 87656 336116
rect 81072 335996 81124 336048
rect 93124 335996 93176 336048
rect 150532 335996 150584 336048
rect 199476 335996 199528 336048
rect 113088 335384 113140 335436
rect 150440 335384 150492 335436
rect 94136 335316 94188 335368
rect 248512 335316 248564 335368
rect 125048 335248 125100 335300
rect 144184 335248 144236 335300
rect 251916 334636 251968 334688
rect 348424 334636 348476 334688
rect 64512 334568 64564 334620
rect 106924 334568 106976 334620
rect 188436 334568 188488 334620
rect 313280 334568 313332 334620
rect 52184 334024 52236 334076
rect 125508 334024 125560 334076
rect 145288 334024 145340 334076
rect 163320 334024 163372 334076
rect 116768 333956 116820 334008
rect 192668 333956 192720 334008
rect 66168 333208 66220 333260
rect 124220 333208 124272 333260
rect 150440 333208 150492 333260
rect 228364 333208 228416 333260
rect 60464 332596 60516 332648
rect 140780 332596 140832 332648
rect 150348 332596 150400 332648
rect 159364 332596 159416 332648
rect 198832 332528 198884 332580
rect 202328 332528 202380 332580
rect 202788 332528 202840 332580
rect 335360 332528 335412 332580
rect 202236 332324 202288 332376
rect 202788 332324 202840 332376
rect 72976 332120 73028 332172
rect 73804 332120 73856 332172
rect 75828 332120 75880 332172
rect 76564 332120 76616 332172
rect 90456 332120 90508 332172
rect 90916 332120 90968 332172
rect 91836 332120 91888 332172
rect 93216 332120 93268 332172
rect 100024 332120 100076 332172
rect 100576 332120 100628 332172
rect 110880 332120 110932 332172
rect 111616 332120 111668 332172
rect 118884 331984 118936 332036
rect 119896 331984 119948 332036
rect 129280 331916 129332 331968
rect 145288 331916 145340 331968
rect 167828 331916 167880 331968
rect 191104 331916 191156 331968
rect 103244 331848 103296 331900
rect 129096 331848 129148 331900
rect 140780 331848 140832 331900
rect 157340 331848 157392 331900
rect 187240 331848 187292 331900
rect 249800 331848 249852 331900
rect 70676 331780 70728 331832
rect 72424 331780 72476 331832
rect 77668 331780 77720 331832
rect 77944 331780 77996 331832
rect 97080 331712 97132 331764
rect 97908 331712 97960 331764
rect 88248 331576 88300 331628
rect 90364 331576 90416 331628
rect 80336 331508 80388 331560
rect 81348 331508 81400 331560
rect 95608 331508 95660 331560
rect 96528 331508 96580 331560
rect 88984 331440 89036 331492
rect 89628 331440 89680 331492
rect 98552 331440 98604 331492
rect 99196 331440 99248 331492
rect 123300 331440 123352 331492
rect 124128 331440 124180 331492
rect 129924 331440 129976 331492
rect 130384 331440 130436 331492
rect 131488 331440 131540 331492
rect 132408 331440 132460 331492
rect 132776 331440 132828 331492
rect 133696 331440 133748 331492
rect 135720 331440 135772 331492
rect 141424 331440 141476 331492
rect 50988 331304 51040 331356
rect 69388 331304 69440 331356
rect 109408 331304 109460 331356
rect 110328 331304 110380 331356
rect 138664 331304 138716 331356
rect 139308 331304 139360 331356
rect 143816 331304 143868 331356
rect 144828 331304 144880 331356
rect 52276 331236 52328 331288
rect 77668 331236 77720 331288
rect 126888 331236 126940 331288
rect 129740 331236 129792 331288
rect 146760 331236 146812 331288
rect 176108 331236 176160 331288
rect 195428 331236 195480 331288
rect 198740 331236 198792 331288
rect 50528 331168 50580 331220
rect 50804 331168 50856 331220
rect 136548 331168 136600 331220
rect 153200 330556 153252 330608
rect 155960 330556 156012 330608
rect 157340 330556 157392 330608
rect 167920 330556 167972 330608
rect 33784 330488 33836 330540
rect 50528 330488 50580 330540
rect 125508 330488 125560 330540
rect 159456 330488 159508 330540
rect 160100 330488 160152 330540
rect 162124 330488 162176 330540
rect 225604 330488 225656 330540
rect 153200 330420 153252 330472
rect 151176 329808 151228 329860
rect 157984 329808 158036 329860
rect 70032 329740 70084 329792
rect 71044 329740 71096 329792
rect 153200 329740 153252 329792
rect 198096 329740 198148 329792
rect 67272 329672 67324 329724
rect 69756 329672 69808 329724
rect 20 328448 72 328500
rect 94228 329060 94280 329112
rect 115388 329060 115440 329112
rect 132224 329060 132276 329112
rect 145380 329060 145432 329112
rect 152188 329060 152240 329112
rect 155868 329060 155920 329112
rect 156328 329060 156380 329112
rect 157064 329060 157116 329112
rect 164792 329060 164844 329112
rect 182180 329060 182232 329112
rect 186964 329060 187016 329112
rect 220176 329060 220228 329112
rect 226984 329060 227036 329112
rect 322204 329060 322256 329112
rect 156880 328584 156932 328636
rect 40684 327700 40736 327752
rect 156696 328448 156748 328500
rect 159456 328448 159508 328500
rect 159548 328448 159600 328500
rect 164976 328448 165028 328500
rect 156880 328312 156932 328364
rect 156696 328244 156748 328296
rect 215116 327768 215168 327820
rect 292580 327768 292632 327820
rect 163320 327700 163372 327752
rect 186964 327700 187016 327752
rect 272616 327700 272668 327752
rect 362960 327700 363012 327752
rect 156696 327088 156748 327140
rect 236736 327088 236788 327140
rect 240048 327088 240100 327140
rect 272616 327088 272668 327140
rect 180064 326408 180116 326460
rect 206468 326408 206520 326460
rect 157064 326340 157116 326392
rect 195244 326340 195296 326392
rect 214564 326340 214616 326392
rect 344284 326340 344336 326392
rect 48228 325660 48280 325712
rect 66260 325660 66312 325712
rect 158720 325660 158772 325712
rect 171140 325660 171192 325712
rect 204996 325660 205048 325712
rect 269120 325660 269172 325712
rect 188528 325592 188580 325644
rect 214564 325592 214616 325644
rect 214564 325116 214616 325168
rect 215116 325116 215168 325168
rect 170496 324980 170548 325032
rect 186320 324980 186372 325032
rect 162124 324912 162176 324964
rect 234436 324912 234488 324964
rect 251916 324912 251968 324964
rect 219716 324300 219768 324352
rect 220176 324300 220228 324352
rect 276664 324300 276716 324352
rect 158812 324164 158864 324216
rect 160744 324164 160796 324216
rect 158720 323008 158772 323060
rect 214656 323008 214708 323060
rect 203616 322940 203668 322992
rect 280804 322940 280856 322992
rect 64788 322872 64840 322924
rect 65800 322872 65852 322924
rect 158720 322804 158772 322856
rect 161572 322804 161624 322856
rect 65800 322396 65852 322448
rect 66536 322396 66588 322448
rect 159456 322260 159508 322312
rect 220176 322260 220228 322312
rect 238024 322260 238076 322312
rect 259644 322260 259696 322312
rect 162952 322192 163004 322244
rect 246304 322192 246356 322244
rect 273996 322192 274048 322244
rect 317604 322192 317656 322244
rect 326988 322192 327040 322244
rect 340236 322192 340288 322244
rect 254676 321580 254728 321632
rect 325700 321580 325752 321632
rect 326988 321580 327040 321632
rect 4804 321512 4856 321564
rect 66812 321512 66864 321564
rect 174912 320900 174964 320952
rect 240876 320900 240928 320952
rect 158168 320832 158220 320884
rect 228548 320832 228600 320884
rect 166908 320560 166960 320612
rect 170496 320560 170548 320612
rect 158720 320152 158772 320204
rect 163688 320152 163740 320204
rect 240876 320152 240928 320204
rect 356704 320152 356756 320204
rect 158812 320084 158864 320136
rect 166908 320084 166960 320136
rect 167644 319472 167696 319524
rect 200488 319472 200540 319524
rect 4068 319404 4120 319456
rect 11704 319404 11756 319456
rect 53748 319404 53800 319456
rect 66444 319404 66496 319456
rect 171140 319404 171192 319456
rect 210424 319404 210476 319456
rect 213368 319404 213420 319456
rect 283564 319404 283616 319456
rect 327816 319404 327868 319456
rect 371424 319404 371476 319456
rect 202788 318792 202840 318844
rect 308404 318792 308456 318844
rect 64604 318588 64656 318640
rect 66444 318588 66496 318640
rect 160836 318112 160888 318164
rect 166448 318112 166500 318164
rect 167920 318112 167972 318164
rect 193956 318112 194008 318164
rect 194048 318112 194100 318164
rect 216036 318112 216088 318164
rect 54944 318044 54996 318096
rect 64144 318044 64196 318096
rect 156788 318044 156840 318096
rect 167828 318044 167880 318096
rect 170588 318044 170640 318096
rect 199568 318044 199620 318096
rect 213276 318044 213328 318096
rect 251272 318044 251324 318096
rect 340880 317500 340932 317552
rect 342168 317500 342220 317552
rect 396724 317500 396776 317552
rect 228456 317432 228508 317484
rect 347044 317432 347096 317484
rect 186320 317364 186372 317416
rect 204996 317364 205048 317416
rect 262404 317364 262456 317416
rect 262864 317364 262916 317416
rect 4804 316684 4856 316736
rect 64512 316684 64564 316736
rect 66904 316684 66956 316736
rect 160008 316684 160060 316736
rect 161296 316684 161348 316736
rect 166356 316684 166408 316736
rect 165068 316480 165120 316532
rect 165528 316480 165580 316532
rect 208124 316072 208176 316124
rect 209780 316072 209832 316124
rect 210976 316072 211028 316124
rect 240140 316072 240192 316124
rect 262404 316072 262456 316124
rect 165068 316004 165120 316056
rect 246396 316004 246448 316056
rect 158812 315936 158864 315988
rect 168288 315936 168340 315988
rect 168288 315324 168340 315376
rect 182824 315324 182876 315376
rect 204904 315324 204956 315376
rect 232688 315324 232740 315376
rect 177488 315256 177540 315308
rect 223028 315256 223080 315308
rect 232596 315256 232648 315308
rect 244372 315256 244424 315308
rect 52092 314644 52144 314696
rect 56508 314644 56560 314696
rect 66812 314644 66864 314696
rect 195980 314644 196032 314696
rect 198740 314644 198792 314696
rect 222476 314644 222528 314696
rect 223028 314644 223080 314696
rect 255504 314644 255556 314696
rect 60372 314576 60424 314628
rect 66904 314576 66956 314628
rect 223488 313896 223540 313948
rect 240140 313896 240192 313948
rect 302332 313896 302384 313948
rect 358820 313896 358872 313948
rect 238576 313352 238628 313404
rect 271880 313352 271932 313404
rect 272524 313352 272576 313404
rect 158812 313284 158864 313336
rect 192484 313284 192536 313336
rect 241980 313284 242032 313336
rect 242256 313284 242308 313336
rect 302332 313284 302384 313336
rect 161572 312536 161624 312588
rect 235356 312536 235408 312588
rect 293224 312536 293276 312588
rect 338764 312536 338816 312588
rect 202144 311856 202196 311908
rect 209228 311856 209280 311908
rect 227812 311856 227864 311908
rect 228548 311856 228600 311908
rect 282920 311856 282972 311908
rect 238116 311788 238168 311840
rect 239404 311788 239456 311840
rect 187608 311176 187660 311228
rect 194600 311176 194652 311228
rect 238024 311176 238076 311228
rect 239404 311176 239456 311228
rect 239588 311176 239640 311228
rect 254676 311176 254728 311228
rect 11704 311108 11756 311160
rect 67088 311108 67140 311160
rect 67456 311108 67508 311160
rect 197176 311108 197228 311160
rect 287704 311108 287756 311160
rect 158904 310496 158956 310548
rect 194600 310496 194652 310548
rect 158812 310428 158864 310480
rect 164240 310428 164292 310480
rect 165528 310428 165580 310480
rect 238668 310428 238720 310480
rect 240232 310428 240284 310480
rect 165528 309816 165580 309868
rect 177488 309816 177540 309868
rect 35164 309748 35216 309800
rect 62764 309748 62816 309800
rect 66812 309748 66864 309800
rect 171968 309748 172020 309800
rect 223488 309748 223540 309800
rect 262128 309748 262180 309800
rect 313924 309748 313976 309800
rect 208492 309136 208544 309188
rect 209228 309136 209280 309188
rect 279424 309136 279476 309188
rect 158812 308932 158864 308984
rect 162860 308932 162912 308984
rect 166540 308932 166592 308984
rect 282184 307844 282236 307896
rect 199568 307776 199620 307828
rect 200028 307776 200080 307828
rect 239036 307776 239088 307828
rect 381544 307776 381596 307828
rect 61752 307708 61804 307760
rect 66904 307708 66956 307760
rect 197084 307096 197136 307148
rect 204352 307096 204404 307148
rect 190276 307028 190328 307080
rect 204260 307028 204312 307080
rect 207756 306416 207808 306468
rect 244004 306416 244056 306468
rect 158812 306348 158864 306400
rect 170404 306348 170456 306400
rect 209412 306348 209464 306400
rect 267096 306348 267148 306400
rect 3332 306280 3384 306332
rect 33784 306280 33836 306332
rect 310428 305600 310480 305652
rect 363236 305600 363288 305652
rect 199476 305056 199528 305108
rect 200120 305056 200172 305108
rect 201408 305056 201460 305108
rect 212724 305056 212776 305108
rect 267832 305056 267884 305108
rect 56416 304988 56468 305040
rect 66812 304988 66864 305040
rect 158812 304988 158864 305040
rect 236000 304988 236052 305040
rect 236092 304988 236144 305040
rect 236736 304988 236788 305040
rect 294604 304920 294656 304972
rect 367100 304920 367152 304972
rect 175188 304308 175240 304360
rect 188436 304308 188488 304360
rect 192760 304308 192812 304360
rect 220176 304308 220228 304360
rect 234528 304308 234580 304360
rect 280988 304308 281040 304360
rect 184296 304240 184348 304292
rect 208952 304240 209004 304292
rect 209044 304240 209096 304292
rect 215208 304240 215260 304292
rect 358084 304240 358136 304292
rect 158812 303968 158864 304020
rect 160836 303968 160888 304020
rect 158812 303628 158864 303680
rect 175188 303628 175240 303680
rect 231676 303628 231728 303680
rect 234528 303628 234580 303680
rect 64696 303560 64748 303612
rect 66904 303560 66956 303612
rect 193404 302880 193456 302932
rect 212724 302880 212776 302932
rect 322204 302880 322256 302932
rect 355324 302880 355376 302932
rect 202236 302268 202288 302320
rect 274088 302268 274140 302320
rect 215300 302200 215352 302252
rect 215852 302200 215904 302252
rect 288440 302200 288492 302252
rect 58992 302132 59044 302184
rect 66904 302132 66956 302184
rect 164976 301520 165028 301572
rect 251364 301520 251416 301572
rect 262956 301520 263008 301572
rect 293960 301520 294012 301572
rect 327724 301520 327776 301572
rect 330484 301520 330536 301572
rect 160008 301452 160060 301504
rect 165620 301452 165672 301504
rect 166080 301452 166132 301504
rect 193864 301452 193916 301504
rect 221556 301452 221608 301504
rect 238024 301452 238076 301504
rect 353944 301452 353996 301504
rect 64696 300840 64748 300892
rect 66812 300840 66864 300892
rect 158996 300296 159048 300348
rect 160100 300296 160152 300348
rect 160928 300296 160980 300348
rect 163688 300160 163740 300212
rect 245752 300160 245804 300212
rect 158812 300092 158864 300144
rect 244464 300092 244516 300144
rect 249156 299480 249208 299532
rect 443000 299480 443052 299532
rect 56324 299412 56376 299464
rect 66628 299412 66680 299464
rect 158812 299412 158864 299464
rect 173256 299412 173308 299464
rect 180248 298800 180300 298852
rect 230388 298800 230440 298852
rect 243452 298800 243504 298852
rect 245660 298800 245712 298852
rect 201316 298732 201368 298784
rect 254676 298732 254728 298784
rect 298100 298732 298152 298784
rect 369860 298732 369912 298784
rect 194324 298120 194376 298172
rect 200304 298120 200356 298172
rect 201316 298120 201368 298172
rect 57888 298052 57940 298104
rect 58992 298052 59044 298104
rect 193956 297508 194008 297560
rect 204260 297508 204312 297560
rect 167828 297440 167880 297492
rect 180248 297440 180300 297492
rect 183376 297440 183428 297492
rect 203524 297440 203576 297492
rect 58992 297372 59044 297424
rect 66812 297372 66864 297424
rect 165160 297372 165212 297424
rect 193404 297372 193456 297424
rect 246396 297372 246448 297424
rect 256700 297372 256752 297424
rect 158812 296692 158864 296744
rect 168288 296692 168340 296744
rect 231124 296692 231176 296744
rect 247132 296692 247184 296744
rect 166816 296012 166868 296064
rect 187056 296012 187108 296064
rect 158812 295944 158864 295996
rect 209044 295944 209096 295996
rect 214564 295400 214616 295452
rect 224316 295400 224368 295452
rect 273168 295400 273220 295452
rect 278228 295400 278280 295452
rect 30288 295332 30340 295384
rect 67180 295332 67232 295384
rect 189908 295332 189960 295384
rect 190368 295332 190420 295384
rect 439412 295332 439464 295384
rect 158812 295264 158864 295316
rect 177396 295264 177448 295316
rect 235264 295264 235316 295316
rect 392676 295264 392728 295316
rect 392676 294584 392728 294636
rect 414664 294584 414716 294636
rect 177304 294040 177356 294092
rect 202236 294040 202288 294092
rect 195336 293972 195388 294024
rect 259736 293972 259788 294024
rect 26148 293904 26200 293956
rect 66812 293904 66864 293956
rect 158812 292612 158864 292664
rect 193864 292612 193916 292664
rect 3608 292544 3660 292596
rect 18604 292544 18656 292596
rect 158904 292544 158956 292596
rect 220176 292544 220228 292596
rect 221556 292544 221608 292596
rect 222108 292544 222160 292596
rect 253204 292612 253256 292664
rect 234436 292544 234488 292596
rect 295432 292544 295484 292596
rect 53564 292476 53616 292528
rect 66812 292476 66864 292528
rect 247132 291796 247184 291848
rect 253940 291796 253992 291848
rect 256056 291796 256108 291848
rect 263784 291796 263836 291848
rect 187516 291320 187568 291372
rect 192576 291320 192628 291372
rect 195152 291252 195204 291304
rect 247316 291252 247368 291304
rect 158812 291184 158864 291236
rect 247132 291184 247184 291236
rect 60464 291116 60516 291168
rect 66352 291116 66404 291168
rect 59176 291048 59228 291100
rect 67088 291048 67140 291100
rect 199568 290776 199620 290828
rect 201500 290776 201552 290828
rect 162216 290436 162268 290488
rect 195152 290436 195204 290488
rect 295892 290436 295944 290488
rect 371240 290436 371292 290488
rect 210424 289892 210476 289944
rect 248420 289892 248472 289944
rect 158812 289824 158864 289876
rect 216680 289824 216732 289876
rect 229744 289824 229796 289876
rect 255320 289824 255372 289876
rect 258908 289824 258960 289876
rect 322296 289824 322348 289876
rect 186964 289756 187016 289808
rect 188436 289756 188488 289808
rect 64144 289212 64196 289264
rect 66812 289212 66864 289264
rect 158812 289212 158864 289264
rect 162768 289212 162820 289264
rect 169024 289076 169076 289128
rect 181444 289076 181496 289128
rect 216680 289076 216732 289128
rect 224868 289076 224920 289128
rect 240508 289076 240560 289128
rect 258908 289076 258960 289128
rect 200028 288464 200080 288516
rect 201684 288464 201736 288516
rect 176108 288396 176160 288448
rect 216680 288396 216732 288448
rect 224868 288396 224920 288448
rect 247500 288396 247552 288448
rect 332600 288396 332652 288448
rect 447140 288396 447192 288448
rect 158904 288328 158956 288380
rect 231124 288328 231176 288380
rect 259552 288192 259604 288244
rect 260104 288192 260156 288244
rect 66168 287784 66220 287836
rect 67364 287784 67416 287836
rect 164976 287648 165028 287700
rect 195152 287648 195204 287700
rect 235356 287648 235408 287700
rect 245844 287648 245896 287700
rect 303620 287648 303672 287700
rect 364340 287648 364392 287700
rect 376116 287648 376168 287700
rect 392584 287648 392636 287700
rect 233148 287104 233200 287156
rect 260104 287104 260156 287156
rect 158812 287036 158864 287088
rect 162124 287036 162176 287088
rect 198740 287036 198792 287088
rect 223580 287036 223632 287088
rect 245844 287036 245896 287088
rect 303620 287036 303672 287088
rect 57612 286968 57664 287020
rect 66812 286968 66864 287020
rect 232688 286968 232740 287020
rect 234252 286968 234304 287020
rect 218612 286628 218664 286680
rect 220084 286628 220136 286680
rect 224224 286356 224276 286408
rect 225052 286356 225104 286408
rect 158812 286288 158864 286340
rect 165068 286288 165120 286340
rect 172060 286288 172112 286340
rect 195336 286288 195388 286340
rect 356704 286084 356756 286136
rect 363604 286084 363656 286136
rect 166448 285948 166500 286000
rect 171876 285948 171928 286000
rect 201408 285812 201460 285864
rect 205548 285812 205600 285864
rect 204996 285744 205048 285796
rect 207020 285744 207072 285796
rect 212908 285744 212960 285796
rect 218060 285744 218112 285796
rect 227628 285744 227680 285796
rect 228916 285744 228968 285796
rect 237380 285744 237432 285796
rect 238484 285744 238536 285796
rect 245016 285744 245068 285796
rect 63408 285676 63460 285728
rect 66260 285676 66312 285728
rect 166356 285676 166408 285728
rect 171968 285676 172020 285728
rect 191104 285676 191156 285728
rect 210884 285676 210936 285728
rect 211804 285676 211856 285728
rect 213828 285676 213880 285728
rect 215208 285676 215260 285728
rect 219164 285676 219216 285728
rect 224316 285676 224368 285728
rect 226524 285676 226576 285728
rect 228364 285676 228416 285728
rect 229284 285676 229336 285728
rect 234436 285676 234488 285728
rect 235172 285676 235224 285728
rect 237564 285676 237616 285728
rect 238576 285676 238628 285728
rect 242348 285676 242400 285728
rect 267004 285676 267056 285728
rect 200120 285268 200172 285320
rect 200948 285268 201000 285320
rect 220820 285268 220872 285320
rect 221280 285268 221332 285320
rect 158168 284928 158220 284980
rect 177580 284928 177632 284980
rect 237472 284928 237524 284980
rect 243912 284928 243964 284980
rect 254676 284928 254728 284980
rect 261576 284928 261628 284980
rect 185676 284384 185728 284436
rect 216772 284384 216824 284436
rect 247040 284384 247092 284436
rect 247684 284384 247736 284436
rect 254584 284384 254636 284436
rect 57888 284316 57940 284368
rect 66812 284316 66864 284368
rect 173256 284316 173308 284368
rect 198740 284316 198792 284368
rect 204628 284316 204680 284368
rect 206652 284316 206704 284368
rect 428464 284316 428516 284368
rect 203340 284248 203392 284300
rect 332600 284248 332652 284300
rect 333888 284248 333940 284300
rect 358176 284248 358228 284300
rect 199476 283908 199528 283960
rect 201408 283908 201460 283960
rect 170588 283568 170640 283620
rect 198832 283568 198884 283620
rect 246304 283568 246356 283620
rect 246856 283568 246908 283620
rect 251180 283568 251232 283620
rect 280988 282956 281040 283008
rect 281724 282956 281776 283008
rect 59176 282888 59228 282940
rect 66812 282888 66864 282940
rect 263600 282888 263652 282940
rect 264888 282888 264940 282940
rect 380164 282888 380216 282940
rect 183284 282820 183336 282872
rect 195152 282820 195204 282872
rect 160100 282140 160152 282192
rect 176660 282140 176712 282192
rect 247500 282140 247552 282192
rect 263600 282140 263652 282192
rect 245936 281664 245988 281716
rect 251088 281664 251140 281716
rect 253204 281664 253256 281716
rect 255504 281664 255556 281716
rect 176660 281528 176712 281580
rect 177948 281528 178000 281580
rect 197360 281528 197412 281580
rect 250628 281460 250680 281512
rect 255504 281460 255556 281512
rect 166540 281392 166592 281444
rect 197360 281392 197412 281444
rect 160836 280780 160888 280832
rect 197176 280780 197228 280832
rect 197452 280780 197504 280832
rect 286416 280780 286468 280832
rect 318064 280780 318116 280832
rect 279056 280576 279108 280628
rect 283564 280576 283616 280628
rect 158812 280236 158864 280288
rect 160928 280236 160980 280288
rect 17868 280168 17920 280220
rect 67548 280168 67600 280220
rect 246120 280168 246172 280220
rect 318800 280168 318852 280220
rect 165528 279760 165580 279812
rect 168564 279760 168616 279812
rect 170404 279488 170456 279540
rect 179420 279488 179472 279540
rect 245936 279488 245988 279540
rect 309784 279488 309836 279540
rect 159364 279420 159416 279472
rect 191840 279420 191892 279472
rect 286324 279420 286376 279472
rect 294604 279420 294656 279472
rect 304264 279420 304316 279472
rect 449900 279420 449952 279472
rect 245936 278944 245988 278996
rect 249156 278944 249208 278996
rect 60280 278740 60332 278792
rect 66628 278740 66680 278792
rect 179420 278740 179472 278792
rect 180708 278740 180760 278792
rect 197360 278740 197412 278792
rect 52184 278672 52236 278724
rect 66812 278672 66864 278724
rect 192668 278672 192720 278724
rect 197176 278672 197228 278724
rect 197452 278672 197504 278724
rect 195888 278604 195940 278656
rect 197360 278604 197412 278656
rect 245936 277992 245988 278044
rect 249892 277992 249944 278044
rect 378232 277992 378284 278044
rect 382924 277992 382976 278044
rect 158628 277380 158680 277432
rect 167644 277380 167696 277432
rect 244372 277380 244424 277432
rect 285036 277380 285088 277432
rect 60556 277312 60608 277364
rect 66260 277312 66312 277364
rect 158812 277312 158864 277364
rect 165160 277312 165212 277364
rect 160928 276632 160980 276684
rect 183284 276632 183336 276684
rect 245752 276632 245804 276684
rect 293960 276632 294012 276684
rect 360200 276632 360252 276684
rect 183284 276088 183336 276140
rect 61844 276020 61896 276072
rect 66812 276020 66864 276072
rect 186228 276020 186280 276072
rect 187240 276020 187292 276072
rect 197452 276020 197504 276072
rect 166908 275952 166960 276004
rect 172520 275952 172572 276004
rect 197268 275952 197320 276004
rect 197544 275952 197596 276004
rect 245936 275952 245988 276004
rect 257344 275952 257396 276004
rect 268384 275952 268436 276004
rect 338856 275952 338908 276004
rect 158812 275884 158864 275936
rect 162216 275884 162268 275936
rect 159824 275272 159876 275324
rect 177396 275272 177448 275324
rect 245936 275272 245988 275324
rect 252836 275272 252888 275324
rect 252836 274660 252888 274712
rect 307116 274660 307168 274712
rect 61936 274592 61988 274644
rect 65892 274592 65944 274644
rect 158812 274592 158864 274644
rect 176108 274592 176160 274644
rect 183468 274524 183520 274576
rect 185032 274524 185084 274576
rect 267188 273980 267240 274032
rect 354128 273980 354180 274032
rect 181720 273912 181772 273964
rect 199476 273912 199528 273964
rect 322204 273912 322256 273964
rect 436744 273912 436796 273964
rect 191840 273436 191892 273488
rect 193036 273436 193088 273488
rect 197452 273436 197504 273488
rect 158812 273232 158864 273284
rect 173348 273232 173400 273284
rect 175096 273164 175148 273216
rect 197452 273164 197504 273216
rect 245844 273164 245896 273216
rect 248604 273164 248656 273216
rect 251272 273164 251324 273216
rect 180248 272484 180300 272536
rect 191380 272484 191432 272536
rect 245936 272484 245988 272536
rect 251272 272484 251324 272536
rect 252468 272484 252520 272536
rect 280896 272484 280948 272536
rect 294604 272484 294656 272536
rect 307668 272484 307720 272536
rect 385040 272484 385092 272536
rect 176108 272280 176160 272332
rect 178684 272280 178736 272332
rect 63132 271872 63184 271924
rect 66260 271872 66312 271924
rect 252468 271872 252520 271924
rect 306380 271872 306432 271924
rect 307668 271872 307720 271924
rect 245936 271192 245988 271244
rect 248604 271192 248656 271244
rect 61936 271124 61988 271176
rect 66904 271124 66956 271176
rect 184756 271124 184808 271176
rect 199568 271124 199620 271176
rect 245844 271124 245896 271176
rect 305184 271124 305236 271176
rect 380900 271124 380952 271176
rect 158812 270784 158864 270836
rect 162216 270784 162268 270836
rect 54944 270512 54996 270564
rect 66904 270512 66956 270564
rect 164148 270512 164200 270564
rect 197452 270512 197504 270564
rect 184388 270444 184440 270496
rect 185768 270444 185820 270496
rect 245936 270172 245988 270224
rect 248512 270172 248564 270224
rect 4068 269764 4120 269816
rect 32404 269764 32456 269816
rect 260104 269764 260156 269816
rect 367744 269764 367796 269816
rect 163688 269084 163740 269136
rect 197452 269084 197504 269136
rect 12440 269016 12492 269068
rect 14464 269016 14516 269068
rect 63316 269016 63368 269068
rect 64788 269016 64840 269068
rect 158812 269016 158864 269068
rect 170588 269016 170640 269068
rect 172428 269016 172480 269068
rect 178684 269016 178736 269068
rect 181536 269016 181588 269068
rect 184296 269016 184348 269068
rect 194416 269016 194468 269068
rect 194692 269016 194744 269068
rect 291844 268948 291896 269000
rect 293224 268948 293276 269000
rect 161296 268336 161348 268388
rect 187332 268336 187384 268388
rect 311992 268336 312044 268388
rect 367192 268336 367244 268388
rect 194692 267996 194744 268048
rect 198280 267996 198332 268048
rect 64788 267860 64840 267912
rect 66812 267860 66864 267912
rect 187332 267724 187384 267776
rect 197544 267724 197596 267776
rect 244464 267724 244516 267776
rect 311992 267724 312044 267776
rect 187608 267656 187660 267708
rect 197452 267656 197504 267708
rect 245752 267656 245804 267708
rect 259644 267656 259696 267708
rect 194324 267112 194376 267164
rect 197544 267112 197596 267164
rect 3148 266976 3200 267028
rect 12440 266976 12492 267028
rect 259644 266976 259696 267028
rect 336096 266976 336148 267028
rect 191288 266908 191340 266960
rect 193220 266908 193272 266960
rect 12440 266364 12492 266416
rect 13084 266364 13136 266416
rect 256792 266364 256844 266416
rect 158812 266296 158864 266348
rect 172060 266296 172112 266348
rect 246028 266296 246080 266348
rect 358176 266296 358228 266348
rect 583300 266296 583352 266348
rect 180616 265684 180668 265736
rect 181444 265684 181496 265736
rect 189816 265684 189868 265736
rect 196624 265684 196676 265736
rect 167736 265616 167788 265668
rect 194324 265616 194376 265668
rect 245844 265616 245896 265668
rect 252560 265616 252612 265668
rect 276756 265616 276808 265668
rect 292580 265616 292632 265668
rect 54852 264936 54904 264988
rect 66812 264936 66864 264988
rect 158812 264868 158864 264920
rect 188528 264868 188580 264920
rect 190368 264868 190420 264920
rect 197452 264868 197504 264920
rect 257436 264256 257488 264308
rect 291200 264256 291252 264308
rect 55128 264188 55180 264240
rect 62120 264188 62172 264240
rect 170588 264188 170640 264240
rect 177304 264188 177356 264240
rect 259368 264188 259420 264240
rect 377496 264188 377548 264240
rect 62120 263576 62172 263628
rect 63224 263576 63276 263628
rect 66904 263576 66956 263628
rect 182088 263576 182140 263628
rect 197452 263576 197504 263628
rect 158812 263508 158864 263560
rect 166264 263508 166316 263560
rect 245016 262964 245068 263016
rect 246396 262964 246448 263016
rect 43996 262828 44048 262880
rect 52460 262828 52512 262880
rect 172428 262828 172480 262880
rect 194692 262828 194744 262880
rect 52460 262216 52512 262268
rect 53564 262216 53616 262268
rect 66812 262216 66864 262268
rect 159456 262216 159508 262268
rect 181444 262216 181496 262268
rect 182088 262216 182140 262268
rect 193128 262216 193180 262268
rect 194784 262216 194836 262268
rect 156788 262148 156840 262200
rect 159548 262148 159600 262200
rect 158628 262080 158680 262132
rect 178776 262148 178828 262200
rect 245844 262216 245896 262268
rect 248512 262216 248564 262268
rect 258908 262216 258960 262268
rect 356796 262216 356848 262268
rect 198096 262148 198148 262200
rect 254584 261536 254636 261588
rect 300124 261536 300176 261588
rect 32404 261468 32456 261520
rect 51080 261468 51132 261520
rect 188436 261468 188488 261520
rect 196808 261468 196860 261520
rect 57612 260924 57664 260976
rect 66812 260924 66864 260976
rect 51080 260856 51132 260908
rect 52184 260856 52236 260908
rect 66260 260856 66312 260908
rect 167092 260856 167144 260908
rect 197452 260856 197504 260908
rect 246028 260788 246080 260840
rect 255504 260788 255556 260840
rect 317328 260788 317380 260840
rect 318064 260788 318116 260840
rect 157984 260108 158036 260160
rect 191288 260108 191340 260160
rect 303712 260108 303764 260160
rect 374000 260108 374052 260160
rect 158904 259428 158956 259480
rect 166264 259428 166316 259480
rect 188436 259428 188488 259480
rect 197452 259428 197504 259480
rect 245660 259428 245712 259480
rect 303712 259428 303764 259480
rect 182088 259360 182140 259412
rect 185676 259360 185728 259412
rect 245844 259360 245896 259412
rect 260932 259360 260984 259412
rect 262128 259360 262180 259412
rect 262128 258748 262180 258800
rect 292764 258748 292816 258800
rect 361672 258748 361724 258800
rect 165068 258680 165120 258732
rect 174728 258680 174780 258732
rect 288532 258680 288584 258732
rect 369952 258680 370004 258732
rect 175096 258544 175148 258596
rect 176108 258544 176160 258596
rect 191840 258476 191892 258528
rect 197452 258476 197504 258528
rect 34428 258000 34480 258052
rect 61384 258000 61436 258052
rect 66260 258068 66312 258120
rect 158812 258068 158864 258120
rect 182088 258136 182140 258188
rect 189724 258136 189776 258188
rect 191840 258136 191892 258188
rect 185584 258068 185636 258120
rect 191104 258068 191156 258120
rect 245660 258068 245712 258120
rect 288532 258068 288584 258120
rect 245844 258000 245896 258052
rect 256700 258000 256752 258052
rect 273904 257388 273956 257440
rect 348424 257388 348476 257440
rect 162216 257320 162268 257372
rect 184204 257320 184256 257372
rect 250536 257320 250588 257372
rect 441620 257320 441672 257372
rect 159272 257048 159324 257100
rect 160836 257048 160888 257100
rect 189724 256776 189776 256828
rect 197452 256776 197504 256828
rect 64512 256708 64564 256760
rect 66904 256708 66956 256760
rect 184204 256708 184256 256760
rect 184664 256708 184716 256760
rect 197544 256708 197596 256760
rect 256700 256708 256752 256760
rect 260104 256708 260156 256760
rect 178040 256640 178092 256692
rect 179328 256640 179380 256692
rect 197452 256640 197504 256692
rect 245844 256640 245896 256692
rect 254124 256640 254176 256692
rect 245844 256028 245896 256080
rect 258172 256028 258224 256080
rect 162216 255960 162268 256012
rect 178040 255960 178092 256012
rect 254124 255960 254176 256012
rect 309232 255960 309284 256012
rect 363144 255960 363196 256012
rect 60464 255280 60516 255332
rect 66812 255280 66864 255332
rect 158812 255280 158864 255332
rect 173808 255280 173860 255332
rect 257528 255280 257580 255332
rect 300860 255280 300912 255332
rect 194416 255212 194468 255264
rect 197452 255212 197504 255264
rect 246028 255212 246080 255264
rect 251364 255212 251416 255264
rect 252468 255212 252520 255264
rect 245844 255144 245896 255196
rect 247316 255144 247368 255196
rect 252468 254600 252520 254652
rect 322204 254600 322256 254652
rect 158812 254532 158864 254584
rect 189724 254532 189776 254584
rect 258172 254532 258224 254584
rect 384304 254532 384356 254584
rect 3148 253920 3200 253972
rect 10968 253920 11020 253972
rect 11704 253920 11756 253972
rect 63316 253920 63368 253972
rect 66812 253920 66864 253972
rect 158904 253920 158956 253972
rect 162768 253920 162820 253972
rect 247040 253920 247092 253972
rect 247316 253920 247368 253972
rect 246028 253852 246080 253904
rect 267832 253852 267884 253904
rect 269028 253852 269080 253904
rect 314660 253240 314712 253292
rect 359004 253240 359056 253292
rect 39948 253172 40000 253224
rect 60096 253172 60148 253224
rect 185768 253172 185820 253224
rect 197912 253172 197964 253224
rect 198372 253172 198424 253224
rect 269028 253172 269080 253224
rect 300952 253172 301004 253224
rect 372620 253172 372672 253224
rect 158812 252628 158864 252680
rect 176108 252628 176160 252680
rect 60096 252560 60148 252612
rect 60372 252560 60424 252612
rect 66812 252560 66864 252612
rect 159640 252560 159692 252612
rect 195888 252560 195940 252612
rect 197452 252560 197504 252612
rect 245660 252560 245712 252612
rect 314660 252560 314712 252612
rect 246028 252492 246080 252544
rect 263692 252492 263744 252544
rect 245844 252220 245896 252272
rect 249800 252220 249852 252272
rect 251088 252220 251140 252272
rect 159364 251880 159416 251932
rect 173440 251948 173492 252000
rect 173808 251880 173860 251932
rect 194324 251880 194376 251932
rect 291108 251880 291160 251932
rect 302240 251880 302292 251932
rect 309876 251880 309928 251932
rect 345664 251880 345716 251932
rect 162768 251812 162820 251864
rect 183284 251812 183336 251864
rect 183560 251812 183612 251864
rect 263692 251812 263744 251864
rect 460940 251812 460992 251864
rect 65892 251744 65944 251796
rect 66996 251744 67048 251796
rect 194324 251608 194376 251660
rect 197084 251608 197136 251660
rect 191380 251200 191432 251252
rect 193128 251200 193180 251252
rect 158812 251132 158864 251184
rect 166356 251132 166408 251184
rect 307760 250520 307812 250572
rect 356060 250520 356112 250572
rect 160928 250452 160980 250504
rect 167736 250452 167788 250504
rect 173348 250452 173400 250504
rect 191748 250452 191800 250504
rect 317328 250452 317380 250504
rect 368480 250452 368532 250504
rect 252468 249840 252520 249892
rect 285128 249840 285180 249892
rect 191104 249772 191156 249824
rect 197452 249772 197504 249824
rect 247316 249772 247368 249824
rect 316040 249772 316092 249824
rect 317328 249772 317380 249824
rect 246028 249704 246080 249756
rect 251824 249704 251876 249756
rect 252468 249704 252520 249756
rect 191748 249500 191800 249552
rect 197452 249500 197504 249552
rect 181536 249364 181588 249416
rect 189816 249364 189868 249416
rect 284944 249092 284996 249144
rect 307852 249092 307904 249144
rect 265716 249024 265768 249076
rect 429844 249024 429896 249076
rect 193128 248684 193180 248736
rect 197452 248684 197504 248736
rect 175924 248480 175976 248532
rect 181720 248480 181772 248532
rect 67548 248412 67600 248464
rect 67916 248412 67968 248464
rect 158812 248412 158864 248464
rect 187148 248412 187200 248464
rect 67548 248276 67600 248328
rect 67916 248276 67968 248328
rect 159548 247052 159600 247104
rect 196716 247120 196768 247172
rect 197268 247120 197320 247172
rect 195336 247052 195388 247104
rect 197728 247052 197780 247104
rect 245016 247052 245068 247104
rect 245660 247052 245712 247104
rect 245844 247052 245896 247104
rect 267832 247052 267884 247104
rect 60648 246984 60700 247036
rect 66812 246984 66864 247036
rect 158812 246372 158864 246424
rect 176200 246372 176252 246424
rect 184204 246372 184256 246424
rect 245660 246372 245712 246424
rect 253112 246372 253164 246424
rect 257344 246372 257396 246424
rect 269120 246372 269172 246424
rect 274088 246372 274140 246424
rect 291200 246372 291252 246424
rect 162124 246304 162176 246356
rect 199476 246304 199528 246356
rect 246304 246304 246356 246356
rect 283564 246304 283616 246356
rect 64604 245624 64656 245676
rect 66812 245624 66864 245676
rect 194232 245624 194284 245676
rect 194600 245624 194652 245676
rect 48136 245556 48188 245608
rect 66904 245556 66956 245608
rect 180524 245556 180576 245608
rect 181628 245556 181680 245608
rect 260748 244944 260800 244996
rect 313280 244944 313332 244996
rect 352656 244944 352708 244996
rect 158812 244876 158864 244928
rect 171784 244876 171836 244928
rect 180156 244876 180208 244928
rect 189080 244876 189132 244928
rect 190368 244876 190420 244928
rect 197360 244876 197412 244928
rect 270408 244876 270460 244928
rect 583024 244876 583076 244928
rect 67088 244400 67140 244452
rect 67364 244400 67416 244452
rect 158812 244264 158864 244316
rect 177304 244264 177356 244316
rect 269948 244264 270000 244316
rect 270408 244264 270460 244316
rect 59268 244196 59320 244248
rect 67456 244196 67508 244248
rect 246396 244196 246448 244248
rect 249984 244196 250036 244248
rect 262128 243380 262180 243432
rect 262404 243380 262456 243432
rect 158812 242972 158864 243024
rect 181720 242972 181772 243024
rect 190184 242972 190236 243024
rect 197360 242972 197412 243024
rect 245752 242972 245804 243024
rect 262128 242972 262180 243024
rect 156972 242904 157024 242956
rect 191196 242904 191248 242956
rect 262772 242904 262824 242956
rect 409880 242904 409932 242956
rect 161020 242224 161072 242276
rect 164148 242224 164200 242276
rect 177488 242224 177540 242276
rect 156880 242156 156932 242208
rect 187516 242156 187568 242208
rect 199568 242156 199620 242208
rect 310612 242156 310664 242208
rect 345756 242156 345808 242208
rect 153108 241476 153160 241528
rect 156696 241476 156748 241528
rect 246120 241476 246172 241528
rect 310612 241476 310664 241528
rect 57796 241408 57848 241460
rect 83326 241408 83378 241460
rect 111110 241408 111162 241460
rect 159640 241408 159692 241460
rect 67088 241340 67140 241392
rect 73804 241340 73856 241392
rect 3332 241068 3384 241120
rect 7564 241068 7616 241120
rect 159456 240796 159508 240848
rect 170588 240796 170640 240848
rect 171876 240796 171928 240848
rect 187056 240796 187108 240848
rect 195796 240796 195848 240848
rect 197912 240796 197964 240848
rect 288348 240796 288400 240848
rect 298744 240796 298796 240848
rect 98368 240728 98420 240780
rect 160928 240728 160980 240780
rect 165160 240728 165212 240780
rect 179420 240728 179472 240780
rect 245660 240728 245712 240780
rect 452660 240728 452712 240780
rect 200120 240184 200172 240236
rect 77300 240116 77352 240168
rect 77852 240116 77904 240168
rect 89720 240116 89772 240168
rect 90364 240116 90416 240168
rect 91100 240116 91152 240168
rect 91836 240116 91888 240168
rect 139400 240116 139452 240168
rect 140044 240116 140096 240168
rect 186320 240116 186372 240168
rect 202880 240116 202932 240168
rect 203432 240116 203484 240168
rect 220728 240116 220780 240168
rect 220912 240116 220964 240168
rect 223304 240116 223356 240168
rect 232136 240116 232188 240168
rect 245660 240184 245712 240236
rect 287244 240116 287296 240168
rect 288348 240116 288400 240168
rect 69480 240048 69532 240100
rect 72516 240048 72568 240100
rect 72608 240048 72660 240100
rect 73068 240048 73120 240100
rect 81900 240048 81952 240100
rect 82728 240048 82780 240100
rect 85580 240048 85632 240100
rect 86868 240048 86920 240100
rect 93032 240048 93084 240100
rect 93768 240048 93820 240100
rect 103796 240048 103848 240100
rect 104808 240048 104860 240100
rect 114652 240048 114704 240100
rect 115204 240048 115256 240100
rect 119344 240048 119396 240100
rect 119988 240048 120040 240100
rect 127164 240048 127216 240100
rect 128268 240048 128320 240100
rect 131856 240048 131908 240100
rect 132316 240048 132368 240100
rect 142896 240048 142948 240100
rect 143448 240048 143500 240100
rect 143632 240048 143684 240100
rect 144276 240048 144328 240100
rect 153292 240048 153344 240100
rect 153844 240048 153896 240100
rect 195244 240048 195296 240100
rect 201132 240048 201184 240100
rect 228732 240048 228784 240100
rect 67364 239980 67416 240032
rect 69664 239980 69716 240032
rect 199844 239980 199896 240032
rect 201040 239980 201092 240032
rect 232596 239980 232648 240032
rect 237472 239980 237524 240032
rect 80704 239912 80756 239964
rect 81256 239912 81308 239964
rect 88800 239912 88852 239964
rect 89536 239912 89588 239964
rect 110696 239912 110748 239964
rect 111708 239912 111760 239964
rect 153752 239912 153804 239964
rect 154488 239912 154540 239964
rect 242624 240048 242676 240100
rect 257528 239912 257580 239964
rect 99656 239776 99708 239828
rect 100576 239776 100628 239828
rect 133328 239708 133380 239760
rect 133788 239708 133840 239760
rect 84108 239436 84160 239488
rect 97356 239436 97408 239488
rect 108948 239436 109000 239488
rect 206008 239436 206060 239488
rect 305092 239436 305144 239488
rect 322940 239436 322992 239488
rect 68928 239368 68980 239420
rect 191840 239368 191892 239420
rect 224408 239368 224460 239420
rect 232044 239368 232096 239420
rect 317512 239368 317564 239420
rect 342260 239368 342312 239420
rect 92572 239232 92624 239284
rect 93124 239232 93176 239284
rect 105544 239232 105596 239284
rect 106188 239232 106240 239284
rect 120816 239232 120868 239284
rect 121368 239232 121420 239284
rect 128912 239232 128964 239284
rect 129556 239232 129608 239284
rect 141424 239232 141476 239284
rect 141976 239232 142028 239284
rect 144184 239232 144236 239284
rect 144828 239232 144880 239284
rect 147128 239232 147180 239284
rect 147588 239232 147640 239284
rect 117320 239164 117372 239216
rect 117964 239164 118016 239216
rect 115112 239096 115164 239148
rect 115848 239096 115900 239148
rect 273168 238824 273220 238876
rect 283196 238824 283248 238876
rect 240324 238756 240376 238808
rect 240876 238756 240928 238808
rect 317512 238756 317564 238808
rect 13084 238688 13136 238740
rect 92572 238688 92624 238740
rect 222292 238688 222344 238740
rect 273168 238688 273220 238740
rect 50896 238620 50948 238672
rect 75920 238620 75972 238672
rect 121644 238620 121696 238672
rect 183376 238620 183428 238672
rect 206008 238620 206060 238672
rect 219900 238620 219952 238672
rect 113180 238552 113232 238604
rect 241796 238620 241848 238672
rect 252652 238620 252704 238672
rect 239220 238144 239272 238196
rect 242716 238144 242768 238196
rect 259368 238076 259420 238128
rect 262956 238076 263008 238128
rect 199384 238008 199436 238060
rect 200212 238008 200264 238060
rect 224776 238008 224828 238060
rect 232964 238008 233016 238060
rect 285128 238008 285180 238060
rect 385684 238008 385736 238060
rect 191840 237668 191892 237720
rect 194416 237668 194468 237720
rect 199384 237668 199436 237720
rect 237472 237532 237524 237584
rect 239404 237532 239456 237584
rect 236828 237464 236880 237516
rect 238024 237464 238076 237516
rect 75920 237396 75972 237448
rect 76564 237396 76616 237448
rect 92572 237396 92624 237448
rect 93124 237396 93176 237448
rect 207112 237396 207164 237448
rect 207940 237396 207992 237448
rect 214196 237396 214248 237448
rect 214656 237396 214708 237448
rect 215668 237396 215720 237448
rect 216496 237396 216548 237448
rect 55036 237328 55088 237380
rect 77392 237328 77444 237380
rect 199568 237328 199620 237380
rect 202972 237328 203024 237380
rect 155960 237260 156012 237312
rect 160744 237260 160796 237312
rect 149060 236784 149112 236836
rect 149244 236784 149296 236836
rect 129004 236716 129056 236768
rect 136824 236716 136876 236768
rect 139492 236716 139544 236768
rect 156972 236716 157024 236768
rect 177304 236716 177356 236768
rect 192944 236716 192996 236768
rect 67732 236648 67784 236700
rect 236644 236648 236696 236700
rect 248604 236648 248656 236700
rect 313372 236648 313424 236700
rect 333980 236648 334032 236700
rect 342904 236648 342956 236700
rect 363696 236648 363748 236700
rect 284944 236036 284996 236088
rect 286416 236036 286468 236088
rect 202972 235968 203024 236020
rect 203524 235968 203576 236020
rect 204076 235968 204128 236020
rect 226984 235968 227036 236020
rect 239404 235968 239456 236020
rect 313372 235968 313424 236020
rect 46848 235900 46900 235952
rect 143632 235900 143684 235952
rect 144184 235900 144236 235952
rect 149060 235900 149112 235952
rect 167644 235900 167696 235952
rect 57704 235832 57756 235884
rect 103520 235832 103572 235884
rect 104716 235832 104768 235884
rect 125600 235832 125652 235884
rect 139492 235832 139544 235884
rect 199476 235832 199528 235884
rect 223764 235832 223816 235884
rect 201132 235560 201184 235612
rect 206376 235560 206428 235612
rect 139584 235220 139636 235272
rect 150440 235220 150492 235272
rect 182088 235220 182140 235272
rect 196624 235220 196676 235272
rect 270408 235220 270460 235272
rect 294696 235220 294748 235272
rect 174636 235084 174688 235136
rect 177304 235084 177356 235136
rect 195980 234880 196032 234932
rect 199384 234880 199436 234932
rect 214748 234676 214800 234728
rect 215116 234676 215168 234728
rect 233332 234676 233384 234728
rect 240784 234676 240836 234728
rect 246028 234676 246080 234728
rect 155224 234608 155276 234660
rect 184756 234608 184808 234660
rect 185032 234608 185084 234660
rect 223764 234608 223816 234660
rect 224224 234608 224276 234660
rect 230204 234608 230256 234660
rect 231952 234608 232004 234660
rect 434812 234608 434864 234660
rect 149244 234540 149296 234592
rect 231860 234540 231912 234592
rect 267648 234540 267700 234592
rect 269764 234540 269816 234592
rect 324320 234540 324372 234592
rect 325608 234540 325660 234592
rect 327724 234540 327776 234592
rect 158076 234472 158128 234524
rect 162308 234472 162360 234524
rect 201316 234472 201368 234524
rect 218152 234472 218204 234524
rect 219900 234472 219952 234524
rect 138020 233928 138072 233980
rect 148324 233928 148376 233980
rect 60280 233860 60332 233912
rect 147680 233860 147732 233912
rect 176108 233860 176160 233912
rect 191196 233860 191248 233912
rect 104900 233180 104952 233232
rect 188436 233180 188488 233232
rect 191288 233180 191340 233232
rect 222844 233180 222896 233232
rect 223396 233180 223448 233232
rect 192484 233112 192536 233164
rect 206836 233112 206888 233164
rect 232964 232568 233016 232620
rect 242164 232568 242216 232620
rect 61936 232500 61988 232552
rect 123484 232500 123536 232552
rect 150440 232500 150492 232552
rect 191656 232500 191708 232552
rect 226156 232500 226208 232552
rect 284392 232500 284444 232552
rect 285036 232500 285088 232552
rect 378784 232500 378836 232552
rect 114284 231752 114336 231804
rect 139492 231820 139544 231872
rect 147680 231752 147732 231804
rect 173256 231752 173308 231804
rect 191656 231752 191708 231804
rect 224408 231752 224460 231804
rect 240048 231752 240100 231804
rect 291292 231752 291344 231804
rect 291844 231752 291896 231804
rect 156604 231684 156656 231736
rect 157984 231684 158036 231736
rect 129556 231208 129608 231260
rect 143356 231208 143408 231260
rect 100576 231140 100628 231192
rect 108304 231140 108356 231192
rect 139124 231140 139176 231192
rect 156880 231140 156932 231192
rect 65892 231072 65944 231124
rect 139216 231072 139268 231124
rect 164148 231072 164200 231124
rect 197268 231072 197320 231124
rect 198556 231072 198608 231124
rect 266360 231072 266412 231124
rect 180064 230460 180116 230512
rect 181628 230460 181680 230512
rect 143356 230392 143408 230444
rect 160100 230392 160152 230444
rect 184664 230392 184716 230444
rect 185676 230392 185728 230444
rect 194232 230392 194284 230444
rect 214748 230392 214800 230444
rect 233056 230392 233108 230444
rect 233424 230392 233476 230444
rect 270408 230392 270460 230444
rect 271144 230392 271196 230444
rect 139492 230324 139544 230376
rect 152740 230324 152792 230376
rect 197268 230324 197320 230376
rect 204996 230324 205048 230376
rect 86960 229780 87012 229832
rect 105544 229780 105596 229832
rect 81256 229712 81308 229764
rect 97264 229712 97316 229764
rect 100760 229712 100812 229764
rect 140780 229712 140832 229764
rect 177396 229712 177448 229764
rect 194232 229712 194284 229764
rect 217324 229712 217376 229764
rect 227260 229712 227312 229764
rect 249800 229780 249852 229832
rect 266360 229780 266412 229832
rect 270408 229780 270460 229832
rect 230388 229712 230440 229764
rect 231124 229712 231176 229764
rect 233424 229712 233476 229764
rect 295340 229712 295392 229764
rect 206836 229100 206888 229152
rect 211804 229100 211856 229152
rect 95332 229032 95384 229084
rect 244280 229032 244332 229084
rect 194232 228964 194284 229016
rect 220084 228964 220136 229016
rect 244280 228760 244332 228812
rect 245016 228760 245068 228812
rect 64512 228352 64564 228404
rect 115020 228352 115072 228404
rect 115848 228352 115900 228404
rect 144736 228352 144788 228404
rect 178040 228352 178092 228404
rect 224408 228352 224460 228404
rect 327816 228352 327868 228404
rect 144092 228284 144144 228336
rect 77208 227672 77260 227724
rect 165160 227672 165212 227724
rect 190460 227672 190512 227724
rect 268384 227672 268436 227724
rect 111708 227604 111760 227656
rect 142160 227604 142212 227656
rect 221648 227604 221700 227656
rect 276020 227604 276072 227656
rect 147680 226992 147732 227044
rect 155224 226992 155276 227044
rect 177488 226992 177540 227044
rect 221556 226992 221608 227044
rect 276020 226992 276072 227044
rect 290096 226992 290148 227044
rect 154580 226312 154632 226364
rect 156788 226312 156840 226364
rect 74540 226244 74592 226296
rect 139124 226244 139176 226296
rect 139216 226244 139268 226296
rect 147680 226244 147732 226296
rect 147772 226244 147824 226296
rect 164884 226244 164936 226296
rect 181720 226244 181772 226296
rect 247132 226244 247184 226296
rect 249800 225632 249852 225684
rect 280160 225632 280212 225684
rect 290464 225632 290516 225684
rect 77300 225564 77352 225616
rect 215944 225564 215996 225616
rect 238024 225564 238076 225616
rect 296812 225564 296864 225616
rect 297364 225564 297416 225616
rect 305644 225564 305696 225616
rect 334624 225564 334676 225616
rect 298468 224952 298520 225004
rect 436100 224952 436152 225004
rect 140780 224272 140832 224324
rect 211068 224272 211120 224324
rect 211436 224272 211488 224324
rect 67824 224204 67876 224256
rect 142804 224204 142856 224256
rect 151728 224204 151780 224256
rect 195244 224204 195296 224256
rect 200764 224204 200816 224256
rect 202236 224204 202288 224256
rect 212448 224204 212500 224256
rect 246120 224204 246172 224256
rect 148324 223524 148376 223576
rect 154580 223524 154632 223576
rect 155224 223524 155276 223576
rect 174544 223524 174596 223576
rect 224316 223524 224368 223576
rect 224868 223524 224920 223576
rect 132316 223456 132368 223508
rect 181536 223456 181588 223508
rect 191196 223456 191248 223508
rect 195704 223456 195756 223508
rect 297916 222844 297968 222896
rect 349804 222844 349856 222896
rect 195428 222164 195480 222216
rect 207940 222164 207992 222216
rect 130936 222096 130988 222148
rect 163504 222096 163556 222148
rect 164148 222096 164200 222148
rect 195244 222096 195296 222148
rect 240876 222096 240928 222148
rect 164148 221484 164200 221536
rect 195244 221484 195296 221536
rect 269028 221484 269080 221536
rect 342904 221484 342956 221536
rect 194324 221416 194376 221468
rect 273904 221416 273956 221468
rect 320640 221416 320692 221468
rect 454040 221416 454092 221468
rect 276756 220804 276808 220856
rect 277400 220804 277452 220856
rect 59176 220736 59228 220788
rect 217140 220736 217192 220788
rect 195704 220668 195756 220720
rect 212448 220668 212500 220720
rect 60464 220056 60516 220108
rect 156512 220056 156564 220108
rect 192944 220056 192996 220108
rect 238760 220056 238812 220108
rect 272708 220056 272760 220108
rect 156696 219988 156748 220040
rect 211988 219444 212040 219496
rect 325056 219444 325108 219496
rect 73804 219376 73856 219428
rect 184296 219376 184348 219428
rect 195888 219376 195940 219428
rect 270500 219376 270552 219428
rect 126980 219308 127032 219360
rect 217324 219308 217376 219360
rect 221372 219308 221424 219360
rect 263784 219308 263836 219360
rect 267096 218696 267148 218748
rect 275376 218696 275428 218748
rect 192668 218016 192720 218068
rect 195244 218016 195296 218068
rect 270500 218016 270552 218068
rect 271144 218016 271196 218068
rect 83556 217948 83608 218000
rect 201500 217948 201552 218000
rect 202052 217948 202104 218000
rect 202328 217948 202380 218000
rect 231124 217948 231176 218000
rect 193036 217676 193088 217728
rect 198096 217676 198148 217728
rect 202052 217336 202104 217388
rect 285680 217336 285732 217388
rect 82728 217268 82780 217320
rect 158720 217268 158772 217320
rect 235356 217268 235408 217320
rect 388536 217268 388588 217320
rect 198004 216656 198056 216708
rect 198740 216656 198792 216708
rect 69756 216588 69808 216640
rect 233516 216588 233568 216640
rect 132408 216520 132460 216572
rect 195336 216520 195388 216572
rect 214564 216520 214616 216572
rect 248972 216520 249024 216572
rect 249708 216520 249760 216572
rect 233516 216044 233568 216096
rect 234436 216044 234488 216096
rect 249708 215908 249760 215960
rect 456800 215908 456852 215960
rect 3332 215228 3384 215280
rect 39304 215228 39356 215280
rect 124220 215228 124272 215280
rect 222384 215228 222436 215280
rect 223396 215228 223448 215280
rect 141976 215160 142028 215212
rect 168380 215160 168432 215212
rect 67640 214548 67692 214600
rect 133144 214548 133196 214600
rect 168380 214548 168432 214600
rect 169576 214548 169628 214600
rect 217416 214548 217468 214600
rect 431868 214548 431920 214600
rect 434720 214548 434772 214600
rect 223396 213936 223448 213988
rect 231952 213936 232004 213988
rect 81440 213868 81492 213920
rect 191104 213868 191156 213920
rect 213460 213868 213512 213920
rect 299572 213868 299624 213920
rect 300216 213868 300268 213920
rect 147496 213800 147548 213852
rect 244464 213800 244516 213852
rect 196716 213188 196768 213240
rect 212540 213188 212592 213240
rect 213460 213188 213512 213240
rect 254032 213188 254084 213240
rect 389824 213188 389876 213240
rect 64604 212440 64656 212492
rect 206468 212440 206520 212492
rect 136640 212372 136692 212424
rect 240140 212372 240192 212424
rect 240784 212372 240836 212424
rect 162768 211080 162820 211132
rect 163688 211080 163740 211132
rect 192484 211080 192536 211132
rect 259460 211080 259512 211132
rect 260748 211080 260800 211132
rect 212540 211012 212592 211064
rect 213644 211012 213696 211064
rect 218428 211012 218480 211064
rect 218796 211012 218848 211064
rect 274640 211012 274692 211064
rect 124312 210468 124364 210520
rect 162768 210468 162820 210520
rect 274640 210468 274692 210520
rect 290004 210468 290056 210520
rect 72516 210400 72568 210452
rect 182180 210400 182232 210452
rect 187056 210400 187108 210452
rect 212540 210400 212592 210452
rect 260748 210400 260800 210452
rect 356704 210400 356756 210452
rect 106188 209720 106240 209772
rect 216772 209720 216824 209772
rect 63408 209652 63460 209704
rect 173808 209652 173860 209704
rect 223396 209108 223448 209160
rect 282276 209108 282328 209160
rect 217416 209040 217468 209092
rect 237472 209040 237524 209092
rect 242164 209040 242216 209092
rect 251916 209040 251968 209092
rect 272708 209040 272760 209092
rect 438124 209040 438176 209092
rect 95148 208292 95200 208344
rect 193864 208292 193916 208344
rect 203524 208020 203576 208072
rect 211896 208020 211948 208072
rect 212448 207680 212500 207732
rect 235264 207680 235316 207732
rect 93952 207612 94004 207664
rect 95148 207612 95200 207664
rect 133788 207612 133840 207664
rect 229192 207612 229244 207664
rect 245844 207612 245896 207664
rect 250536 207612 250588 207664
rect 308404 207612 308456 207664
rect 114468 206932 114520 206984
rect 242900 206932 242952 206984
rect 440240 206932 440292 206984
rect 440884 206932 440936 206984
rect 582748 206932 582800 206984
rect 105544 206864 105596 206916
rect 214472 206864 214524 206916
rect 264980 206252 265032 206304
rect 371884 206252 371936 206304
rect 242900 206116 242952 206168
rect 243912 206116 243964 206168
rect 214472 205640 214524 205692
rect 216036 205640 216088 205692
rect 216128 205640 216180 205692
rect 216496 205640 216548 205692
rect 245844 205640 245896 205692
rect 97264 205572 97316 205624
rect 205824 205572 205876 205624
rect 205824 205096 205876 205148
rect 206560 205096 206612 205148
rect 87144 204892 87196 204944
rect 184664 204892 184716 204944
rect 185584 204892 185636 204944
rect 207296 204892 207348 204944
rect 280896 204892 280948 204944
rect 207020 204280 207072 204332
rect 207388 204280 207440 204332
rect 215300 204280 215352 204332
rect 70400 204212 70452 204264
rect 216128 204212 216180 204264
rect 184756 203600 184808 203652
rect 227720 203600 227772 203652
rect 102048 203532 102100 203584
rect 171784 203532 171836 203584
rect 215300 203532 215352 203584
rect 284944 203532 284996 203584
rect 3056 202784 3108 202836
rect 129004 202784 129056 202836
rect 156696 202784 156748 202836
rect 177764 202784 177816 202836
rect 207020 202784 207072 202836
rect 126888 202716 126940 202768
rect 248512 202716 248564 202768
rect 211068 202104 211120 202156
rect 240232 202104 240284 202156
rect 273996 201764 274048 201816
rect 278228 201764 278280 201816
rect 97908 201424 97960 201476
rect 165068 201424 165120 201476
rect 168288 201424 168340 201476
rect 211988 201424 212040 201476
rect 195336 200812 195388 200864
rect 218704 200812 218756 200864
rect 224316 200812 224368 200864
rect 236000 200812 236052 200864
rect 122748 200744 122800 200796
rect 178776 200744 178828 200796
rect 214656 200744 214708 200796
rect 306472 200744 306524 200796
rect 323676 200744 323728 200796
rect 431224 200744 431276 200796
rect 79968 200064 80020 200116
rect 194508 200064 194560 200116
rect 194416 199452 194468 199504
rect 287244 199452 287296 199504
rect 54944 199384 54996 199436
rect 177856 199384 177908 199436
rect 178868 199384 178920 199436
rect 194508 199384 194560 199436
rect 217324 199384 217376 199436
rect 239404 199384 239456 199436
rect 385776 199384 385828 199436
rect 53564 198636 53616 198688
rect 168288 198636 168340 198688
rect 178960 198636 179012 198688
rect 195244 198636 195296 198688
rect 139400 198568 139452 198620
rect 166908 198568 166960 198620
rect 195428 198024 195480 198076
rect 206284 198024 206336 198076
rect 206560 198024 206612 198076
rect 288624 198024 288676 198076
rect 166172 197956 166224 198008
rect 218796 197956 218848 198008
rect 220360 197956 220412 198008
rect 407120 197956 407172 198008
rect 64788 197276 64840 197328
rect 221648 197276 221700 197328
rect 221556 196664 221608 196716
rect 244372 196664 244424 196716
rect 135168 196596 135220 196648
rect 181628 196596 181680 196648
rect 189724 196596 189776 196648
rect 250444 196596 250496 196648
rect 251916 196596 251968 196648
rect 300308 196596 300360 196648
rect 155224 195916 155276 195968
rect 163504 195916 163556 195968
rect 163596 195304 163648 195356
rect 176016 195304 176068 195356
rect 177856 195304 177908 195356
rect 206560 195304 206612 195356
rect 280804 195304 280856 195356
rect 303896 195304 303948 195356
rect 89628 195236 89680 195288
rect 166356 195236 166408 195288
rect 206468 195236 206520 195288
rect 241612 195236 241664 195288
rect 270408 195236 270460 195288
rect 302240 195236 302292 195288
rect 61844 194488 61896 194540
rect 220176 194488 220228 194540
rect 223488 193876 223540 193928
rect 238760 193876 238812 193928
rect 144828 193808 144880 193860
rect 163596 193808 163648 193860
rect 198096 193808 198148 193860
rect 227076 193808 227128 193860
rect 395896 193808 395948 193860
rect 582932 193808 582984 193860
rect 226340 193196 226392 193248
rect 432696 193196 432748 193248
rect 57612 193128 57664 193180
rect 166172 193128 166224 193180
rect 93124 193060 93176 193112
rect 196716 193060 196768 193112
rect 202144 192516 202196 192568
rect 239404 192516 239456 192568
rect 185676 192448 185728 192500
rect 230664 192448 230716 192500
rect 400864 192448 400916 192500
rect 415400 192448 415452 192500
rect 200028 192380 200080 192432
rect 201500 192380 201552 192432
rect 156604 191768 156656 191820
rect 226340 191768 226392 191820
rect 221464 191088 221516 191140
rect 447324 191088 447376 191140
rect 118608 190476 118660 190528
rect 170496 190476 170548 190528
rect 159364 190408 159416 190460
rect 225604 190408 225656 190460
rect 264244 189728 264296 189780
rect 281632 189728 281684 189780
rect 122748 189048 122800 189100
rect 174544 189048 174596 189100
rect 224224 189048 224276 189100
rect 243084 189048 243136 189100
rect 2780 188844 2832 188896
rect 4804 188844 4856 188896
rect 188436 188368 188488 188420
rect 204536 188368 204588 188420
rect 206376 188368 206428 188420
rect 233424 188368 233476 188420
rect 32404 188300 32456 188352
rect 159364 188300 159416 188352
rect 162768 188300 162820 188352
rect 177580 188300 177632 188352
rect 201500 188300 201552 188352
rect 249800 188300 249852 188352
rect 268384 188300 268436 188352
rect 296904 188300 296956 188352
rect 300308 188300 300360 188352
rect 310704 188300 310756 188352
rect 125508 187688 125560 187740
rect 202144 187688 202196 187740
rect 282184 187144 282236 187196
rect 284576 187144 284628 187196
rect 191748 186940 191800 186992
rect 235356 186940 235408 186992
rect 126888 186396 126940 186448
rect 164884 186396 164936 186448
rect 110328 186328 110380 186380
rect 187148 186328 187200 186380
rect 204536 186260 204588 186312
rect 224224 186260 224276 186312
rect 191104 185648 191156 185700
rect 204996 185648 205048 185700
rect 215300 185648 215352 185700
rect 227812 185648 227864 185700
rect 181536 185580 181588 185632
rect 216036 185580 216088 185632
rect 226340 185580 226392 185632
rect 249892 185580 249944 185632
rect 267004 185580 267056 185632
rect 279148 185580 279200 185632
rect 130936 184968 130988 185020
rect 169208 184968 169260 185020
rect 148876 184900 148928 184952
rect 191104 184900 191156 184952
rect 272432 184900 272484 184952
rect 302424 184900 302476 184952
rect 207020 184832 207072 184884
rect 226340 184832 226392 184884
rect 271236 184832 271288 184884
rect 279608 184832 279660 184884
rect 196624 184152 196676 184204
rect 231124 184152 231176 184204
rect 257436 184152 257488 184204
rect 280252 184152 280304 184204
rect 334808 184152 334860 184204
rect 396908 184152 396960 184204
rect 133788 183608 133840 183660
rect 162124 183608 162176 183660
rect 124864 183540 124916 183592
rect 200764 183540 200816 183592
rect 224316 182860 224368 182912
rect 232044 182860 232096 182912
rect 180708 182792 180760 182844
rect 215116 182792 215168 182844
rect 215944 182792 215996 182844
rect 241520 182792 241572 182844
rect 270316 182792 270368 182844
rect 303804 182792 303856 182844
rect 114376 182248 114428 182300
rect 164976 182248 165028 182300
rect 103336 182180 103388 182232
rect 171876 182180 171928 182232
rect 211896 182112 211948 182164
rect 272432 182112 272484 182164
rect 269856 181500 269908 181552
rect 283104 181500 283156 181552
rect 273904 181432 273956 181484
rect 294052 181432 294104 181484
rect 124036 180888 124088 180940
rect 166540 180888 166592 180940
rect 132408 180820 132460 180872
rect 211804 180820 211856 180872
rect 226984 180820 227036 180872
rect 229284 180820 229336 180872
rect 204996 180752 205048 180804
rect 218796 180752 218848 180804
rect 260104 180140 260156 180192
rect 285864 180140 285916 180192
rect 220084 180072 220136 180124
rect 234712 180072 234764 180124
rect 262864 180072 262916 180124
rect 291384 180072 291436 180124
rect 119528 179460 119580 179512
rect 198096 179460 198148 179512
rect 129464 179392 129516 179444
rect 214196 179392 214248 179444
rect 215944 179392 215996 179444
rect 230848 179392 230900 179444
rect 230388 179324 230440 179376
rect 258080 179324 258132 179376
rect 259276 179324 259328 179376
rect 215116 178712 215168 178764
rect 240324 178712 240376 178764
rect 271144 178712 271196 178764
rect 283012 178712 283064 178764
rect 283564 178712 283616 178764
rect 298192 178712 298244 178764
rect 177948 178644 178000 178696
rect 229560 178644 229612 178696
rect 262128 178644 262180 178696
rect 280344 178644 280396 178696
rect 280896 178644 280948 178696
rect 299572 178644 299624 178696
rect 115848 178100 115900 178152
rect 170588 178100 170640 178152
rect 113732 178032 113784 178084
rect 177488 178032 177540 178084
rect 120816 177964 120868 178016
rect 124864 177964 124916 178016
rect 275468 177964 275520 178016
rect 284300 177964 284352 178016
rect 282276 177896 282328 177948
rect 288716 177896 288768 177948
rect 226340 177556 226392 177608
rect 230572 177556 230624 177608
rect 181628 177352 181680 177404
rect 207664 177352 207716 177404
rect 284944 177352 284996 177404
rect 289820 177352 289872 177404
rect 181444 177284 181496 177336
rect 234620 177284 234672 177336
rect 235264 177284 235316 177336
rect 243176 177284 243228 177336
rect 276756 177284 276808 177336
rect 280804 177284 280856 177336
rect 298744 177284 298796 177336
rect 371976 177284 372028 177336
rect 158996 176740 159048 176792
rect 166264 176740 166316 176792
rect 127072 176672 127124 176724
rect 165436 176672 165488 176724
rect 231124 176672 231176 176724
rect 231860 176672 231912 176724
rect 135720 176604 135772 176656
rect 213920 176604 213972 176656
rect 228364 175992 228416 176044
rect 234804 175992 234856 176044
rect 134432 175924 134484 175976
rect 165528 175924 165580 175976
rect 218704 175924 218756 175976
rect 233240 175924 233292 175976
rect 239404 175924 239456 175976
rect 281908 175924 281960 175976
rect 305184 175924 305236 175976
rect 316132 175924 316184 175976
rect 333888 175924 333940 175976
rect 401692 175924 401744 175976
rect 278228 175788 278280 175840
rect 279332 175788 279384 175840
rect 215392 175244 215444 175296
rect 229008 175244 229060 175296
rect 239496 175244 239548 175296
rect 264980 175244 265032 175296
rect 281540 175244 281592 175296
rect 305184 175244 305236 175296
rect 305644 175244 305696 175296
rect 162124 175176 162176 175228
rect 214012 175176 214064 175228
rect 230480 175176 230532 175228
rect 244924 175176 244976 175228
rect 281816 175176 281868 175228
rect 305276 175176 305328 175228
rect 165528 175108 165580 175160
rect 213920 175108 213972 175160
rect 229100 174564 229152 174616
rect 229284 174564 229336 174616
rect 215300 173884 215352 173936
rect 229008 173952 229060 174004
rect 230020 173952 230072 174004
rect 230940 173952 230992 174004
rect 245016 173952 245068 174004
rect 264980 173952 265032 174004
rect 238208 173884 238260 173936
rect 265072 173884 265124 173936
rect 169208 173816 169260 173868
rect 213920 173816 213972 173868
rect 211804 173748 211856 173800
rect 214472 173748 214524 173800
rect 231676 173136 231728 173188
rect 244464 173136 244516 173188
rect 300124 173136 300176 173188
rect 419632 173136 419684 173188
rect 250536 172592 250588 172644
rect 265072 172592 265124 172644
rect 236920 172524 236972 172576
rect 264980 172524 265032 172576
rect 166356 172456 166408 172508
rect 215300 172456 215352 172508
rect 231400 172456 231452 172508
rect 248604 172456 248656 172508
rect 190368 172388 190420 172440
rect 216772 172388 216824 172440
rect 231768 172388 231820 172440
rect 242992 172388 243044 172440
rect 254584 171164 254636 171216
rect 265072 171164 265124 171216
rect 249340 171096 249392 171148
rect 264980 171096 265032 171148
rect 289820 171776 289872 171828
rect 354128 171776 354180 171828
rect 417424 171776 417476 171828
rect 164884 171028 164936 171080
rect 213920 171028 213972 171080
rect 210516 170960 210568 171012
rect 214012 170960 214064 171012
rect 280068 170892 280120 170944
rect 230756 170620 230808 170672
rect 233240 170620 233292 170672
rect 231124 170348 231176 170400
rect 247040 170348 247092 170400
rect 342996 170348 343048 170400
rect 392768 170348 392820 170400
rect 247684 169804 247736 169856
rect 264980 169804 265032 169856
rect 240876 169736 240928 169788
rect 265072 169736 265124 169788
rect 166540 169668 166592 169720
rect 214012 169668 214064 169720
rect 281540 169668 281592 169720
rect 284668 169668 284720 169720
rect 202144 169600 202196 169652
rect 213920 169600 213972 169652
rect 231768 169532 231820 169584
rect 236000 169532 236052 169584
rect 231768 169124 231820 169176
rect 234712 169124 234764 169176
rect 242256 168444 242308 168496
rect 264980 168444 265032 168496
rect 235264 168376 235316 168428
rect 265072 168376 265124 168428
rect 174544 168308 174596 168360
rect 213920 168308 213972 168360
rect 231492 168308 231544 168360
rect 234804 168308 234856 168360
rect 200764 168240 200816 168292
rect 214012 168240 214064 168292
rect 234712 167968 234764 168020
rect 237380 167968 237432 168020
rect 308404 167628 308456 167680
rect 434720 167628 434772 167680
rect 262956 167084 263008 167136
rect 265348 167084 265400 167136
rect 233976 167016 234028 167068
rect 264980 167016 265032 167068
rect 170496 166948 170548 167000
rect 214012 166948 214064 167000
rect 281908 166948 281960 167000
rect 291476 166948 291528 167000
rect 198096 166880 198148 166932
rect 213920 166880 213972 166932
rect 231308 166880 231360 166932
rect 234620 166880 234672 166932
rect 231768 166676 231820 166728
rect 234712 166676 234764 166728
rect 249064 165656 249116 165708
rect 265072 165656 265124 165708
rect 237012 165588 237064 165640
rect 264980 165588 265032 165640
rect 170588 165520 170640 165572
rect 213920 165520 213972 165572
rect 231492 165180 231544 165232
rect 234620 165180 234672 165232
rect 230940 165112 230992 165164
rect 233332 165112 233384 165164
rect 282184 164908 282236 164960
rect 310704 164908 310756 164960
rect 300216 164840 300268 164892
rect 381728 164840 381780 164892
rect 257344 164296 257396 164348
rect 264980 164296 265032 164348
rect 247776 164228 247828 164280
rect 265072 164228 265124 164280
rect 282828 164228 282880 164280
rect 287244 164228 287296 164280
rect 3332 164160 3384 164212
rect 29644 164160 29696 164212
rect 176108 164160 176160 164212
rect 214012 164160 214064 164212
rect 231032 164160 231084 164212
rect 248420 164160 248472 164212
rect 177488 164092 177540 164144
rect 213920 164092 213972 164144
rect 167828 163480 167880 163532
rect 175924 163480 175976 163532
rect 245108 163480 245160 163532
rect 265440 163480 265492 163532
rect 281816 163480 281868 163532
rect 295340 163480 295392 163532
rect 341616 163480 341668 163532
rect 444564 163480 444616 163532
rect 282828 163072 282880 163124
rect 288716 163072 288768 163124
rect 252192 162868 252244 162920
rect 265072 162868 265124 162920
rect 166448 162800 166500 162852
rect 213920 162800 213972 162852
rect 242440 162800 242492 162852
rect 243084 162800 243136 162852
rect 243544 162800 243596 162852
rect 244372 162800 244424 162852
rect 281632 162800 281684 162852
rect 303896 162800 303948 162852
rect 187148 162732 187200 162784
rect 214012 162732 214064 162784
rect 231676 162732 231728 162784
rect 241612 162732 241664 162784
rect 256148 162120 256200 162172
rect 264980 162120 265032 162172
rect 281908 161780 281960 161832
rect 286324 161780 286376 161832
rect 235540 161440 235592 161492
rect 265072 161440 265124 161492
rect 165528 161372 165580 161424
rect 214012 161372 214064 161424
rect 282828 161372 282880 161424
rect 317512 161372 317564 161424
rect 173348 161304 173400 161356
rect 213920 161304 213972 161356
rect 231032 161032 231084 161084
rect 233516 161032 233568 161084
rect 249708 160692 249760 160744
rect 262956 160692 263008 160744
rect 356796 160692 356848 160744
rect 395436 160692 395488 160744
rect 282828 160420 282880 160472
rect 287336 160420 287388 160472
rect 263048 160148 263100 160200
rect 265440 160148 265492 160200
rect 229744 160080 229796 160132
rect 231952 160080 232004 160132
rect 245200 160080 245252 160132
rect 264980 160080 265032 160132
rect 167644 160012 167696 160064
rect 213920 160012 213972 160064
rect 282828 160012 282880 160064
rect 293960 160012 294012 160064
rect 230572 159400 230624 159452
rect 240232 159400 240284 159452
rect 232688 159332 232740 159384
rect 265256 159332 265308 159384
rect 307116 159332 307168 159384
rect 409972 159332 410024 159384
rect 241060 158720 241112 158772
rect 264980 158720 265032 158772
rect 171876 158652 171928 158704
rect 213920 158652 213972 158704
rect 231768 158652 231820 158704
rect 241704 158652 241756 158704
rect 282092 158652 282144 158704
rect 292764 158652 292816 158704
rect 180248 158584 180300 158636
rect 214012 158584 214064 158636
rect 231492 158584 231544 158636
rect 234252 158584 234304 158636
rect 322296 157972 322348 158024
rect 430580 157972 430632 158024
rect 242164 157428 242216 157480
rect 264980 157428 265032 157480
rect 238300 157360 238352 157412
rect 265072 157360 265124 157412
rect 281540 157360 281592 157412
rect 283196 157360 283248 157412
rect 169116 157292 169168 157344
rect 213920 157292 213972 157344
rect 231768 157292 231820 157344
rect 244280 157292 244332 157344
rect 180156 157224 180208 157276
rect 214012 157224 214064 157276
rect 318064 156612 318116 156664
rect 422300 156612 422352 156664
rect 250628 156000 250680 156052
rect 265072 156000 265124 156052
rect 246304 155932 246356 155984
rect 264980 155932 265032 155984
rect 170404 155864 170456 155916
rect 214012 155864 214064 155916
rect 231768 155864 231820 155916
rect 238760 155864 238812 155916
rect 282276 155864 282328 155916
rect 311992 155864 312044 155916
rect 178868 155796 178920 155848
rect 213920 155796 213972 155848
rect 239680 155184 239732 155236
rect 249708 155184 249760 155236
rect 358084 155184 358136 155236
rect 436836 155184 436888 155236
rect 250444 154640 250496 154692
rect 264980 154640 265032 154692
rect 233884 154572 233936 154624
rect 265072 154572 265124 154624
rect 282828 154504 282880 154556
rect 306472 154504 306524 154556
rect 282092 154436 282144 154488
rect 302240 154436 302292 154488
rect 230664 153824 230716 153876
rect 245844 153824 245896 153876
rect 309784 153824 309836 153876
rect 423036 153824 423088 153876
rect 231216 153688 231268 153740
rect 233424 153688 233476 153740
rect 211896 153280 211948 153332
rect 214012 153280 214064 153332
rect 195428 153212 195480 153264
rect 213920 153212 213972 153264
rect 253204 153212 253256 153264
rect 264980 153212 265032 153264
rect 230480 152464 230532 152516
rect 238852 152464 238904 152516
rect 319444 152464 319496 152516
rect 441804 152464 441856 152516
rect 211988 152056 212040 152108
rect 214012 152056 214064 152108
rect 249248 151852 249300 151904
rect 265072 151852 265124 151904
rect 202236 151784 202288 151836
rect 213920 151784 213972 151836
rect 238116 151784 238168 151836
rect 264980 151784 265032 151836
rect 281908 151716 281960 151768
rect 300860 151716 300912 151768
rect 230480 151580 230532 151632
rect 232136 151580 232188 151632
rect 238392 151104 238444 151156
rect 263048 151104 263100 151156
rect 374736 151104 374788 151156
rect 429936 151104 429988 151156
rect 436744 151104 436796 151156
rect 448612 151104 448664 151156
rect 229928 151036 229980 151088
rect 265716 151036 265768 151088
rect 282276 151036 282328 151088
rect 289912 151036 289964 151088
rect 398748 151036 398800 151088
rect 583024 151036 583076 151088
rect 198096 150492 198148 150544
rect 214012 150492 214064 150544
rect 180340 150424 180392 150476
rect 213920 150424 213972 150476
rect 262956 150424 263008 150476
rect 265348 150424 265400 150476
rect 3608 150356 3660 150408
rect 11704 150356 11756 150408
rect 175924 150356 175976 150408
rect 214012 150356 214064 150408
rect 282736 150356 282788 150408
rect 307852 150356 307904 150408
rect 191104 150288 191156 150340
rect 213920 150288 213972 150340
rect 282828 150288 282880 150340
rect 302424 150288 302476 150340
rect 239404 149676 239456 149728
rect 265624 149676 265676 149728
rect 367744 149676 367796 149728
rect 439596 149676 439648 149728
rect 235448 149064 235500 149116
rect 264980 149064 265032 149116
rect 166264 148996 166316 149048
rect 213920 148996 213972 149048
rect 282828 148996 282880 149048
rect 310612 148996 310664 149048
rect 449900 148996 449952 149048
rect 582840 148996 582892 149048
rect 282184 148928 282236 148980
rect 288532 148928 288584 148980
rect 429844 148384 429896 148436
rect 440424 148384 440476 148436
rect 231124 148316 231176 148368
rect 240876 148316 240928 148368
rect 437664 148316 437716 148368
rect 449900 148316 449952 148368
rect 240968 147704 241020 147756
rect 264980 147704 265032 147756
rect 209228 147636 209280 147688
rect 213920 147636 213972 147688
rect 234068 147636 234120 147688
rect 265072 147636 265124 147688
rect 281724 147568 281776 147620
rect 299572 147568 299624 147620
rect 282828 147500 282880 147552
rect 291384 147500 291436 147552
rect 432696 146956 432748 147008
rect 443276 146956 443328 147008
rect 580908 146956 580960 147008
rect 582748 146956 582800 147008
rect 169024 146888 169076 146940
rect 204996 146888 205048 146940
rect 231860 146888 231912 146940
rect 248512 146888 248564 146940
rect 298836 146888 298888 146940
rect 404728 146888 404780 146940
rect 414664 146888 414716 146940
rect 436376 146888 436428 146940
rect 441804 146820 441856 146872
rect 441988 146820 442040 146872
rect 263048 146344 263100 146396
rect 265164 146344 265216 146396
rect 169116 146276 169168 146328
rect 213920 146276 213972 146328
rect 240876 146276 240928 146328
rect 265072 146276 265124 146328
rect 282828 146208 282880 146260
rect 302332 146208 302384 146260
rect 403624 146208 403676 146260
rect 411904 146208 411956 146260
rect 412548 146208 412600 146260
rect 414480 146208 414532 146260
rect 392584 145528 392636 145580
rect 407304 145528 407356 145580
rect 421472 145528 421524 145580
rect 582564 145528 582616 145580
rect 235356 144984 235408 145036
rect 264980 144984 265032 145036
rect 185676 144916 185728 144968
rect 213920 144916 213972 144968
rect 232872 144916 232924 144968
rect 265072 144916 265124 144968
rect 295984 144916 296036 144968
rect 403440 144916 403492 144968
rect 231768 144848 231820 144900
rect 240784 144848 240836 144900
rect 282828 144848 282880 144900
rect 294052 144848 294104 144900
rect 417424 144848 417476 144900
rect 418068 144848 418120 144900
rect 583300 144848 583352 144900
rect 170404 144168 170456 144220
rect 214012 144168 214064 144220
rect 247868 144168 247920 144220
rect 265164 144168 265216 144220
rect 280896 144168 280948 144220
rect 296812 144168 296864 144220
rect 338764 144168 338816 144220
rect 441712 144168 441764 144220
rect 171876 143556 171928 143608
rect 213920 143556 213972 143608
rect 249156 143556 249208 143608
rect 264980 143556 265032 143608
rect 300860 143488 300912 143540
rect 301504 143488 301556 143540
rect 405004 143488 405056 143540
rect 409052 143488 409104 143540
rect 418896 143488 418948 143540
rect 420000 143488 420052 143540
rect 436836 143488 436888 143540
rect 439320 143488 439372 143540
rect 231768 142808 231820 142860
rect 241520 142808 241572 142860
rect 244280 142808 244332 142860
rect 264980 142808 265032 142860
rect 422944 142808 422996 142860
rect 432236 142808 432288 142860
rect 191104 142196 191156 142248
rect 214012 142196 214064 142248
rect 396724 142196 396776 142248
rect 414204 142196 414256 142248
rect 173256 142128 173308 142180
rect 213920 142128 213972 142180
rect 257620 142128 257672 142180
rect 265072 142128 265124 142180
rect 300860 142128 300912 142180
rect 402612 142128 402664 142180
rect 428464 142128 428516 142180
rect 432880 142128 432932 142180
rect 583024 142128 583076 142180
rect 282828 142060 282880 142112
rect 295524 142060 295576 142112
rect 281908 141720 281960 141772
rect 285864 141720 285916 141772
rect 247960 141448 248012 141500
rect 265808 141448 265860 141500
rect 173164 141380 173216 141432
rect 184296 141380 184348 141432
rect 232596 141380 232648 141432
rect 265164 141380 265216 141432
rect 319444 141380 319496 141432
rect 416780 141380 416832 141432
rect 431224 141380 431276 141432
rect 440332 141380 440384 141432
rect 198188 140836 198240 140888
rect 213920 140836 213972 140888
rect 317420 140836 317472 140888
rect 191288 140768 191340 140820
rect 214012 140768 214064 140820
rect 422576 140836 422628 140888
rect 423036 140836 423088 140888
rect 423680 140768 423732 140820
rect 424508 140768 424560 140820
rect 580264 140768 580316 140820
rect 282736 140700 282788 140752
rect 318800 140700 318852 140752
rect 400220 140700 400272 140752
rect 400956 140700 401008 140752
rect 434720 140700 434772 140752
rect 435180 140700 435232 140752
rect 436100 140700 436152 140752
rect 437020 140700 437072 140752
rect 192484 140020 192536 140072
rect 214196 140020 214248 140072
rect 307116 140020 307168 140072
rect 317696 140020 317748 140072
rect 318708 140020 318760 140072
rect 420276 140020 420328 140072
rect 440240 140020 440292 140072
rect 282828 139544 282880 139596
rect 288440 139544 288492 139596
rect 399852 139544 399904 139596
rect 400404 139544 400456 139596
rect 231216 139476 231268 139528
rect 236920 139476 236972 139528
rect 398012 139476 398064 139528
rect 404360 139476 404412 139528
rect 174544 139408 174596 139460
rect 213920 139408 213972 139460
rect 231400 139408 231452 139460
rect 235264 139408 235316 139460
rect 248052 139408 248104 139460
rect 264980 139408 265032 139460
rect 318708 139408 318760 139460
rect 417148 139408 417200 139460
rect 426808 139408 426860 139460
rect 582656 139408 582708 139460
rect 231768 139340 231820 139392
rect 255412 139340 255464 139392
rect 282828 139340 282880 139392
rect 296904 139340 296956 139392
rect 398104 139340 398156 139392
rect 412732 139340 412784 139392
rect 438216 139340 438268 139392
rect 439504 139340 439556 139392
rect 231308 138796 231360 138848
rect 238208 138796 238260 138848
rect 178776 138660 178828 138712
rect 200764 138660 200816 138712
rect 263140 138048 263192 138100
rect 265072 138048 265124 138100
rect 322296 138048 322348 138100
rect 398104 138048 398156 138100
rect 175924 137980 175976 138032
rect 213920 137980 213972 138032
rect 238024 137980 238076 138032
rect 264980 137980 265032 138032
rect 398656 137980 398708 138032
rect 580172 137980 580224 138032
rect 3332 137912 3384 137964
rect 21364 137912 21416 137964
rect 231584 137912 231636 137964
rect 249800 137912 249852 137964
rect 281632 137912 281684 137964
rect 300952 137912 301004 137964
rect 327724 137912 327776 137964
rect 397552 137912 397604 137964
rect 170680 137232 170732 137284
rect 214380 137232 214432 137284
rect 264520 137232 264572 137284
rect 265624 137232 265676 137284
rect 442908 136688 442960 136740
rect 452752 136688 452804 136740
rect 229744 136620 229796 136672
rect 264980 136620 265032 136672
rect 388444 136620 388496 136672
rect 397552 136620 397604 136672
rect 440424 136620 440476 136672
rect 582564 136620 582616 136672
rect 231492 136552 231544 136604
rect 245016 136552 245068 136604
rect 395436 136552 395488 136604
rect 397644 136552 397696 136604
rect 441988 136552 442040 136604
rect 583392 136552 583444 136604
rect 231768 136484 231820 136536
rect 242992 136484 243044 136536
rect 282276 136008 282328 136060
rect 285680 136008 285732 136060
rect 328368 135872 328420 135924
rect 398012 135872 398064 135924
rect 182916 135328 182968 135380
rect 213920 135328 213972 135380
rect 250812 135328 250864 135380
rect 265072 135328 265124 135380
rect 177488 135260 177540 135312
rect 214012 135260 214064 135312
rect 243544 135260 243596 135312
rect 264980 135260 265032 135312
rect 231492 135192 231544 135244
rect 250536 135192 250588 135244
rect 363604 135192 363656 135244
rect 398656 135192 398708 135244
rect 230756 135056 230808 135108
rect 237012 135056 237064 135108
rect 178684 134580 178736 134632
rect 199476 134580 199528 134632
rect 185584 134512 185636 134564
rect 214104 134512 214156 134564
rect 250720 134512 250772 134564
rect 265256 134512 265308 134564
rect 442908 134512 442960 134564
rect 443092 134512 443144 134564
rect 456892 134512 456944 134564
rect 202144 133900 202196 133952
rect 213920 133900 213972 133952
rect 260196 133900 260248 133952
rect 264980 133900 265032 133952
rect 376116 133900 376168 133952
rect 397552 133900 397604 133952
rect 231676 133832 231728 133884
rect 254584 133832 254636 133884
rect 282828 133832 282880 133884
rect 313372 133832 313424 133884
rect 342904 133832 342956 133884
rect 397644 133832 397696 133884
rect 442908 133832 442960 133884
rect 582472 133832 582524 133884
rect 231768 133764 231820 133816
rect 253296 133764 253348 133816
rect 171784 133152 171836 133204
rect 206468 133152 206520 133204
rect 211804 132540 211856 132592
rect 214472 132540 214524 132592
rect 196808 132472 196860 132524
rect 213920 132472 213972 132524
rect 253572 132472 253624 132524
rect 264980 132472 265032 132524
rect 231768 132404 231820 132456
rect 249340 132404 249392 132456
rect 282644 132404 282696 132456
rect 325700 132404 325752 132456
rect 369124 132404 369176 132456
rect 397552 132404 397604 132456
rect 281724 132336 281776 132388
rect 303620 132336 303672 132388
rect 178776 131724 178828 131776
rect 211988 131724 212040 131776
rect 231676 131724 231728 131776
rect 239680 131724 239732 131776
rect 256700 131724 256752 131776
rect 265164 131724 265216 131776
rect 180248 131112 180300 131164
rect 213920 131112 213972 131164
rect 252008 131112 252060 131164
rect 264980 131112 265032 131164
rect 231768 131044 231820 131096
rect 260104 131044 260156 131096
rect 282276 131044 282328 131096
rect 316040 131044 316092 131096
rect 231400 130976 231452 131028
rect 247684 130976 247736 131028
rect 282828 130976 282880 131028
rect 303804 130976 303856 131028
rect 442908 130772 442960 130824
rect 444380 130772 444432 130824
rect 192576 130432 192628 130484
rect 214472 130432 214524 130484
rect 180156 130364 180208 130416
rect 209228 130364 209280 130416
rect 345756 130364 345808 130416
rect 391204 130364 391256 130416
rect 209136 129752 209188 129804
rect 213920 129752 213972 129804
rect 256056 129752 256108 129804
rect 264980 129752 265032 129804
rect 355324 129752 355376 129804
rect 358820 129752 358872 129804
rect 397552 129752 397604 129804
rect 442908 129752 442960 129804
rect 454132 129752 454184 129804
rect 231768 129684 231820 129736
rect 252100 129684 252152 129736
rect 282092 129684 282144 129736
rect 288624 129684 288676 129736
rect 231400 129616 231452 129668
rect 242256 129616 242308 129668
rect 367836 129072 367888 129124
rect 393320 129072 393372 129124
rect 394608 129072 394660 129124
rect 167736 129004 167788 129056
rect 198096 129004 198148 129056
rect 336004 129004 336056 129056
rect 378876 129004 378928 129056
rect 257528 128392 257580 128444
rect 265072 128392 265124 128444
rect 60648 128324 60700 128376
rect 66168 128324 66220 128376
rect 210608 128324 210660 128376
rect 213920 128324 213972 128376
rect 251916 128324 251968 128376
rect 264980 128324 265032 128376
rect 393964 128324 394016 128376
rect 397552 128324 397604 128376
rect 442172 128324 442224 128376
rect 444472 128324 444524 128376
rect 231768 128256 231820 128308
rect 245108 128256 245160 128308
rect 231308 127984 231360 128036
rect 233976 127984 234028 128036
rect 285680 127644 285732 127696
rect 295984 127644 296036 127696
rect 173348 127576 173400 127628
rect 214564 127576 214616 127628
rect 282828 127576 282880 127628
rect 314660 127576 314712 127628
rect 442908 127168 442960 127220
rect 448520 127168 448572 127220
rect 261484 127032 261536 127084
rect 265072 127032 265124 127084
rect 187148 126964 187200 127016
rect 213920 126964 213972 127016
rect 242256 126964 242308 127016
rect 264980 126964 265032 127016
rect 371884 126964 371936 127016
rect 397552 126964 397604 127016
rect 231676 126896 231728 126948
rect 249064 126896 249116 126948
rect 282276 126896 282328 126948
rect 298192 126896 298244 126948
rect 371240 126896 371292 126948
rect 398104 126896 398156 126948
rect 442908 126896 442960 126948
rect 583116 126896 583168 126948
rect 231768 126828 231820 126880
rect 243636 126828 243688 126880
rect 442816 126828 442868 126880
rect 454040 126828 454092 126880
rect 169024 126216 169076 126268
rect 211896 126216 211948 126268
rect 243728 126216 243780 126268
rect 256700 126216 256752 126268
rect 260380 126216 260432 126268
rect 263140 126216 263192 126268
rect 282000 126216 282052 126268
rect 306380 126216 306432 126268
rect 202420 125604 202472 125656
rect 213920 125604 213972 125656
rect 257436 125604 257488 125656
rect 264980 125604 265032 125656
rect 282368 125536 282420 125588
rect 298100 125536 298152 125588
rect 442908 125536 442960 125588
rect 460940 125536 460992 125588
rect 582748 125536 582800 125588
rect 230756 124924 230808 124976
rect 250628 124924 250680 124976
rect 205088 124856 205140 124908
rect 214012 124856 214064 124908
rect 230664 124856 230716 124908
rect 245200 124856 245252 124908
rect 245292 124856 245344 124908
rect 265716 124856 265768 124908
rect 166264 124176 166316 124228
rect 213920 124176 213972 124228
rect 254768 124176 254820 124228
rect 264980 124176 265032 124228
rect 377404 124176 377456 124228
rect 385040 124176 385092 124228
rect 397552 124176 397604 124228
rect 231768 124108 231820 124160
rect 252192 124108 252244 124160
rect 385684 124108 385736 124160
rect 397644 124108 397696 124160
rect 442632 124108 442684 124160
rect 583484 124108 583536 124160
rect 230572 124040 230624 124092
rect 232688 124040 232740 124092
rect 167644 123428 167696 123480
rect 180340 123428 180392 123480
rect 232780 123428 232832 123480
rect 248052 123428 248104 123480
rect 282736 123428 282788 123480
rect 291292 123428 291344 123480
rect 354036 123428 354088 123480
rect 397552 123428 397604 123480
rect 196716 122884 196768 122936
rect 214012 122884 214064 122936
rect 252100 122884 252152 122936
rect 264980 122884 265032 122936
rect 176016 122816 176068 122868
rect 213920 122816 213972 122868
rect 250812 122816 250864 122868
rect 265072 122816 265124 122868
rect 231768 122748 231820 122800
rect 256148 122748 256200 122800
rect 282828 122748 282880 122800
rect 305000 122748 305052 122800
rect 441896 122612 441948 122664
rect 444564 122612 444616 122664
rect 230940 121864 230992 121916
rect 235540 121864 235592 121916
rect 180340 121524 180392 121576
rect 213920 121524 213972 121576
rect 171784 121456 171836 121508
rect 214012 121456 214064 121508
rect 249064 121456 249116 121508
rect 264980 121456 265032 121508
rect 367744 121456 367796 121508
rect 397552 121456 397604 121508
rect 231676 121388 231728 121440
rect 260288 121388 260340 121440
rect 282828 121388 282880 121440
rect 290004 121388 290056 121440
rect 387064 121388 387116 121440
rect 397644 121388 397696 121440
rect 231768 121320 231820 121372
rect 240784 121320 240836 121372
rect 191196 120164 191248 120216
rect 214012 120164 214064 120216
rect 260104 120164 260156 120216
rect 265072 120164 265124 120216
rect 166356 120096 166408 120148
rect 213920 120096 213972 120148
rect 262772 120096 262824 120148
rect 264980 120096 265032 120148
rect 231768 120028 231820 120080
rect 241060 120028 241112 120080
rect 282828 120028 282880 120080
rect 292580 120028 292632 120080
rect 338856 120028 338908 120080
rect 397644 120028 397696 120080
rect 385776 119960 385828 120012
rect 397552 119960 397604 120012
rect 231032 119892 231084 119944
rect 238300 119892 238352 119944
rect 240876 119348 240928 119400
rect 258908 119348 258960 119400
rect 192576 118736 192628 118788
rect 213920 118736 213972 118788
rect 258724 118736 258776 118788
rect 265072 118736 265124 118788
rect 174636 118668 174688 118720
rect 214012 118668 214064 118720
rect 240784 118668 240836 118720
rect 264980 118668 265032 118720
rect 231768 118600 231820 118652
rect 267280 118600 267332 118652
rect 352656 118600 352708 118652
rect 397552 118600 397604 118652
rect 442908 118532 442960 118584
rect 445852 118532 445904 118584
rect 230940 118396 230992 118448
rect 236736 118396 236788 118448
rect 282552 118396 282604 118448
rect 285772 118396 285824 118448
rect 177396 117988 177448 118040
rect 188344 117988 188396 118040
rect 173164 117920 173216 117972
rect 191104 117920 191156 117972
rect 236920 117920 236972 117972
rect 248420 117920 248472 117972
rect 282184 117920 282236 117972
rect 296720 117920 296772 117972
rect 338120 117512 338172 117564
rect 340236 117512 340288 117564
rect 198096 117376 198148 117428
rect 213920 117376 213972 117428
rect 194048 117308 194100 117360
rect 214012 117308 214064 117360
rect 253480 117308 253532 117360
rect 264980 117308 265032 117360
rect 374736 117308 374788 117360
rect 397644 117308 397696 117360
rect 231492 117240 231544 117292
rect 242164 117240 242216 117292
rect 320916 117240 320968 117292
rect 395896 117240 395948 117292
rect 397552 117240 397604 117292
rect 235540 116560 235592 116612
rect 253572 116560 253624 116612
rect 282276 116560 282328 116612
rect 307760 116560 307812 116612
rect 442908 116288 442960 116340
rect 449900 116288 449952 116340
rect 282828 116084 282880 116136
rect 287152 116084 287204 116136
rect 188436 116016 188488 116068
rect 213920 116016 213972 116068
rect 170588 115948 170640 116000
rect 214012 115948 214064 116000
rect 253296 115948 253348 116000
rect 264980 115948 265032 116000
rect 231492 115880 231544 115932
rect 246488 115880 246540 115932
rect 282460 115880 282512 115932
rect 309140 115880 309192 115932
rect 358176 115880 358228 115932
rect 397552 115880 397604 115932
rect 392676 115812 392728 115864
rect 397644 115812 397696 115864
rect 442908 115812 442960 115864
rect 447324 115812 447376 115864
rect 230664 114928 230716 114980
rect 233884 114928 233936 114980
rect 195336 114588 195388 114640
rect 213920 114588 213972 114640
rect 250536 114588 250588 114640
rect 265072 114588 265124 114640
rect 169208 114520 169260 114572
rect 214012 114520 214064 114572
rect 242164 114520 242216 114572
rect 264980 114520 265032 114572
rect 231768 114452 231820 114504
rect 250444 114452 250496 114504
rect 282828 114452 282880 114504
rect 290096 114452 290148 114504
rect 352564 114452 352616 114504
rect 397552 114452 397604 114504
rect 231676 114384 231728 114436
rect 243820 114384 243872 114436
rect 384304 114384 384356 114436
rect 397644 114384 397696 114436
rect 177580 113840 177632 113892
rect 202144 113840 202196 113892
rect 164884 113772 164936 113824
rect 214748 113772 214800 113824
rect 442908 113364 442960 113416
rect 444380 113364 444432 113416
rect 207756 113160 207808 113212
rect 213920 113160 213972 113212
rect 245108 113160 245160 113212
rect 264980 113160 265032 113212
rect 231768 113092 231820 113144
rect 264428 113092 264480 113144
rect 282828 113092 282880 113144
rect 303712 113092 303764 113144
rect 309876 113092 309928 113144
rect 397552 113092 397604 113144
rect 442908 113092 442960 113144
rect 456800 113092 456852 113144
rect 230940 113024 230992 113076
rect 253204 113024 253256 113076
rect 281816 113024 281868 113076
rect 284484 113024 284536 113076
rect 388536 112412 388588 112464
rect 398748 112412 398800 112464
rect 202604 111868 202656 111920
rect 214012 111868 214064 111920
rect 166540 111800 166592 111852
rect 213920 111800 213972 111852
rect 261576 111800 261628 111852
rect 264980 111800 265032 111852
rect 3148 111732 3200 111784
rect 32404 111732 32456 111784
rect 231768 111732 231820 111784
rect 249248 111732 249300 111784
rect 378784 111732 378836 111784
rect 397460 111732 397512 111784
rect 282828 111528 282880 111580
rect 287060 111528 287112 111580
rect 281540 111392 281592 111444
rect 284576 111392 284628 111444
rect 230756 110848 230808 110900
rect 238116 110848 238168 110900
rect 181628 110508 181680 110560
rect 213920 110508 213972 110560
rect 256240 110508 256292 110560
rect 264980 110508 265032 110560
rect 170496 110440 170548 110492
rect 214012 110440 214064 110492
rect 247684 110440 247736 110492
rect 265072 110440 265124 110492
rect 231676 110372 231728 110424
rect 262956 110372 263008 110424
rect 282828 110372 282880 110424
rect 295432 110372 295484 110424
rect 231768 110304 231820 110356
rect 244924 110304 244976 110356
rect 177672 109080 177724 109132
rect 214012 109080 214064 109132
rect 167644 109012 167696 109064
rect 213920 109012 213972 109064
rect 260288 109012 260340 109064
rect 265072 109012 265124 109064
rect 354036 109012 354088 109064
rect 397552 109012 397604 109064
rect 442172 109012 442224 109064
rect 443368 109012 443420 109064
rect 167552 108944 167604 108996
rect 170680 108944 170732 108996
rect 231768 108944 231820 108996
rect 242348 108944 242400 108996
rect 282368 108944 282420 108996
rect 305092 108944 305144 108996
rect 389824 108944 389876 108996
rect 397460 108944 397512 108996
rect 442448 108944 442500 108996
rect 443276 108944 443328 108996
rect 231308 108876 231360 108928
rect 235448 108876 235500 108928
rect 378784 108264 378836 108316
rect 397644 108264 397696 108316
rect 203708 107720 203760 107772
rect 213920 107720 213972 107772
rect 170772 107652 170824 107704
rect 214012 107652 214064 107704
rect 253204 107652 253256 107704
rect 264980 107652 265032 107704
rect 231768 107584 231820 107636
rect 264520 107584 264572 107636
rect 282828 107584 282880 107636
rect 291200 107584 291252 107636
rect 231676 107516 231728 107568
rect 263048 107516 263100 107568
rect 298100 106904 298152 106956
rect 367836 106904 367888 106956
rect 185768 106360 185820 106412
rect 213920 106360 213972 106412
rect 377404 106360 377456 106412
rect 397460 106360 397512 106412
rect 166448 106292 166500 106344
rect 214012 106292 214064 106344
rect 262956 106292 263008 106344
rect 265256 106292 265308 106344
rect 370596 106292 370648 106344
rect 397552 106292 397604 106344
rect 231308 106224 231360 106276
rect 240968 106224 241020 106276
rect 294696 106224 294748 106276
rect 397460 106224 397512 106276
rect 442724 106224 442776 106276
rect 452660 106224 452712 106276
rect 231584 106156 231636 106208
rect 234068 106156 234120 106208
rect 173440 105544 173492 105596
rect 202604 105544 202656 105596
rect 236736 105544 236788 105596
rect 246580 105544 246632 105596
rect 374644 105544 374696 105596
rect 397920 105544 397972 105596
rect 231216 105068 231268 105120
rect 231492 105068 231544 105120
rect 202328 104932 202380 104984
rect 213920 104932 213972 104984
rect 263324 104932 263376 104984
rect 265164 104932 265216 104984
rect 178684 104864 178736 104916
rect 214012 104864 214064 104916
rect 245200 104864 245252 104916
rect 264980 104864 265032 104916
rect 442356 104864 442408 104916
rect 445852 104864 445904 104916
rect 231768 104796 231820 104848
rect 247868 104796 247920 104848
rect 281540 104796 281592 104848
rect 284392 104796 284444 104848
rect 347044 104796 347096 104848
rect 397460 104796 397512 104848
rect 391204 104728 391256 104780
rect 397552 104728 397604 104780
rect 231676 104660 231728 104712
rect 236828 104660 236880 104712
rect 167736 104184 167788 104236
rect 185676 104184 185728 104236
rect 171968 104116 172020 104168
rect 195428 104116 195480 104168
rect 263048 104116 263100 104168
rect 265072 104116 265124 104168
rect 238116 103504 238168 103556
rect 264980 103504 265032 103556
rect 230756 103436 230808 103488
rect 249156 103436 249208 103488
rect 359464 103436 359516 103488
rect 397460 103436 397512 103488
rect 231308 102824 231360 102876
rect 235356 102824 235408 102876
rect 256148 102756 256200 102808
rect 263324 102756 263376 102808
rect 325056 102756 325108 102808
rect 366916 102756 366968 102808
rect 198188 102144 198240 102196
rect 213920 102144 213972 102196
rect 249248 102144 249300 102196
rect 264980 102144 265032 102196
rect 449164 102076 449216 102128
rect 583208 102076 583260 102128
rect 231584 102008 231636 102060
rect 257620 102008 257672 102060
rect 230572 101872 230624 101924
rect 232596 101872 232648 101924
rect 442172 101600 442224 101652
rect 445944 101600 445996 101652
rect 363696 101532 363748 101584
rect 439320 101532 439372 101584
rect 329104 101396 329156 101448
rect 360844 101396 360896 101448
rect 176108 100784 176160 100836
rect 214012 100784 214064 100836
rect 262772 100784 262824 100836
rect 265164 100784 265216 100836
rect 169300 100716 169352 100768
rect 213920 100716 213972 100768
rect 255964 100716 256016 100768
rect 264980 100716 265032 100768
rect 392584 100716 392636 100768
rect 397460 100716 397512 100768
rect 231676 100648 231728 100700
rect 258816 100648 258868 100700
rect 442908 100648 442960 100700
rect 449164 100648 449216 100700
rect 231768 100580 231820 100632
rect 245292 100580 245344 100632
rect 164976 99968 165028 100020
rect 196808 99968 196860 100020
rect 202880 99968 202932 100020
rect 217232 99968 217284 100020
rect 282000 99968 282052 100020
rect 309232 99968 309284 100020
rect 165068 99832 165120 99884
rect 171876 99832 171928 99884
rect 371976 99424 372028 99476
rect 408408 99424 408460 99476
rect 172060 99356 172112 99408
rect 213920 99356 213972 99408
rect 254676 99356 254728 99408
rect 264980 99356 265032 99408
rect 336096 99356 336148 99408
rect 405832 99356 405884 99408
rect 231676 99288 231728 99340
rect 250720 99288 250772 99340
rect 377496 99288 377548 99340
rect 429016 99288 429068 99340
rect 231768 99220 231820 99272
rect 239496 99220 239548 99272
rect 398656 99220 398708 99272
rect 403256 99220 403308 99272
rect 405832 99220 405884 99272
rect 580172 99356 580224 99408
rect 436836 99288 436888 99340
rect 439504 99288 439556 99340
rect 434168 99152 434220 99204
rect 445760 99288 445812 99340
rect 246304 98608 246356 98660
rect 264520 98608 264572 98660
rect 205180 98064 205232 98116
rect 213920 98064 213972 98116
rect 189816 97996 189868 98048
rect 214012 97996 214064 98048
rect 261668 97996 261720 98048
rect 264980 97996 265032 98048
rect 356704 97928 356756 97980
rect 432880 97928 432932 97980
rect 438032 97928 438084 97980
rect 447140 97928 447192 97980
rect 392768 97860 392820 97912
rect 403900 97860 403952 97912
rect 167828 97248 167880 97300
rect 202236 97248 202288 97300
rect 213460 97248 213512 97300
rect 264980 97248 265032 97300
rect 432696 97180 432748 97232
rect 440424 97180 440476 97232
rect 413284 96908 413336 96960
rect 416136 96908 416188 96960
rect 409052 96840 409104 96892
rect 409972 96840 410024 96892
rect 423220 96840 423272 96892
rect 429292 96840 429344 96892
rect 210424 96704 210476 96756
rect 196808 96636 196860 96688
rect 213920 96636 213972 96688
rect 231676 96636 231728 96688
rect 246488 96636 246540 96688
rect 382924 96568 382976 96620
rect 420000 96568 420052 96620
rect 412916 96364 412968 96416
rect 413376 96364 413428 96416
rect 219164 96024 219216 96076
rect 230480 96024 230532 96076
rect 232596 96024 232648 96076
rect 213184 95956 213236 96008
rect 225604 95956 225656 96008
rect 178868 95888 178920 95940
rect 214656 95888 214708 95940
rect 227076 95888 227128 95940
rect 262772 95888 262824 95940
rect 432604 95820 432656 95872
rect 439136 95820 439188 95872
rect 401324 95208 401376 95260
rect 402980 95208 403032 95260
rect 413376 95208 413428 95260
rect 582748 95208 582800 95260
rect 259368 95140 259420 95192
rect 279424 95140 279476 95192
rect 353944 95140 353996 95192
rect 429660 95140 429712 95192
rect 267832 95072 267884 95124
rect 269120 95072 269172 95124
rect 366916 95072 366968 95124
rect 412272 95072 412324 95124
rect 216220 94528 216272 94580
rect 232780 94528 232832 94580
rect 66076 94460 66128 94512
rect 111156 94460 111208 94512
rect 176200 94460 176252 94512
rect 202420 94460 202472 94512
rect 216680 94460 216732 94512
rect 223488 94460 223540 94512
rect 226984 94460 227036 94512
rect 247960 94460 248012 94512
rect 120632 93916 120684 93968
rect 176016 93916 176068 93968
rect 100668 93848 100720 93900
rect 166540 93848 166592 93900
rect 421288 93848 421340 93900
rect 582840 93848 582892 93900
rect 267740 93780 267792 93832
rect 273996 93780 274048 93832
rect 322204 93780 322256 93832
rect 426440 93780 426492 93832
rect 381728 93712 381780 93764
rect 424508 93712 424560 93764
rect 67364 93168 67416 93220
rect 97264 93168 97316 93220
rect 124128 93168 124180 93220
rect 166264 93168 166316 93220
rect 216036 93168 216088 93220
rect 243452 93168 243504 93220
rect 262128 93168 262180 93220
rect 270592 93168 270644 93220
rect 64788 93100 64840 93152
rect 98644 93100 98696 93152
rect 118240 93100 118292 93152
rect 180340 93100 180392 93152
rect 220084 93100 220136 93152
rect 265900 93100 265952 93152
rect 108120 92488 108172 92540
rect 122104 92488 122156 92540
rect 258816 92488 258868 92540
rect 260380 92488 260432 92540
rect 125784 92420 125836 92472
rect 173256 92420 173308 92472
rect 217232 92420 217284 92472
rect 280436 92420 280488 92472
rect 373264 92420 373316 92472
rect 432236 92420 432288 92472
rect 110144 92352 110196 92404
rect 112444 92352 112496 92404
rect 133144 92352 133196 92404
rect 169116 92352 169168 92404
rect 171876 91808 171928 91860
rect 187148 91808 187200 91860
rect 213184 91808 213236 91860
rect 236920 91808 236972 91860
rect 60648 91740 60700 91792
rect 100024 91740 100076 91792
rect 178040 91740 178092 91792
rect 213368 91740 213420 91792
rect 398748 91740 398800 91792
rect 583024 91740 583076 91792
rect 103428 91128 103480 91180
rect 108304 91128 108356 91180
rect 85120 91060 85172 91112
rect 105544 91060 105596 91112
rect 111248 91060 111300 91112
rect 115296 91060 115348 91112
rect 116768 91060 116820 91112
rect 132868 91060 132920 91112
rect 115756 90992 115808 91044
rect 174636 90992 174688 91044
rect 223488 90992 223540 91044
rect 280344 90992 280396 91044
rect 243452 90924 243504 90976
rect 281724 90924 281776 90976
rect 185584 90380 185636 90432
rect 213460 90380 213512 90432
rect 218704 90380 218756 90432
rect 239680 90380 239732 90432
rect 67548 90312 67600 90364
rect 115204 90312 115256 90364
rect 193864 90312 193916 90364
rect 223028 90312 223080 90364
rect 119896 89632 119948 89684
rect 171784 89632 171836 89684
rect 360844 89632 360896 89684
rect 430304 89632 430356 89684
rect 151636 89564 151688 89616
rect 167828 89564 167880 89616
rect 168380 89564 168432 89616
rect 206376 89564 206428 89616
rect 224224 89020 224276 89072
rect 242440 89020 242492 89072
rect 64696 88952 64748 89004
rect 111064 88952 111116 89004
rect 192668 88952 192720 89004
rect 216128 88952 216180 89004
rect 221464 88952 221516 89004
rect 250812 88952 250864 89004
rect 122288 88272 122340 88324
rect 196716 88272 196768 88324
rect 276020 88272 276072 88324
rect 443368 88272 443420 88324
rect 109224 88204 109276 88256
rect 170588 88204 170640 88256
rect 216312 88204 216364 88256
rect 280528 88204 280580 88256
rect 366364 88204 366416 88256
rect 425152 88204 425204 88256
rect 178960 87660 179012 87712
rect 214840 87660 214892 87712
rect 75276 87592 75328 87644
rect 112536 87592 112588 87644
rect 204904 87592 204956 87644
rect 253480 87592 253532 87644
rect 88064 86912 88116 86964
rect 172060 86912 172112 86964
rect 246488 86912 246540 86964
rect 305644 86912 305696 86964
rect 432696 86912 432748 86964
rect 114376 86844 114428 86896
rect 192576 86844 192628 86896
rect 225604 86844 225656 86896
rect 281632 86844 281684 86896
rect 195244 86232 195296 86284
rect 222844 86232 222896 86284
rect 299664 86232 299716 86284
rect 444472 86232 444524 86284
rect 3516 85484 3568 85536
rect 17224 85484 17276 85536
rect 108672 85484 108724 85536
rect 188436 85484 188488 85536
rect 214564 85484 214616 85536
rect 413376 85484 413428 85536
rect 151728 85416 151780 85468
rect 171968 85416 172020 85468
rect 177396 84804 177448 84856
rect 243728 84804 243780 84856
rect 97908 84124 97960 84176
rect 177672 84124 177724 84176
rect 126796 84056 126848 84108
rect 164884 84056 164936 84108
rect 207664 83444 207716 83496
rect 220176 83444 220228 83496
rect 222936 83444 222988 83496
rect 238208 83444 238260 83496
rect 324964 83444 325016 83496
rect 440332 83444 440384 83496
rect 86776 82764 86828 82816
rect 189816 82764 189868 82816
rect 294604 82764 294656 82816
rect 432604 82764 432656 82816
rect 153108 82696 153160 82748
rect 178776 82696 178828 82748
rect 217324 82152 217376 82204
rect 239588 82152 239640 82204
rect 67456 82084 67508 82136
rect 123484 82084 123536 82136
rect 206284 82084 206336 82136
rect 258816 82084 258868 82136
rect 343548 82084 343600 82136
rect 404360 82084 404412 82136
rect 113088 81336 113140 81388
rect 184388 81336 184440 81388
rect 135168 81268 135220 81320
rect 160744 81268 160796 81320
rect 214656 80724 214708 80776
rect 247776 80724 247828 80776
rect 195244 80656 195296 80708
rect 235540 80656 235592 80708
rect 304264 80656 304316 80708
rect 360936 80656 360988 80708
rect 111156 79976 111208 80028
rect 176108 79976 176160 80028
rect 331220 79976 331272 80028
rect 331864 79976 331916 80028
rect 436744 79976 436796 80028
rect 107568 79908 107620 79960
rect 169208 79908 169260 79960
rect 214564 79296 214616 79348
rect 254768 79296 254820 79348
rect 101956 78616 102008 78668
rect 173440 78616 173492 78668
rect 108948 77936 109000 77988
rect 238300 77936 238352 77988
rect 125416 77188 125468 77240
rect 176200 77188 176252 77240
rect 122104 77120 122156 77172
rect 164976 77120 165028 77172
rect 332600 76508 332652 76560
rect 393412 76508 393464 76560
rect 98644 75828 98696 75880
rect 214748 75828 214800 75880
rect 244924 75828 244976 75880
rect 247040 75828 247092 75880
rect 439228 75828 439280 75880
rect 115296 75760 115348 75812
rect 177580 75760 177632 75812
rect 67640 74468 67692 74520
rect 174728 74468 174780 74520
rect 100668 74400 100720 74452
rect 170496 74400 170548 74452
rect 335360 73788 335412 73840
rect 441712 73788 441764 73840
rect 107568 72496 107620 72548
rect 229744 72496 229796 72548
rect 122748 72428 122800 72480
rect 261576 72428 261628 72480
rect 344284 72428 344336 72480
rect 414204 72428 414256 72480
rect 100024 71680 100076 71732
rect 202328 71680 202380 71732
rect 126888 71612 126940 71664
rect 173164 71612 173216 71664
rect 99196 70320 99248 70372
rect 171876 70320 171928 70372
rect 48136 69640 48188 69692
rect 249248 69640 249300 69692
rect 336740 69640 336792 69692
rect 440240 69640 440292 69692
rect 115204 68960 115256 69012
rect 196808 68960 196860 69012
rect 106096 68892 106148 68944
rect 180248 68892 180300 68944
rect 330484 67668 330536 67720
rect 335360 67668 335412 67720
rect 334624 67600 334676 67652
rect 336740 67600 336792 67652
rect 103336 67532 103388 67584
rect 199384 67532 199436 67584
rect 337476 67532 337528 67584
rect 401968 67532 402020 67584
rect 124036 67464 124088 67516
rect 178868 67464 178920 67516
rect 323676 66852 323728 66904
rect 337476 66852 337528 66904
rect 110144 66172 110196 66224
rect 192668 66172 192720 66224
rect 151544 66104 151596 66156
rect 169024 66104 169076 66156
rect 292488 65492 292540 65544
rect 428372 65492 428424 65544
rect 102048 64812 102100 64864
rect 205088 64812 205140 64864
rect 112536 64744 112588 64796
rect 178960 64744 179012 64796
rect 284944 64132 284996 64184
rect 352748 64132 352800 64184
rect 89628 63452 89680 63504
rect 162124 63452 162176 63504
rect 292672 63452 292724 63504
rect 425704 63452 425756 63504
rect 124128 63384 124180 63436
rect 193956 63384 194008 63436
rect 266360 62772 266412 62824
rect 292672 62772 292724 62824
rect 104164 62024 104216 62076
rect 203524 62024 203576 62076
rect 262956 61412 263008 61464
rect 399484 61412 399536 61464
rect 59268 61344 59320 61396
rect 263048 61344 263100 61396
rect 116584 60664 116636 60716
rect 210516 60664 210568 60716
rect 84108 59984 84160 60036
rect 242256 59984 242308 60036
rect 3056 59304 3108 59356
rect 40684 59304 40736 59356
rect 108304 59304 108356 59356
rect 209136 59304 209188 59356
rect 311900 59304 311952 59356
rect 407120 59304 407172 59356
rect 115848 58624 115900 58676
rect 247684 58624 247736 58676
rect 248328 58624 248380 58676
rect 311900 58624 311952 58676
rect 107476 57876 107528 57928
rect 211804 57876 211856 57928
rect 220176 57264 220228 57316
rect 259460 57264 259512 57316
rect 342996 57264 343048 57316
rect 104808 57196 104860 57248
rect 260288 57196 260340 57248
rect 346400 57196 346452 57248
rect 446036 57196 446088 57248
rect 123484 56516 123536 56568
rect 213276 56516 213328 56568
rect 91008 55836 91060 55888
rect 264428 55836 264480 55888
rect 112444 55156 112496 55208
rect 198096 55156 198148 55208
rect 382924 54544 382976 54596
rect 422576 54544 422628 54596
rect 89628 54476 89680 54528
rect 243544 54476 243596 54528
rect 335360 54476 335412 54528
rect 383016 54476 383068 54528
rect 340788 53728 340840 53780
rect 435456 53728 435508 53780
rect 340144 53252 340196 53304
rect 340788 53252 340840 53304
rect 146944 53116 146996 53168
rect 227076 53116 227128 53168
rect 41328 53048 41380 53100
rect 231124 53048 231176 53100
rect 117136 52368 117188 52420
rect 191196 52368 191248 52420
rect 250536 51756 250588 51808
rect 416780 51756 416832 51808
rect 17868 51688 17920 51740
rect 254676 51688 254728 51740
rect 106188 51008 106240 51060
rect 195336 51008 195388 51060
rect 136548 50940 136600 50992
rect 180156 50940 180208 50992
rect 52368 50328 52420 50380
rect 135260 50328 135312 50380
rect 186964 50328 187016 50380
rect 302976 50328 303028 50380
rect 321560 50328 321612 50380
rect 408500 50328 408552 50380
rect 86868 49648 86920 49700
rect 205180 49648 205232 49700
rect 114468 48968 114520 49020
rect 236644 48968 236696 49020
rect 297364 48968 297416 49020
rect 444380 48968 444432 49020
rect 129648 48220 129700 48272
rect 192484 48220 192536 48272
rect 227076 47608 227128 47660
rect 269120 47608 269172 47660
rect 133144 47540 133196 47592
rect 217324 47540 217376 47592
rect 268384 47540 268436 47592
rect 454132 47540 454184 47592
rect 300768 46860 300820 46912
rect 400680 46860 400732 46912
rect 85488 46248 85540 46300
rect 267004 46248 267056 46300
rect 71044 46180 71096 46232
rect 258724 46180 258776 46232
rect 269764 46180 269816 46232
rect 299480 46180 299532 46232
rect 300768 46180 300820 46232
rect 3516 45500 3568 45552
rect 43444 45500 43496 45552
rect 95056 44820 95108 44872
rect 253204 44820 253256 44872
rect 257344 44820 257396 44872
rect 400864 44820 400916 44872
rect 12256 43392 12308 43444
rect 245016 43392 245068 43444
rect 246396 43392 246448 43444
rect 405740 43392 405792 43444
rect 283564 42712 283616 42764
rect 452752 42712 452804 42764
rect 37188 42100 37240 42152
rect 147036 42100 147088 42152
rect 147128 42100 147180 42152
rect 230480 42100 230532 42152
rect 105544 42032 105596 42084
rect 250444 42032 250496 42084
rect 99288 40740 99340 40792
rect 239404 40740 239456 40792
rect 46848 40672 46900 40724
rect 240876 40672 240928 40724
rect 228364 39312 228416 39364
rect 258080 39312 258132 39364
rect 436100 39312 436152 39364
rect 39948 37884 40000 37936
rect 222936 37884 222988 37936
rect 314660 37884 314712 37936
rect 456892 37884 456944 37936
rect 320824 37204 320876 37256
rect 392584 37204 392636 37256
rect 320180 36864 320232 36916
rect 320824 36864 320876 36916
rect 247040 36660 247092 36712
rect 248328 36660 248380 36712
rect 54484 36524 54536 36576
rect 265716 36524 265768 36576
rect 316776 35844 316828 35896
rect 443000 35844 443052 35896
rect 186964 35232 187016 35284
rect 221464 35232 221516 35284
rect 61936 35164 61988 35216
rect 224316 35164 224368 35216
rect 316040 34484 316092 34536
rect 316776 34484 316828 34536
rect 86868 33804 86920 33856
rect 226984 33804 227036 33856
rect 61384 33736 61436 33788
rect 279424 33736 279476 33788
rect 3516 33056 3568 33108
rect 15844 33056 15896 33108
rect 74448 32444 74500 32496
rect 260104 32444 260156 32496
rect 62028 32376 62080 32428
rect 274640 32376 274692 32428
rect 309876 32376 309928 32428
rect 393964 32376 394016 32428
rect 78588 31084 78640 31136
rect 262864 31084 262916 31136
rect 60004 31016 60056 31068
rect 246304 31016 246356 31068
rect 252560 31016 252612 31068
rect 304264 31016 304316 31068
rect 112444 29656 112496 29708
rect 204904 29656 204956 29708
rect 56508 29588 56560 29640
rect 264336 29588 264388 29640
rect 282276 29588 282328 29640
rect 389916 29588 389968 29640
rect 160744 28364 160796 28416
rect 214656 28364 214708 28416
rect 37096 28296 37148 28348
rect 178684 28296 178736 28348
rect 112 28228 164 28280
rect 147128 28228 147180 28280
rect 188344 28228 188396 28280
rect 270500 28228 270552 28280
rect 277400 28228 277452 28280
rect 294604 28228 294656 28280
rect 303620 28228 303672 28280
rect 327080 28228 327132 28280
rect 274640 27548 274692 27600
rect 417424 27548 417476 27600
rect 81348 26936 81400 26988
rect 232504 26936 232556 26988
rect 16488 26868 16540 26920
rect 185584 26868 185636 26920
rect 270500 26188 270552 26240
rect 371884 26188 371936 26240
rect 200764 25576 200816 25628
rect 268476 25576 268528 25628
rect 125508 25508 125560 25560
rect 216036 25508 216088 25560
rect 327080 24148 327132 24200
rect 419356 24148 419408 24200
rect 100668 24080 100720 24132
rect 235264 24080 235316 24132
rect 264336 24080 264388 24132
rect 374736 24080 374788 24132
rect 67180 22788 67232 22840
rect 255964 22788 256016 22840
rect 259552 22788 259604 22840
rect 395344 22788 395396 22840
rect 20628 22720 20680 22772
rect 261484 22720 261536 22772
rect 111616 21428 111668 21480
rect 238024 21428 238076 21480
rect 57888 21360 57940 21412
rect 251916 21360 251968 21412
rect 257436 21360 257488 21412
rect 447232 21360 447284 21412
rect 334716 20612 334768 20664
rect 335268 20612 335320 20664
rect 429292 20612 429344 20664
rect 45468 20000 45520 20052
rect 133144 20000 133196 20052
rect 189724 20000 189776 20052
rect 215944 20000 215996 20052
rect 88248 19932 88300 19984
rect 249064 19932 249116 19984
rect 250444 19932 250496 19984
rect 385040 19932 385092 19984
rect 323584 19320 323636 19372
rect 327080 19320 327132 19372
rect 222844 18640 222896 18692
rect 245660 18640 245712 18692
rect 103428 18572 103480 18624
rect 236736 18572 236788 18624
rect 409972 18572 410024 18624
rect 50988 17892 51040 17944
rect 296720 17892 296772 17944
rect 297364 17892 297416 17944
rect 28816 17212 28868 17264
rect 242164 17212 242216 17264
rect 243544 17212 243596 17264
rect 413284 17212 413336 17264
rect 249156 16532 249208 16584
rect 370596 16532 370648 16584
rect 126244 15920 126296 15972
rect 214564 15920 214616 15972
rect 9588 15852 9640 15904
rect 198004 15852 198056 15904
rect 341524 15852 341576 15904
rect 342352 15852 342404 15904
rect 407764 15852 407816 15904
rect 248420 15172 248472 15224
rect 249156 15172 249208 15224
rect 255872 15104 255924 15156
rect 311164 15104 311216 15156
rect 96252 14424 96304 14476
rect 218704 14424 218756 14476
rect 196624 13744 196676 13796
rect 264336 13744 264388 13796
rect 280896 13744 280948 13796
rect 367744 13744 367796 13796
rect 112812 13132 112864 13184
rect 160744 13132 160796 13184
rect 45284 13064 45336 13116
rect 224224 13064 224276 13116
rect 288348 13064 288400 13116
rect 414664 13064 414716 13116
rect 280712 12452 280764 12504
rect 280896 12452 280948 12504
rect 348056 12384 348108 12436
rect 448520 12384 448572 12436
rect 268476 12316 268528 12368
rect 349804 12316 349856 12368
rect 267740 11908 267792 11960
rect 268476 11908 268528 11960
rect 135260 11772 135312 11824
rect 136456 11772 136508 11824
rect 106832 11704 106884 11756
rect 227076 11704 227128 11756
rect 242164 11704 242216 11756
rect 264244 11704 264296 11756
rect 71504 10344 71556 10396
rect 195244 10344 195296 10396
rect 311440 10344 311492 10396
rect 378784 10344 378836 10396
rect 54944 10276 54996 10328
rect 238116 10276 238168 10328
rect 261760 10276 261812 10328
rect 449900 10276 449952 10328
rect 180432 9596 180484 9648
rect 242900 9596 242952 9648
rect 243544 9596 243596 9648
rect 257344 9596 257396 9648
rect 258724 9596 258776 9648
rect 334624 9596 334676 9648
rect 337476 9596 337528 9648
rect 349988 9596 350040 9648
rect 350448 9596 350500 9648
rect 439412 9596 439464 9648
rect 91560 8984 91612 9036
rect 202236 8984 202288 9036
rect 332692 8984 332744 9036
rect 349988 8984 350040 9036
rect 26516 8916 26568 8968
rect 146944 8916 146996 8968
rect 328000 8916 328052 8968
rect 358820 8916 358872 8968
rect 59636 7624 59688 7676
rect 112444 7624 112496 7676
rect 117596 7624 117648 7676
rect 206284 7624 206336 7676
rect 329196 7624 329248 7676
rect 381636 7624 381688 7676
rect 66720 7556 66772 7608
rect 240784 7556 240836 7608
rect 288992 7556 289044 7608
rect 354036 7556 354088 7608
rect 308404 6808 308456 6860
rect 309784 6808 309836 6860
rect 325056 6808 325108 6860
rect 411628 6808 411680 6860
rect 24216 6196 24268 6248
rect 191104 6196 191156 6248
rect 62028 6128 62080 6180
rect 233884 6128 233936 6180
rect 278044 6128 278096 6180
rect 285404 6128 285456 6180
rect 427912 6128 427964 6180
rect 282828 5516 282880 5568
rect 283564 5516 283616 5568
rect 324504 5516 324556 5568
rect 325056 5516 325108 5568
rect 306748 5448 306800 5500
rect 307024 5448 307076 5500
rect 396724 5448 396776 5500
rect 105728 4768 105780 4820
rect 186964 4768 187016 4820
rect 232596 4156 232648 4208
rect 235816 4156 235868 4208
rect 247776 4088 247828 4140
rect 250536 4088 250588 4140
rect 265348 4088 265400 4140
rect 269764 4088 269816 4140
rect 279424 4088 279476 4140
rect 286324 4088 286376 4140
rect 305552 4088 305604 4140
rect 307116 4088 307168 4140
rect 315304 4088 315356 4140
rect 319720 4088 319772 4140
rect 326344 4088 326396 4140
rect 326804 4088 326856 4140
rect 329104 4088 329156 4140
rect 268384 4020 268436 4072
rect 268844 4020 268896 4072
rect 302884 4020 302936 4072
rect 309876 4020 309928 4072
rect 345756 4020 345808 4072
rect 402980 4020 403032 4072
rect 254676 3748 254728 3800
rect 258080 3748 258132 3800
rect 351184 3612 351236 3664
rect 351644 3612 351696 3664
rect 11152 3544 11204 3596
rect 12256 3544 12308 3596
rect 20536 3544 20588 3596
rect 2872 3476 2924 3528
rect 4068 3476 4120 3528
rect 8760 3476 8812 3528
rect 9588 3476 9640 3528
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 15936 3476 15988 3528
rect 16488 3476 16540 3528
rect 17040 3476 17092 3528
rect 17868 3476 17920 3528
rect 18236 3476 18288 3528
rect 19248 3476 19300 3528
rect 19432 3476 19484 3528
rect 20628 3476 20680 3528
rect 25320 3544 25372 3596
rect 26148 3544 26200 3596
rect 27712 3544 27764 3596
rect 28816 3544 28868 3596
rect 32404 3544 32456 3596
rect 33048 3544 33100 3596
rect 33600 3544 33652 3596
rect 34428 3544 34480 3596
rect 34796 3544 34848 3596
rect 35808 3544 35860 3596
rect 35992 3544 36044 3596
rect 37096 3544 37148 3596
rect 40684 3544 40736 3596
rect 41328 3544 41380 3596
rect 41880 3544 41932 3596
rect 42708 3544 42760 3596
rect 43076 3544 43128 3596
rect 44088 3544 44140 3596
rect 44272 3544 44324 3596
rect 45376 3544 45428 3596
rect 54484 3544 54536 3596
rect 64328 3544 64380 3596
rect 64788 3544 64840 3596
rect 48964 3476 49016 3528
rect 49608 3476 49660 3528
rect 50160 3476 50212 3528
rect 50896 3476 50948 3528
rect 52552 3476 52604 3528
rect 53656 3476 53708 3528
rect 56048 3476 56100 3528
rect 56508 3476 56560 3528
rect 57244 3476 57296 3528
rect 57796 3476 57848 3528
rect 58440 3476 58492 3528
rect 59268 3476 59320 3528
rect 60832 3476 60884 3528
rect 61936 3476 61988 3528
rect 63224 3476 63276 3528
rect 71044 3544 71096 3596
rect 78496 3544 78548 3596
rect 65524 3476 65576 3528
rect 66168 3476 66220 3528
rect 67916 3476 67968 3528
rect 68928 3476 68980 3528
rect 69112 3476 69164 3528
rect 70216 3476 70268 3528
rect 72608 3476 72660 3528
rect 73068 3476 73120 3528
rect 73804 3476 73856 3528
rect 74448 3476 74500 3528
rect 75000 3476 75052 3528
rect 75828 3476 75880 3528
rect 76196 3476 76248 3528
rect 77208 3476 77260 3528
rect 77392 3476 77444 3528
rect 78588 3476 78640 3528
rect 80888 3544 80940 3596
rect 81348 3544 81400 3596
rect 83280 3544 83332 3596
rect 84108 3544 84160 3596
rect 87604 3544 87656 3596
rect 84476 3476 84528 3528
rect 85488 3476 85540 3528
rect 89168 3476 89220 3528
rect 89628 3476 89680 3528
rect 90364 3476 90416 3528
rect 91008 3476 91060 3528
rect 92756 3476 92808 3528
rect 93768 3476 93820 3528
rect 93952 3476 94004 3528
rect 95056 3476 95108 3528
rect 97448 3476 97500 3528
rect 97908 3476 97960 3528
rect 98644 3476 98696 3528
rect 99288 3476 99340 3528
rect 99840 3476 99892 3528
rect 100668 3476 100720 3528
rect 101036 3476 101088 3528
rect 102048 3476 102100 3528
rect 106924 3476 106976 3528
rect 107568 3476 107620 3528
rect 108120 3476 108172 3528
rect 108948 3476 109000 3528
rect 109316 3476 109368 3528
rect 126244 3544 126296 3596
rect 124680 3476 124732 3528
rect 125508 3476 125560 3528
rect 125876 3476 125928 3528
rect 126888 3476 126940 3528
rect 129372 3476 129424 3528
rect 130384 3476 130436 3528
rect 140044 3476 140096 3528
rect 141424 3476 141476 3528
rect 143540 3476 143592 3528
rect 144828 3476 144880 3528
rect 251180 3476 251232 3528
rect 251916 3476 251968 3528
rect 258264 3476 258316 3528
rect 258724 3476 258776 3528
rect 272432 3476 272484 3528
rect 273260 3476 273312 3528
rect 273628 3476 273680 3528
rect 274548 3476 274600 3528
rect 292488 3476 292540 3528
rect 294880 3476 294932 3528
rect 296720 3476 296772 3528
rect 297272 3476 297324 3528
rect 307944 3476 307996 3528
rect 309140 3476 309192 3528
rect 313832 3476 313884 3528
rect 314568 3476 314620 3528
rect 316040 3476 316092 3528
rect 317328 3476 317380 3528
rect 324412 3476 324464 3528
rect 325608 3476 325660 3528
rect 332600 3476 332652 3528
rect 333888 3476 333940 3528
rect 339868 3476 339920 3528
rect 340788 3476 340840 3528
rect 340972 3476 341024 3528
rect 342352 3476 342404 3528
rect 582196 3476 582248 3528
rect 583576 3476 583628 3528
rect 106832 3408 106884 3460
rect 114008 3408 114060 3460
rect 114468 3408 114520 3460
rect 115204 3408 115256 3460
rect 115848 3408 115900 3460
rect 116400 3408 116452 3460
rect 117228 3408 117280 3460
rect 122288 3408 122340 3460
rect 122748 3408 122800 3460
rect 123484 3408 123536 3460
rect 220084 3408 220136 3460
rect 245660 3408 245712 3460
rect 257068 3408 257120 3460
rect 276112 3408 276164 3460
rect 277124 3408 277176 3460
rect 282184 3408 282236 3460
rect 312636 3408 312688 3460
rect 323676 3408 323728 3460
rect 349252 3408 349304 3460
rect 360844 3408 360896 3460
rect 4068 3340 4120 3392
rect 240508 3340 240560 3392
rect 246396 3340 246448 3392
rect 241704 3272 241756 3324
rect 244924 3272 244976 3324
rect 110512 3068 110564 3120
rect 111524 3068 111576 3120
rect 581000 3068 581052 3120
rect 583760 3068 583812 3120
rect 245200 2932 245252 2984
rect 247040 2932 247092 2984
rect 271788 2728 271840 2780
rect 445852 2728 445904 2780
rect 51356 2116 51408 2168
rect 60004 2116 60056 2168
rect 102232 2116 102284 2168
rect 213184 2116 213236 2168
rect 239312 2116 239364 2168
rect 270592 2116 270644 2168
rect 271788 2116 271840 2168
rect 7656 2048 7708 2100
rect 105544 2048 105596 2100
rect 118792 2048 118844 2100
rect 242164 2048 242216 2100
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 702506 8156 703520
rect 24320 702642 24348 703520
rect 24308 702636 24360 702642
rect 24308 702578 24360 702584
rect 8116 702500 8168 702506
rect 8116 702442 8168 702448
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 2778 658200 2834 658209
rect 2778 658135 2834 658144
rect 2792 657014 2820 658135
rect 2780 657008 2832 657014
rect 2780 656950 2832 656956
rect 3056 580780 3108 580786
rect 3056 580722 3108 580728
rect 3068 580009 3096 580722
rect 3054 580000 3110 580009
rect 3054 579935 3110 579944
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 2778 553888 2834 553897
rect 2778 553823 2780 553832
rect 2832 553823 2834 553832
rect 2780 553794 2832 553800
rect 3436 543046 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 14464 670744 14516 670750
rect 14464 670686 14516 670692
rect 4804 657008 4856 657014
rect 4804 656950 4856 656956
rect 3516 632120 3568 632126
rect 3514 632088 3516 632097
rect 3568 632088 3570 632097
rect 3514 632023 3570 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 4816 591326 4844 656950
rect 4804 591320 4856 591326
rect 4804 591262 4856 591268
rect 7564 589348 7616 589354
rect 7564 589290 7616 589296
rect 7576 580786 7604 589290
rect 7564 580780 7616 580786
rect 7564 580722 7616 580728
rect 4804 553852 4856 553858
rect 4804 553794 4856 553800
rect 3424 543040 3476 543046
rect 3424 542982 3476 542988
rect 4816 540258 4844 553794
rect 14476 541686 14504 670686
rect 21364 632120 21416 632126
rect 21364 632062 21416 632068
rect 21376 576162 21404 632062
rect 22744 618316 22796 618322
rect 22744 618258 22796 618264
rect 21364 576156 21416 576162
rect 21364 576098 21416 576104
rect 14464 541680 14516 541686
rect 14464 541622 14516 541628
rect 4804 540252 4856 540258
rect 4804 540194 4856 540200
rect 7564 538892 7616 538898
rect 7564 538834 7616 538840
rect 4802 534712 4858 534721
rect 4802 534647 4858 534656
rect 3424 532024 3476 532030
rect 3424 531966 3476 531972
rect 3436 527921 3464 531966
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 2780 501900 2832 501906
rect 2780 501842 2832 501848
rect 2792 501809 2820 501842
rect 2778 501800 2834 501809
rect 2778 501735 2834 501744
rect 2778 462632 2834 462641
rect 2778 462567 2780 462576
rect 2832 462567 2834 462576
rect 2780 462538 2832 462544
rect 3436 451926 3464 527847
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 4816 501906 4844 534647
rect 4804 501900 4856 501906
rect 4804 501842 4856 501848
rect 3514 475688 3570 475697
rect 3514 475623 3570 475632
rect 3528 474026 3556 475623
rect 7576 474026 7604 538834
rect 12348 537600 12400 537606
rect 12348 537542 12400 537548
rect 3516 474020 3568 474026
rect 3516 473962 3568 473968
rect 7564 474020 7616 474026
rect 7564 473962 7616 473968
rect 4804 462596 4856 462602
rect 4804 462538 4856 462544
rect 3424 451920 3476 451926
rect 3424 451862 3476 451868
rect 4816 450566 4844 462538
rect 4804 450560 4856 450566
rect 4804 450502 4856 450508
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 12360 447166 12388 537542
rect 22756 536081 22784 618258
rect 40052 594114 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 62028 703044 62080 703050
rect 62028 702986 62080 702992
rect 40040 594108 40092 594114
rect 40040 594050 40092 594056
rect 55128 587920 55180 587926
rect 55128 587862 55180 587868
rect 50896 582412 50948 582418
rect 50896 582354 50948 582360
rect 39948 576156 40000 576162
rect 39948 576098 40000 576104
rect 39960 575550 39988 576098
rect 39948 575544 40000 575550
rect 39948 575486 40000 575492
rect 37188 561740 37240 561746
rect 37188 561682 37240 561688
rect 34520 543040 34572 543046
rect 34520 542982 34572 542988
rect 34532 542434 34560 542982
rect 34520 542428 34572 542434
rect 34520 542370 34572 542376
rect 35808 542428 35860 542434
rect 35808 542370 35860 542376
rect 22742 536072 22798 536081
rect 22742 536007 22798 536016
rect 34428 523728 34480 523734
rect 34428 523670 34480 523676
rect 14464 514820 14516 514826
rect 14464 514762 14516 514768
rect 14476 455394 14504 514762
rect 15844 474020 15896 474026
rect 15844 473962 15896 473968
rect 14464 455388 14516 455394
rect 14464 455330 14516 455336
rect 11704 447160 11756 447166
rect 11704 447102 11756 447108
rect 12348 447160 12400 447166
rect 12348 447102 12400 447108
rect 7564 445800 7616 445806
rect 7564 445742 7616 445748
rect 3424 423632 3476 423638
rect 3422 423600 3424 423609
rect 3476 423600 3478 423609
rect 3422 423535 3478 423544
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3436 389201 3464 410479
rect 7576 397594 7604 445742
rect 11716 423638 11744 447102
rect 14464 428460 14516 428466
rect 14464 428402 14516 428408
rect 11704 423632 11756 423638
rect 11704 423574 11756 423580
rect 3516 397588 3568 397594
rect 3516 397530 3568 397536
rect 7564 397588 7616 397594
rect 7564 397530 7616 397536
rect 3528 397497 3556 397530
rect 3514 397488 3570 397497
rect 3514 397423 3570 397432
rect 3422 389192 3478 389201
rect 3422 389127 3478 389136
rect 7564 386436 7616 386442
rect 7564 386378 7616 386384
rect 4802 385656 4858 385665
rect 4802 385591 4858 385600
rect 3608 381540 3660 381546
rect 3608 381482 3660 381488
rect 2964 371408 3016 371414
rect 2962 371376 2964 371385
rect 3016 371376 3018 371385
rect 2962 371311 3018 371320
rect 3424 358624 3476 358630
rect 3424 358566 3476 358572
rect 3436 358465 3464 358566
rect 3422 358456 3478 358465
rect 3422 358391 3478 358400
rect 3424 355428 3476 355434
rect 3424 355370 3476 355376
rect 20 328500 72 328506
rect 20 328442 72 328448
rect 32 6769 60 328442
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3146 267200 3202 267209
rect 3146 267135 3202 267144
rect 3160 267034 3188 267135
rect 3148 267028 3200 267034
rect 3148 266970 3200 266976
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3160 253978 3188 254079
rect 3148 253972 3200 253978
rect 3148 253914 3200 253920
rect 3332 241120 3384 241126
rect 3330 241088 3332 241097
rect 3384 241088 3386 241097
rect 3330 241023 3386 241032
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 2780 188896 2832 188902
rect 2778 188864 2780 188873
rect 2832 188864 2834 188873
rect 2778 188799 2834 188808
rect 3332 164212 3384 164218
rect 3332 164154 3384 164160
rect 3344 162897 3372 164154
rect 3330 162888 3386 162897
rect 3330 162823 3386 162832
rect 3332 137964 3384 137970
rect 3332 137906 3384 137912
rect 3344 136785 3372 137906
rect 3330 136776 3386 136785
rect 3330 136711 3386 136720
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 112 28280 164 28286
rect 112 28222 164 28228
rect 18 6760 74 6769
rect 18 6695 74 6704
rect 124 490 152 28222
rect 3436 19417 3464 355370
rect 3514 353968 3570 353977
rect 3514 353903 3570 353912
rect 3528 97617 3556 353903
rect 3620 345409 3648 381482
rect 4816 371414 4844 385591
rect 4804 371408 4856 371414
rect 4804 371350 4856 371356
rect 3606 345400 3662 345409
rect 3606 345335 3662 345344
rect 4816 321570 4844 371350
rect 7576 358630 7604 386378
rect 11704 377460 11756 377466
rect 11704 377402 11756 377408
rect 7564 358624 7616 358630
rect 7564 358566 7616 358572
rect 7562 329896 7618 329905
rect 7562 329831 7618 329840
rect 4804 321564 4856 321570
rect 4804 321506 4856 321512
rect 4068 319456 4120 319462
rect 4068 319398 4120 319404
rect 4080 319297 4108 319398
rect 4066 319288 4122 319297
rect 4066 319223 4122 319232
rect 3606 293176 3662 293185
rect 3606 293111 3662 293120
rect 3620 292602 3648 293111
rect 3608 292596 3660 292602
rect 3608 292538 3660 292544
rect 4080 269822 4108 319223
rect 4804 316736 4856 316742
rect 4804 316678 4856 316684
rect 4068 269816 4120 269822
rect 4068 269758 4120 269764
rect 4816 188902 4844 316678
rect 7576 241126 7604 329831
rect 11716 319462 11744 377402
rect 11704 319456 11756 319462
rect 11704 319398 11756 319404
rect 11704 311160 11756 311166
rect 11704 311102 11756 311108
rect 11716 253978 11744 311102
rect 14476 269074 14504 428402
rect 15856 388482 15884 473962
rect 25504 448588 25556 448594
rect 25504 448530 25556 448536
rect 15844 388476 15896 388482
rect 15844 388418 15896 388424
rect 25516 369850 25544 448530
rect 25504 369844 25556 369850
rect 25504 369786 25556 369792
rect 26148 369844 26200 369850
rect 26148 369786 26200 369792
rect 21362 335472 21418 335481
rect 21362 335407 21418 335416
rect 18604 292596 18656 292602
rect 18604 292538 18656 292544
rect 17868 280220 17920 280226
rect 17868 280162 17920 280168
rect 12440 269068 12492 269074
rect 12440 269010 12492 269016
rect 14464 269068 14516 269074
rect 14464 269010 14516 269016
rect 12452 267034 12480 269010
rect 12440 267028 12492 267034
rect 12440 266970 12492 266976
rect 12452 266422 12480 266970
rect 12440 266416 12492 266422
rect 12440 266358 12492 266364
rect 13084 266416 13136 266422
rect 13084 266358 13136 266364
rect 10968 253972 11020 253978
rect 10968 253914 11020 253920
rect 11704 253972 11756 253978
rect 11704 253914 11756 253920
rect 7564 241120 7616 241126
rect 7564 241062 7616 241068
rect 10980 227089 11008 253914
rect 13096 238746 13124 266358
rect 13084 238740 13136 238746
rect 13084 238682 13136 238688
rect 11702 229120 11758 229129
rect 11702 229055 11758 229064
rect 10966 227080 11022 227089
rect 10966 227015 11022 227024
rect 4804 188896 4856 188902
rect 4804 188838 4856 188844
rect 11716 150414 11744 229055
rect 15842 213208 15898 213217
rect 15842 213143 15898 213152
rect 3608 150408 3660 150414
rect 3608 150350 3660 150356
rect 11704 150408 11756 150414
rect 11704 150350 11756 150356
rect 3620 149841 3648 150350
rect 3606 149832 3662 149841
rect 3606 149767 3662 149776
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 12346 80744 12402 80753
rect 12346 80679 12402 80688
rect 5446 79520 5502 79529
rect 5446 79455 5502 79464
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 4066 36544 4122 36553
rect 4066 36479 4122 36488
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 1674 4856 1730 4865
rect 1674 4791 1730 4800
rect 400 598 612 626
rect 400 490 428 598
rect 124 462 428 490
rect 584 480 612 598
rect 1688 480 1716 4791
rect 4080 3534 4108 36479
rect 5460 6914 5488 79455
rect 10966 55856 11022 55865
rect 10966 55791 11022 55800
rect 6826 39264 6882 39273
rect 6826 39199 6882 39208
rect 6840 6914 6868 39199
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 5276 6886 5488 6914
rect 6472 6886 6868 6914
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 2884 480 2912 3470
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 4080 480 4108 3334
rect 5276 480 5304 6886
rect 6472 480 6500 6886
rect 9600 3534 9628 15846
rect 10980 3534 11008 55791
rect 12256 43444 12308 43450
rect 12256 43386 12308 43392
rect 12268 16574 12296 43386
rect 12176 16546 12296 16574
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 7668 480 7696 2042
rect 8772 480 8800 3470
rect 9968 480 9996 3470
rect 11164 480 11192 3538
rect 12176 3482 12204 16546
rect 12360 6914 12388 80679
rect 13726 77888 13782 77897
rect 13726 77823 13782 77832
rect 13740 6914 13768 77823
rect 15106 76528 15162 76537
rect 15106 76463 15162 76472
rect 15120 6914 15148 76463
rect 15856 33114 15884 213143
rect 17880 190369 17908 280162
rect 18616 241505 18644 292538
rect 18602 241496 18658 241505
rect 18602 241431 18658 241440
rect 17866 190360 17922 190369
rect 17866 190295 17922 190304
rect 17880 189145 17908 190295
rect 17222 189136 17278 189145
rect 17222 189071 17278 189080
rect 17866 189136 17922 189145
rect 17866 189071 17922 189080
rect 17236 85542 17264 189071
rect 21376 137970 21404 335407
rect 26160 293962 26188 369786
rect 33784 330540 33836 330546
rect 33784 330482 33836 330488
rect 33796 306338 33824 330482
rect 33784 306332 33836 306338
rect 33784 306274 33836 306280
rect 30288 295384 30340 295390
rect 30288 295326 30340 295332
rect 26148 293956 26200 293962
rect 26148 293898 26200 293904
rect 30300 191729 30328 295326
rect 32404 269816 32456 269822
rect 32404 269758 32456 269764
rect 32416 261526 32444 269758
rect 32404 261520 32456 261526
rect 32404 261462 32456 261468
rect 34440 258058 34468 523670
rect 35820 396778 35848 542370
rect 37200 429146 37228 561682
rect 39960 449886 39988 575486
rect 48136 569220 48188 569226
rect 48136 569162 48188 569168
rect 43444 565888 43496 565894
rect 43444 565830 43496 565836
rect 41328 560312 41380 560318
rect 41328 560254 41380 560260
rect 41340 534070 41368 560254
rect 43456 536790 43484 565830
rect 43996 554804 44048 554810
rect 43996 554746 44048 554752
rect 43444 536784 43496 536790
rect 43444 536726 43496 536732
rect 41328 534064 41380 534070
rect 41328 534006 41380 534012
rect 39948 449880 40000 449886
rect 39948 449822 40000 449828
rect 39946 445768 40002 445777
rect 39946 445703 40002 445712
rect 36728 429140 36780 429146
rect 36728 429082 36780 429088
rect 37188 429140 37240 429146
rect 37188 429082 37240 429088
rect 36740 428466 36768 429082
rect 36728 428460 36780 428466
rect 36728 428402 36780 428408
rect 35808 396772 35860 396778
rect 35808 396714 35860 396720
rect 39302 330032 39358 330041
rect 39302 329967 39358 329976
rect 35164 309800 35216 309806
rect 35164 309742 35216 309748
rect 34428 258052 34480 258058
rect 34428 257994 34480 258000
rect 29642 191720 29698 191729
rect 29642 191655 29698 191664
rect 30286 191720 30342 191729
rect 30286 191655 30342 191664
rect 29656 190505 29684 191655
rect 29642 190496 29698 190505
rect 29642 190431 29698 190440
rect 29656 164218 29684 190431
rect 32404 188352 32456 188358
rect 32404 188294 32456 188300
rect 29644 164212 29696 164218
rect 29644 164154 29696 164160
rect 21364 137964 21416 137970
rect 21364 137906 21416 137912
rect 32416 111790 32444 188294
rect 32404 111784 32456 111790
rect 32404 111726 32456 111732
rect 17224 85536 17276 85542
rect 17224 85478 17276 85484
rect 34426 83464 34482 83473
rect 34426 83399 34482 83408
rect 26146 79384 26202 79393
rect 26146 79319 26202 79328
rect 23386 64152 23442 64161
rect 23386 64087 23442 64096
rect 19246 62792 19302 62801
rect 19246 62727 19302 62736
rect 17868 51740 17920 51746
rect 17868 51682 17920 51688
rect 15844 33108 15896 33114
rect 15844 33050 15896 33056
rect 16488 26920 16540 26926
rect 16488 26862 16540 26868
rect 12268 6886 12388 6914
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 12268 3602 12296 6886
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12176 3454 12388 3482
rect 12360 480 12388 3454
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 16500 3534 16528 26862
rect 17880 3534 17908 51682
rect 19260 3534 19288 62727
rect 22006 53136 22062 53145
rect 22006 53071 22062 53080
rect 20628 22772 20680 22778
rect 20628 22714 20680 22720
rect 20536 3596 20588 3602
rect 20536 3538 20588 3544
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 15948 480 15976 3470
rect 17052 480 17080 3470
rect 18248 480 18276 3470
rect 19444 480 19472 3470
rect 20548 1850 20576 3538
rect 20640 3534 20668 22714
rect 22020 6914 22048 53071
rect 23400 6914 23428 64087
rect 21836 6886 22048 6914
rect 23032 6886 23428 6914
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20548 1822 20668 1850
rect 20640 480 20668 1822
rect 21836 480 21864 6886
rect 23032 480 23060 6886
rect 24216 6248 24268 6254
rect 24216 6190 24268 6196
rect 24228 480 24256 6190
rect 26160 3602 26188 79319
rect 30286 72448 30342 72457
rect 30286 72383 30342 72392
rect 28906 35184 28962 35193
rect 28906 35119 28962 35128
rect 28816 17264 28868 17270
rect 28816 17206 28868 17212
rect 26516 8968 26568 8974
rect 26516 8910 26568 8916
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 26148 3596 26200 3602
rect 26148 3538 26200 3544
rect 25332 480 25360 3538
rect 26528 480 26556 8910
rect 28828 3602 28856 17206
rect 27712 3596 27764 3602
rect 27712 3538 27764 3544
rect 28816 3596 28868 3602
rect 28816 3538 28868 3544
rect 27724 480 27752 3538
rect 28920 480 28948 35119
rect 30300 6914 30328 72383
rect 31666 58576 31722 58585
rect 31666 58511 31722 58520
rect 31680 6914 31708 58511
rect 33046 47560 33102 47569
rect 33046 47495 33102 47504
rect 30116 6886 30328 6914
rect 31312 6886 31708 6914
rect 30116 480 30144 6886
rect 31312 480 31340 6886
rect 33060 3602 33088 47495
rect 34440 3602 34468 83399
rect 35176 71913 35204 309742
rect 39316 215286 39344 329967
rect 39960 253230 39988 445703
rect 41340 425746 41368 534006
rect 41328 425740 41380 425746
rect 41328 425682 41380 425688
rect 44008 418810 44036 554746
rect 44086 536072 44142 536081
rect 44086 536007 44142 536016
rect 43996 418804 44048 418810
rect 43996 418746 44048 418752
rect 43994 382936 44050 382945
rect 43994 382871 44050 382880
rect 40684 327752 40736 327758
rect 40684 327694 40736 327700
rect 39948 253224 40000 253230
rect 39948 253166 40000 253172
rect 39304 215280 39356 215286
rect 39304 215222 39356 215228
rect 35162 71904 35218 71913
rect 35162 71839 35218 71848
rect 38566 65512 38622 65521
rect 38566 65447 38622 65456
rect 35806 57216 35862 57225
rect 35806 57151 35862 57160
rect 35820 3602 35848 57151
rect 37188 42152 37240 42158
rect 37188 42094 37240 42100
rect 37096 28348 37148 28354
rect 37096 28290 37148 28296
rect 37108 3602 37136 28290
rect 32404 3596 32456 3602
rect 32404 3538 32456 3544
rect 33048 3596 33100 3602
rect 33048 3538 33100 3544
rect 33600 3596 33652 3602
rect 33600 3538 33652 3544
rect 34428 3596 34480 3602
rect 34428 3538 34480 3544
rect 34796 3596 34848 3602
rect 34796 3538 34848 3544
rect 35808 3596 35860 3602
rect 35808 3538 35860 3544
rect 35992 3596 36044 3602
rect 35992 3538 36044 3544
rect 37096 3596 37148 3602
rect 37096 3538 37148 3544
rect 32416 480 32444 3538
rect 33612 480 33640 3538
rect 34808 480 34836 3538
rect 36004 480 36032 3538
rect 37200 480 37228 42094
rect 38580 6914 38608 65447
rect 40696 59362 40724 327694
rect 44008 262886 44036 382871
rect 44100 380866 44128 536007
rect 48148 442950 48176 569162
rect 48226 539608 48282 539617
rect 48226 539543 48282 539552
rect 48136 442944 48188 442950
rect 48136 442886 48188 442892
rect 46848 433356 46900 433362
rect 46848 433298 46900 433304
rect 44088 380860 44140 380866
rect 44088 380802 44140 380808
rect 43996 262880 44048 262886
rect 43996 262822 44048 262828
rect 46860 235958 46888 433298
rect 48136 402960 48188 402966
rect 48136 402902 48188 402908
rect 48148 343641 48176 402902
rect 48240 393310 48268 539543
rect 50908 525094 50936 582354
rect 53656 565888 53708 565894
rect 53656 565830 53708 565836
rect 52276 563100 52328 563106
rect 52276 563042 52328 563048
rect 50988 545148 51040 545154
rect 50988 545090 51040 545096
rect 51000 529922 51028 545090
rect 50988 529916 51040 529922
rect 50988 529858 51040 529864
rect 50896 525088 50948 525094
rect 50896 525030 50948 525036
rect 49608 508564 49660 508570
rect 49608 508506 49660 508512
rect 48228 393304 48280 393310
rect 48228 393246 48280 393252
rect 48134 343632 48190 343641
rect 48134 343567 48190 343576
rect 48148 245614 48176 343567
rect 48228 325712 48280 325718
rect 48228 325654 48280 325660
rect 48136 245608 48188 245614
rect 48136 245550 48188 245556
rect 46848 235952 46900 235958
rect 46848 235894 46900 235900
rect 43442 233880 43498 233889
rect 43442 233815 43498 233824
rect 40684 59356 40736 59362
rect 40684 59298 40736 59304
rect 41328 53100 41380 53106
rect 41328 53042 41380 53048
rect 39948 37936 40000 37942
rect 39948 37878 40000 37884
rect 39960 6914 39988 37878
rect 38396 6886 38608 6914
rect 39592 6886 39988 6914
rect 38396 480 38424 6886
rect 39592 480 39620 6886
rect 41340 3602 41368 53042
rect 43456 45558 43484 233815
rect 48136 69692 48188 69698
rect 48136 69634 48188 69640
rect 43444 45552 43496 45558
rect 43444 45494 43496 45500
rect 44086 43480 44142 43489
rect 44086 43415 44142 43424
rect 42706 11656 42762 11665
rect 42706 11591 42762 11600
rect 42720 3602 42748 11591
rect 44100 3602 44128 43415
rect 46848 40724 46900 40730
rect 46848 40666 46900 40672
rect 45468 20052 45520 20058
rect 45468 19994 45520 20000
rect 45284 13116 45336 13122
rect 45284 13058 45336 13064
rect 40684 3596 40736 3602
rect 40684 3538 40736 3544
rect 41328 3596 41380 3602
rect 41328 3538 41380 3544
rect 41880 3596 41932 3602
rect 41880 3538 41932 3544
rect 42708 3596 42760 3602
rect 42708 3538 42760 3544
rect 43076 3596 43128 3602
rect 43076 3538 43128 3544
rect 44088 3596 44140 3602
rect 44088 3538 44140 3544
rect 44272 3596 44324 3602
rect 44272 3538 44324 3544
rect 40696 480 40724 3538
rect 41892 480 41920 3538
rect 43088 480 43116 3538
rect 44284 480 44312 3538
rect 45296 3482 45324 13058
rect 45480 6914 45508 19994
rect 46860 6914 46888 40666
rect 48148 6914 48176 69634
rect 48240 54505 48268 325654
rect 49620 240145 49648 508506
rect 50804 450016 50856 450022
rect 50804 449958 50856 449964
rect 50816 331226 50844 449958
rect 50908 449206 50936 525030
rect 50896 449200 50948 449206
rect 50896 449142 50948 449148
rect 51000 402974 51028 529858
rect 52184 517540 52236 517546
rect 52184 517482 52236 517488
rect 50908 402946 51028 402974
rect 52196 402966 52224 517482
rect 52288 431254 52316 563042
rect 52368 546508 52420 546514
rect 52368 546450 52420 546456
rect 52380 518906 52408 546450
rect 52368 518900 52420 518906
rect 52368 518842 52420 518848
rect 52380 517546 52408 518842
rect 52368 517540 52420 517546
rect 52368 517482 52420 517488
rect 52368 460216 52420 460222
rect 52368 460158 52420 460164
rect 52276 431248 52328 431254
rect 52276 431190 52328 431196
rect 52276 421592 52328 421598
rect 52276 421534 52328 421540
rect 52184 402960 52236 402966
rect 50908 400926 50936 402946
rect 52184 402902 52236 402908
rect 52196 402286 52224 402902
rect 52184 402280 52236 402286
rect 52184 402222 52236 402228
rect 50896 400920 50948 400926
rect 50896 400862 50948 400868
rect 50528 331220 50580 331226
rect 50528 331162 50580 331168
rect 50804 331220 50856 331226
rect 50804 331162 50856 331168
rect 50540 330546 50568 331162
rect 50528 330540 50580 330546
rect 50528 330482 50580 330488
rect 49606 240136 49662 240145
rect 49606 240071 49662 240080
rect 50908 238678 50936 400862
rect 52288 373994 52316 421534
rect 52104 373966 52316 373994
rect 52104 372570 52132 373966
rect 52092 372564 52144 372570
rect 52092 372506 52144 372512
rect 50988 331356 51040 331362
rect 50988 331298 51040 331304
rect 50896 238672 50948 238678
rect 50896 238614 50948 238620
rect 50894 66872 50950 66881
rect 50894 66807 50950 66816
rect 48226 54496 48282 54505
rect 48226 54431 48282 54440
rect 49606 39400 49662 39409
rect 49606 39335 49662 39344
rect 45388 6886 45508 6914
rect 46676 6886 46888 6914
rect 47872 6886 48176 6914
rect 45388 3602 45416 6886
rect 45376 3596 45428 3602
rect 45376 3538 45428 3544
rect 45296 3454 45508 3482
rect 45480 480 45508 3454
rect 46676 480 46704 6886
rect 47872 480 47900 6886
rect 49620 3534 49648 39335
rect 50908 3534 50936 66807
rect 51000 17950 51028 331298
rect 52104 314702 52132 372506
rect 52184 334076 52236 334082
rect 52184 334018 52236 334024
rect 52092 314696 52144 314702
rect 52092 314638 52144 314644
rect 52196 278730 52224 334018
rect 52276 331288 52328 331294
rect 52276 331230 52328 331236
rect 52184 278724 52236 278730
rect 52184 278666 52236 278672
rect 51080 261520 51132 261526
rect 51080 261462 51132 261468
rect 51092 260914 51120 261462
rect 51080 260908 51132 260914
rect 51080 260850 51132 260856
rect 52184 260908 52236 260914
rect 52184 260850 52236 260856
rect 52196 232665 52224 260850
rect 52182 232656 52238 232665
rect 52182 232591 52238 232600
rect 52288 26217 52316 331230
rect 52380 50386 52408 460158
rect 53564 444508 53616 444514
rect 53564 444450 53616 444456
rect 53576 372638 53604 444450
rect 53668 436082 53696 565830
rect 55036 543788 55088 543794
rect 55036 543730 55088 543736
rect 53748 519580 53800 519586
rect 53748 519522 53800 519528
rect 53656 436076 53708 436082
rect 53656 436018 53708 436024
rect 53564 372632 53616 372638
rect 53564 372574 53616 372580
rect 53576 292534 53604 372574
rect 53656 340196 53708 340202
rect 53656 340138 53708 340144
rect 53564 292528 53616 292534
rect 53564 292470 53616 292476
rect 52460 262880 52512 262886
rect 52460 262822 52512 262828
rect 52472 262274 52500 262822
rect 52460 262268 52512 262274
rect 52460 262210 52512 262216
rect 53564 262268 53616 262274
rect 53564 262210 53616 262216
rect 53576 198694 53604 262210
rect 53668 241505 53696 340138
rect 53760 319462 53788 519522
rect 55048 399498 55076 543730
rect 55140 457502 55168 587862
rect 59084 586560 59136 586566
rect 59084 586502 59136 586508
rect 57888 585200 57940 585206
rect 57888 585142 57940 585148
rect 55864 564460 55916 564466
rect 55864 564402 55916 564408
rect 55128 457496 55180 457502
rect 55128 457438 55180 457444
rect 55126 444544 55182 444553
rect 55126 444479 55182 444488
rect 55036 399492 55088 399498
rect 55036 399434 55088 399440
rect 55048 379409 55076 399434
rect 55034 379400 55090 379409
rect 55034 379335 55090 379344
rect 54944 360868 54996 360874
rect 54944 360810 54996 360816
rect 53748 319456 53800 319462
rect 53748 319398 53800 319404
rect 53654 241496 53710 241505
rect 53654 241431 53710 241440
rect 53564 198688 53616 198694
rect 53564 198630 53616 198636
rect 53760 75177 53788 319398
rect 54956 318102 54984 360810
rect 54944 318096 54996 318102
rect 54944 318038 54996 318044
rect 54944 270564 54996 270570
rect 54944 270506 54996 270512
rect 54852 264988 54904 264994
rect 54852 264930 54904 264936
rect 54864 186289 54892 264930
rect 54956 199442 54984 270506
rect 55048 237386 55076 379335
rect 55140 264246 55168 444479
rect 55876 433294 55904 564402
rect 57796 554056 57848 554062
rect 57796 553998 57848 554004
rect 56508 459604 56560 459610
rect 56508 459546 56560 459552
rect 55864 433288 55916 433294
rect 55864 433230 55916 433236
rect 56322 373280 56378 373289
rect 56322 373215 56378 373224
rect 56336 299470 56364 373215
rect 56520 366382 56548 459546
rect 57704 453348 57756 453354
rect 57704 453290 57756 453296
rect 57716 385014 57744 453290
rect 57808 416090 57836 553998
rect 57900 447817 57928 585142
rect 59096 468518 59124 586502
rect 61936 579692 61988 579698
rect 61936 579634 61988 579640
rect 61844 574116 61896 574122
rect 61844 574058 61896 574064
rect 59176 558340 59228 558346
rect 59176 558282 59228 558288
rect 59084 468512 59136 468518
rect 59084 468454 59136 468460
rect 57886 447808 57942 447817
rect 57886 447743 57942 447752
rect 57888 436076 57940 436082
rect 57888 436018 57940 436024
rect 57900 434790 57928 436018
rect 57888 434784 57940 434790
rect 57888 434726 57940 434732
rect 57796 416084 57848 416090
rect 57796 416026 57848 416032
rect 57796 414724 57848 414730
rect 57796 414666 57848 414672
rect 57704 385008 57756 385014
rect 57704 384950 57756 384956
rect 56508 366376 56560 366382
rect 56508 366318 56560 366324
rect 57702 347032 57758 347041
rect 57702 346967 57758 346976
rect 57610 336016 57666 336025
rect 57610 335951 57666 335960
rect 56508 314696 56560 314702
rect 56508 314638 56560 314644
rect 56416 305040 56468 305046
rect 56416 304982 56468 304988
rect 56324 299464 56376 299470
rect 56324 299406 56376 299412
rect 55128 264240 55180 264246
rect 55128 264182 55180 264188
rect 55036 237380 55088 237386
rect 55036 237322 55088 237328
rect 56428 222057 56456 304982
rect 56414 222048 56470 222057
rect 56414 221983 56470 221992
rect 56520 219337 56548 314638
rect 57624 287026 57652 335951
rect 57612 287020 57664 287026
rect 57612 286962 57664 286968
rect 57612 260976 57664 260982
rect 57612 260918 57664 260924
rect 56506 219328 56562 219337
rect 56506 219263 56562 219272
rect 54944 199436 54996 199442
rect 54944 199378 54996 199384
rect 57624 193186 57652 260918
rect 57716 235890 57744 346967
rect 57808 241466 57836 414666
rect 57900 298110 57928 434726
rect 59084 425740 59136 425746
rect 59084 425682 59136 425688
rect 59096 425134 59124 425682
rect 59084 425128 59136 425134
rect 59084 425070 59136 425076
rect 59096 374678 59124 425070
rect 59188 421598 59216 558282
rect 60648 549296 60700 549302
rect 60648 549238 60700 549244
rect 59268 547936 59320 547942
rect 59268 547878 59320 547884
rect 59176 421592 59228 421598
rect 59176 421534 59228 421540
rect 59176 418804 59228 418810
rect 59176 418746 59228 418752
rect 59188 416838 59216 418746
rect 59176 416832 59228 416838
rect 59176 416774 59228 416780
rect 59188 396030 59216 416774
rect 59280 405822 59308 547878
rect 60660 522986 60688 549238
rect 60648 522980 60700 522986
rect 60648 522922 60700 522928
rect 60464 440292 60516 440298
rect 60464 440234 60516 440240
rect 59268 405816 59320 405822
rect 59268 405758 59320 405764
rect 59176 396024 59228 396030
rect 59176 395966 59228 395972
rect 59084 374672 59136 374678
rect 59084 374614 59136 374620
rect 58990 334656 59046 334665
rect 58990 334591 59046 334600
rect 59004 302190 59032 334591
rect 59082 332616 59138 332625
rect 59082 332551 59138 332560
rect 58992 302184 59044 302190
rect 58992 302126 59044 302132
rect 57888 298104 57940 298110
rect 57888 298046 57940 298052
rect 58992 298104 59044 298110
rect 58992 298046 59044 298052
rect 59004 297430 59032 298046
rect 58992 297424 59044 297430
rect 58992 297366 59044 297372
rect 57888 284368 57940 284374
rect 57888 284310 57940 284316
rect 57796 241460 57848 241466
rect 57796 241402 57848 241408
rect 57704 235884 57756 235890
rect 57704 235826 57756 235832
rect 57612 193180 57664 193186
rect 57612 193122 57664 193128
rect 54850 186280 54906 186289
rect 54850 186215 54906 186224
rect 53746 75168 53802 75177
rect 53746 75103 53802 75112
rect 53746 68232 53802 68241
rect 53746 68167 53802 68176
rect 52368 50380 52420 50386
rect 52368 50322 52420 50328
rect 53654 50280 53710 50289
rect 53654 50215 53710 50224
rect 52274 26208 52330 26217
rect 52274 26143 52330 26152
rect 50988 17944 51040 17950
rect 50988 17886 51040 17892
rect 53668 3534 53696 50215
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 49608 3528 49660 3534
rect 49608 3470 49660 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50896 3528 50948 3534
rect 50896 3470 50948 3476
rect 52552 3528 52604 3534
rect 52552 3470 52604 3476
rect 53656 3528 53708 3534
rect 53656 3470 53708 3476
rect 48976 480 49004 3470
rect 50172 480 50200 3470
rect 51356 2168 51408 2174
rect 51356 2110 51408 2116
rect 51368 480 51396 2110
rect 52564 480 52592 3470
rect 53760 480 53788 68167
rect 57794 59936 57850 59945
rect 57794 59871 57850 59880
rect 54484 36576 54536 36582
rect 54484 36518 54536 36524
rect 54496 3602 54524 36518
rect 56508 29640 56560 29646
rect 56508 29582 56560 29588
rect 54944 10328 54996 10334
rect 54944 10270 54996 10276
rect 54484 3596 54536 3602
rect 54484 3538 54536 3544
rect 54956 480 54984 10270
rect 56520 3534 56548 29582
rect 57808 3534 57836 59871
rect 57900 21418 57928 284310
rect 59004 230489 59032 297366
rect 58990 230480 59046 230489
rect 58990 230415 59046 230424
rect 59096 222193 59124 332551
rect 59188 291106 59216 395966
rect 59266 371376 59322 371385
rect 59266 371311 59322 371320
rect 59176 291100 59228 291106
rect 59176 291042 59228 291048
rect 59176 282940 59228 282946
rect 59176 282882 59228 282888
rect 59082 222184 59138 222193
rect 59082 222119 59138 222128
rect 59188 220794 59216 282882
rect 59280 244254 59308 371311
rect 60372 342916 60424 342922
rect 60372 342858 60424 342864
rect 60384 314634 60412 342858
rect 60476 338201 60504 440234
rect 60660 407182 60688 522922
rect 61856 456113 61884 574058
rect 61948 525162 61976 579634
rect 62040 558346 62068 702986
rect 67640 702704 67692 702710
rect 67640 702646 67692 702652
rect 66168 699712 66220 699718
rect 66168 699654 66220 699660
rect 65982 590744 66038 590753
rect 65982 590679 66038 590688
rect 64696 581052 64748 581058
rect 64696 580994 64748 581000
rect 63316 571396 63368 571402
rect 63316 571338 63368 571344
rect 62028 558340 62080 558346
rect 62028 558282 62080 558288
rect 62040 557598 62068 558282
rect 62028 557592 62080 557598
rect 62028 557534 62080 557540
rect 61936 525156 61988 525162
rect 61936 525098 61988 525104
rect 61936 504416 61988 504422
rect 61936 504358 61988 504364
rect 61842 456104 61898 456113
rect 61842 456039 61898 456048
rect 61752 453416 61804 453422
rect 61752 453358 61804 453364
rect 60648 407176 60700 407182
rect 60648 407118 60700 407124
rect 60556 378208 60608 378214
rect 60556 378150 60608 378156
rect 60462 338192 60518 338201
rect 60462 338127 60518 338136
rect 60464 332648 60516 332654
rect 60464 332590 60516 332596
rect 60372 314628 60424 314634
rect 60372 314570 60424 314576
rect 60476 291174 60504 332590
rect 60464 291168 60516 291174
rect 60464 291110 60516 291116
rect 60280 278792 60332 278798
rect 60280 278734 60332 278740
rect 60096 253224 60148 253230
rect 60096 253166 60148 253172
rect 60108 252618 60136 253166
rect 60096 252612 60148 252618
rect 60096 252554 60148 252560
rect 59268 244248 59320 244254
rect 59268 244190 59320 244196
rect 60292 233918 60320 278734
rect 60568 277370 60596 378150
rect 60660 376038 60688 407118
rect 61764 391377 61792 453358
rect 61844 423700 61896 423706
rect 61844 423642 61896 423648
rect 61750 391368 61806 391377
rect 61750 391303 61806 391312
rect 60648 376032 60700 376038
rect 60648 375974 60700 375980
rect 60646 374096 60702 374105
rect 60646 374031 60702 374040
rect 60556 277364 60608 277370
rect 60556 277306 60608 277312
rect 60464 255332 60516 255338
rect 60464 255274 60516 255280
rect 60372 252612 60424 252618
rect 60372 252554 60424 252560
rect 60280 233912 60332 233918
rect 60280 233854 60332 233860
rect 60384 223417 60412 252554
rect 60370 223408 60426 223417
rect 60370 223343 60426 223352
rect 59176 220788 59228 220794
rect 59176 220730 59228 220736
rect 60476 220114 60504 255274
rect 60660 247042 60688 374031
rect 61660 365016 61712 365022
rect 61660 364958 61712 364964
rect 61672 287054 61700 364958
rect 61856 362234 61884 423642
rect 61844 362228 61896 362234
rect 61844 362170 61896 362176
rect 61750 338328 61806 338337
rect 61750 338263 61806 338272
rect 61764 307766 61792 338263
rect 61752 307760 61804 307766
rect 61752 307702 61804 307708
rect 61672 287026 61884 287054
rect 61856 276078 61884 287026
rect 61844 276072 61896 276078
rect 61844 276014 61896 276020
rect 61384 258052 61436 258058
rect 61384 257994 61436 258000
rect 60648 247036 60700 247042
rect 60648 246978 60700 246984
rect 60464 220108 60516 220114
rect 60464 220050 60516 220056
rect 60648 128376 60700 128382
rect 60648 128318 60700 128324
rect 60660 91798 60688 128318
rect 60648 91792 60700 91798
rect 60648 91734 60700 91740
rect 59268 61396 59320 61402
rect 59268 61338 59320 61344
rect 57888 21412 57940 21418
rect 57888 21354 57940 21360
rect 59280 3534 59308 61338
rect 61396 33794 61424 257994
rect 61856 194546 61884 276014
rect 61948 274650 61976 504358
rect 63224 461644 63276 461650
rect 63224 461586 63276 461592
rect 62028 456068 62080 456074
rect 62028 456010 62080 456016
rect 62040 386374 62068 456010
rect 63132 405816 63184 405822
rect 63132 405758 63184 405764
rect 62028 386368 62080 386374
rect 62028 386310 62080 386316
rect 63144 356794 63172 405758
rect 63236 391241 63264 461586
rect 63328 454714 63356 571338
rect 64708 530602 64736 580994
rect 65890 573472 65946 573481
rect 65890 573407 65946 573416
rect 64788 567248 64840 567254
rect 64788 567190 64840 567196
rect 64696 530596 64748 530602
rect 64696 530538 64748 530544
rect 63408 520940 63460 520946
rect 63408 520882 63460 520888
rect 63316 454708 63368 454714
rect 63316 454650 63368 454656
rect 63316 437572 63368 437578
rect 63316 437514 63368 437520
rect 63222 391232 63278 391241
rect 63222 391167 63278 391176
rect 63328 384334 63356 437514
rect 63316 384328 63368 384334
rect 63316 384270 63368 384276
rect 63314 363760 63370 363769
rect 63314 363695 63370 363704
rect 63132 356788 63184 356794
rect 63132 356730 63184 356736
rect 62762 338192 62818 338201
rect 62762 338127 62818 338136
rect 62026 331936 62082 331945
rect 62026 331871 62082 331880
rect 61936 274644 61988 274650
rect 61936 274586 61988 274592
rect 61936 271176 61988 271182
rect 61936 271118 61988 271124
rect 61948 232558 61976 271118
rect 61936 232552 61988 232558
rect 61936 232494 61988 232500
rect 61844 194540 61896 194546
rect 61844 194482 61896 194488
rect 61936 35216 61988 35222
rect 61936 35158 61988 35164
rect 61384 33788 61436 33794
rect 61384 33730 61436 33736
rect 60004 31068 60056 31074
rect 60004 31010 60056 31016
rect 59636 7676 59688 7682
rect 59636 7618 59688 7624
rect 56048 3528 56100 3534
rect 56048 3470 56100 3476
rect 56508 3528 56560 3534
rect 56508 3470 56560 3476
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 57796 3528 57848 3534
rect 57796 3470 57848 3476
rect 58440 3528 58492 3534
rect 58440 3470 58492 3476
rect 59268 3528 59320 3534
rect 59268 3470 59320 3476
rect 56060 480 56088 3470
rect 57256 480 57284 3470
rect 58452 480 58480 3470
rect 59648 480 59676 7618
rect 60016 2174 60044 31010
rect 61948 3534 61976 35158
rect 62040 32434 62068 331871
rect 62776 309806 62804 338127
rect 62764 309800 62816 309806
rect 62764 309742 62816 309748
rect 63132 271924 63184 271930
rect 63132 271866 63184 271872
rect 62120 264240 62172 264246
rect 62120 264182 62172 264188
rect 62132 263634 62160 264182
rect 62120 263628 62172 263634
rect 62120 263570 62172 263576
rect 63144 242049 63172 271866
rect 63328 269074 63356 363695
rect 63420 285734 63448 520882
rect 64694 454744 64750 454753
rect 64694 454679 64750 454688
rect 64604 447840 64656 447846
rect 64604 447782 64656 447788
rect 64616 389162 64644 447782
rect 64604 389156 64656 389162
rect 64604 389098 64656 389104
rect 64708 388929 64736 454679
rect 64800 437578 64828 567190
rect 65904 539714 65932 573407
rect 65892 539708 65944 539714
rect 65892 539650 65944 539656
rect 65996 463010 66024 590679
rect 66074 559600 66130 559609
rect 66074 559535 66130 559544
rect 65984 463004 66036 463010
rect 65984 462946 66036 462952
rect 65984 446412 66036 446418
rect 65984 446354 66036 446360
rect 64788 437572 64840 437578
rect 64788 437514 64840 437520
rect 65892 431248 65944 431254
rect 65892 431190 65944 431196
rect 65800 393304 65852 393310
rect 65798 393272 65800 393281
rect 65852 393272 65854 393281
rect 65798 393207 65854 393216
rect 64694 388920 64750 388929
rect 64694 388855 64750 388864
rect 64788 387116 64840 387122
rect 64788 387058 64840 387064
rect 64604 346452 64656 346458
rect 64604 346394 64656 346400
rect 64512 334620 64564 334626
rect 64512 334562 64564 334568
rect 64144 318096 64196 318102
rect 64144 318038 64196 318044
rect 64156 289270 64184 318038
rect 64524 316742 64552 334562
rect 64616 318646 64644 346394
rect 64696 336796 64748 336802
rect 64696 336738 64748 336744
rect 64604 318640 64656 318646
rect 64604 318582 64656 318588
rect 64512 316736 64564 316742
rect 64512 316678 64564 316684
rect 64708 303618 64736 336738
rect 64800 322930 64828 387058
rect 65904 376689 65932 431190
rect 65996 389230 66024 446354
rect 66088 424289 66116 559535
rect 66180 539034 66208 699654
rect 67456 599004 67508 599010
rect 67456 598946 67508 598952
rect 67364 592680 67416 592686
rect 67364 592622 67416 592628
rect 66810 588432 66866 588441
rect 66810 588367 66866 588376
rect 66824 587926 66852 588367
rect 66812 587920 66864 587926
rect 66812 587862 66864 587868
rect 66260 586560 66312 586566
rect 66258 586528 66260 586537
rect 66312 586528 66314 586537
rect 66258 586463 66314 586472
rect 66902 585712 66958 585721
rect 66902 585647 66958 585656
rect 66916 585206 66944 585647
rect 66904 585200 66956 585206
rect 66904 585142 66956 585148
rect 66810 582992 66866 583001
rect 66810 582927 66866 582936
rect 66824 582418 66852 582927
rect 66812 582412 66864 582418
rect 66812 582354 66864 582360
rect 66534 581768 66590 581777
rect 66534 581703 66590 581712
rect 66548 581058 66576 581703
rect 66536 581052 66588 581058
rect 66536 580994 66588 581000
rect 66810 580272 66866 580281
rect 66810 580207 66866 580216
rect 66824 579698 66852 580207
rect 66812 579692 66864 579698
rect 66812 579634 66864 579640
rect 66810 576192 66866 576201
rect 66810 576127 66866 576136
rect 66824 575550 66852 576127
rect 66812 575544 66864 575550
rect 66812 575486 66864 575492
rect 67376 574977 67404 592622
rect 67362 574968 67418 574977
rect 67362 574903 67418 574912
rect 67376 574122 67404 574903
rect 67364 574116 67416 574122
rect 67364 574058 67416 574064
rect 66810 572112 66866 572121
rect 66810 572047 66866 572056
rect 66824 571402 66852 572047
rect 66812 571396 66864 571402
rect 66812 571338 66864 571344
rect 67468 570761 67496 598946
rect 67548 587920 67600 587926
rect 67548 587862 67600 587868
rect 67086 570752 67142 570761
rect 67086 570687 67142 570696
rect 67454 570752 67510 570761
rect 67454 570687 67510 570696
rect 67100 569226 67128 570687
rect 67362 569392 67418 569401
rect 67362 569327 67418 569336
rect 67088 569220 67140 569226
rect 67088 569162 67140 569168
rect 66810 568032 66866 568041
rect 66810 567967 66866 567976
rect 66824 567254 66852 567967
rect 66812 567248 66864 567254
rect 66812 567190 66864 567196
rect 66810 565040 66866 565049
rect 66810 564975 66866 564984
rect 66824 564466 66852 564975
rect 66812 564460 66864 564466
rect 66812 564402 66864 564408
rect 66810 563680 66866 563689
rect 66810 563615 66866 563624
rect 66824 563106 66852 563615
rect 66812 563100 66864 563106
rect 66812 563042 66864 563048
rect 66810 562320 66866 562329
rect 66810 562255 66866 562264
rect 66824 561746 66852 562255
rect 66812 561740 66864 561746
rect 66812 561682 66864 561688
rect 66810 560960 66866 560969
rect 66810 560895 66866 560904
rect 66824 560318 66852 560895
rect 66812 560312 66864 560318
rect 66812 560254 66864 560260
rect 66810 558240 66866 558249
rect 66810 558175 66866 558184
rect 66824 557598 66852 558175
rect 66812 557592 66864 557598
rect 66812 557534 66864 557540
rect 66810 555520 66866 555529
rect 66810 555455 66866 555464
rect 66824 554810 66852 555455
rect 66812 554804 66864 554810
rect 66812 554746 66864 554752
rect 66626 554160 66682 554169
rect 66626 554095 66682 554104
rect 66640 554062 66668 554095
rect 66628 554056 66680 554062
rect 66628 553998 66680 554004
rect 66810 550080 66866 550089
rect 66810 550015 66866 550024
rect 66824 549302 66852 550015
rect 66812 549296 66864 549302
rect 66812 549238 66864 549244
rect 66810 548720 66866 548729
rect 66810 548655 66866 548664
rect 66824 547942 66852 548655
rect 66812 547936 66864 547942
rect 66812 547878 66864 547884
rect 66810 547360 66866 547369
rect 66810 547295 66866 547304
rect 66824 546514 66852 547295
rect 66812 546508 66864 546514
rect 66812 546450 66864 546456
rect 66810 546000 66866 546009
rect 66810 545935 66866 545944
rect 66824 545154 66852 545935
rect 66812 545148 66864 545154
rect 66812 545090 66864 545096
rect 66810 544640 66866 544649
rect 66810 544575 66866 544584
rect 66824 543794 66852 544575
rect 66812 543788 66864 543794
rect 66812 543730 66864 543736
rect 66810 543280 66866 543289
rect 66810 543215 66866 543224
rect 66824 542434 66852 543215
rect 67376 543017 67404 569327
rect 67560 554169 67588 587862
rect 67652 566681 67680 702646
rect 72988 699718 73016 703520
rect 79324 702636 79376 702642
rect 79324 702578 79376 702584
rect 75184 700324 75236 700330
rect 75184 700266 75236 700272
rect 72976 699712 73028 699718
rect 72976 699654 73028 699660
rect 70308 596216 70360 596222
rect 70308 596158 70360 596164
rect 69112 591320 69164 591326
rect 69112 591262 69164 591268
rect 69124 590782 69152 591262
rect 69112 590776 69164 590782
rect 70320 590753 70348 596158
rect 75196 592686 75224 700266
rect 76746 593464 76802 593473
rect 76746 593399 76802 593408
rect 75184 592680 75236 592686
rect 75184 592622 75236 592628
rect 75644 592136 75696 592142
rect 73986 592104 74042 592113
rect 75644 592078 75696 592084
rect 73986 592039 74042 592048
rect 72148 590844 72200 590850
rect 72148 590786 72200 590792
rect 71688 590776 71740 590782
rect 69112 590718 69164 590724
rect 70306 590744 70362 590753
rect 69124 589084 69152 590718
rect 70124 590708 70176 590714
rect 70306 590679 70362 590688
rect 71134 590744 71190 590753
rect 71688 590718 71740 590724
rect 71134 590679 71190 590688
rect 70124 590650 70176 590656
rect 70136 589084 70164 590650
rect 71148 589084 71176 590679
rect 71700 590034 71728 590718
rect 71688 590028 71740 590034
rect 71688 589970 71740 589976
rect 72160 589084 72188 590786
rect 73066 590744 73122 590753
rect 73066 590679 73122 590688
rect 73080 589084 73108 590679
rect 74000 589084 74028 592039
rect 74448 590708 74500 590714
rect 74448 590650 74500 590656
rect 74460 589937 74488 590650
rect 75656 589966 75684 592078
rect 74908 589960 74960 589966
rect 74446 589928 74502 589937
rect 74908 589902 74960 589908
rect 75644 589960 75696 589966
rect 75644 589902 75696 589908
rect 74446 589863 74502 589872
rect 74920 589354 74948 589902
rect 74908 589348 74960 589354
rect 74908 589290 74960 589296
rect 74920 589084 74948 589290
rect 76760 589084 76788 593399
rect 79336 591530 79364 702578
rect 88248 702568 88300 702574
rect 88248 702510 88300 702516
rect 86868 699712 86920 699718
rect 86868 699654 86920 699660
rect 82820 597576 82872 597582
rect 82820 597518 82872 597524
rect 79968 596828 80020 596834
rect 79968 596770 80020 596776
rect 79324 591524 79376 591530
rect 79324 591466 79376 591472
rect 79980 590850 80008 596770
rect 80704 591524 80756 591530
rect 80704 591466 80756 591472
rect 79968 590844 80020 590850
rect 79968 590786 80020 590792
rect 78588 590776 78640 590782
rect 78588 590718 78640 590724
rect 77666 589384 77722 589393
rect 77666 589319 77722 589328
rect 77680 589084 77708 589319
rect 78600 589084 78628 590718
rect 80716 589966 80744 591466
rect 82266 591016 82322 591025
rect 82266 590951 82322 590960
rect 81898 590744 81954 590753
rect 81898 590679 81954 590688
rect 80704 589960 80756 589966
rect 80704 589902 80756 589908
rect 80716 589098 80744 589902
rect 81346 589520 81402 589529
rect 81346 589455 81402 589464
rect 80454 589070 80744 589098
rect 81360 589084 81388 589455
rect 79690 588704 79746 588713
rect 79534 588662 79690 588690
rect 79690 588639 79746 588648
rect 81912 588606 81940 590679
rect 82280 589084 82308 590951
rect 82832 589098 82860 597518
rect 86880 596834 86908 699654
rect 86868 596828 86920 596834
rect 86868 596770 86920 596776
rect 85948 594856 86000 594862
rect 85948 594798 86000 594804
rect 84108 592068 84160 592074
rect 84108 592010 84160 592016
rect 82832 589070 83122 589098
rect 84120 589084 84148 592010
rect 85028 590708 85080 590714
rect 85028 590650 85080 590656
rect 85040 589084 85068 590650
rect 85960 589084 85988 594798
rect 88260 593434 88288 702510
rect 88800 702500 88852 702506
rect 88800 702442 88852 702448
rect 88812 596174 88840 702442
rect 89180 699718 89208 703520
rect 95148 702636 95200 702642
rect 95148 702578 95200 702584
rect 93768 702500 93820 702506
rect 93768 702442 93820 702448
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 90364 605872 90416 605878
rect 90364 605814 90416 605820
rect 88812 596146 88932 596174
rect 88248 593428 88300 593434
rect 88248 593370 88300 593376
rect 86866 590880 86922 590889
rect 86866 590815 86922 590824
rect 86880 589084 86908 590815
rect 88260 590714 88288 593370
rect 88248 590708 88300 590714
rect 88248 590650 88300 590656
rect 81900 588600 81952 588606
rect 75854 588526 76144 588554
rect 88062 588568 88118 588577
rect 81900 588542 81952 588548
rect 87814 588526 88062 588554
rect 76116 588470 76144 588526
rect 88062 588503 88118 588512
rect 76104 588464 76156 588470
rect 76104 588406 76156 588412
rect 88734 588390 88840 588418
rect 88812 587178 88840 588390
rect 88800 587172 88852 587178
rect 88800 587114 88852 587120
rect 67730 584352 67786 584361
rect 67730 584287 67786 584296
rect 67638 566672 67694 566681
rect 67638 566607 67694 566616
rect 67652 565894 67680 566607
rect 67640 565888 67692 565894
rect 67640 565830 67692 565836
rect 67546 554160 67602 554169
rect 67546 554095 67602 554104
rect 67454 552800 67510 552809
rect 67454 552735 67510 552744
rect 67362 543008 67418 543017
rect 67362 542943 67418 542952
rect 66812 542428 66864 542434
rect 66812 542370 66864 542376
rect 66994 541920 67050 541929
rect 66994 541855 67050 541864
rect 67364 541884 67416 541890
rect 67008 541686 67036 541855
rect 67364 541826 67416 541832
rect 66996 541680 67048 541686
rect 66996 541622 67048 541628
rect 67272 541680 67324 541686
rect 67272 541622 67324 541628
rect 66168 539028 66220 539034
rect 66168 538970 66220 538976
rect 66902 452568 66958 452577
rect 66902 452503 66958 452512
rect 66168 451988 66220 451994
rect 66168 451930 66220 451936
rect 66074 424280 66130 424289
rect 66074 424215 66130 424224
rect 66088 423706 66116 424215
rect 66076 423700 66128 423706
rect 66076 423642 66128 423648
rect 66076 396024 66128 396030
rect 66076 395966 66128 395972
rect 66088 390522 66116 395966
rect 66076 390516 66128 390522
rect 66076 390458 66128 390464
rect 65984 389224 66036 389230
rect 65984 389166 66036 389172
rect 66180 387705 66208 451930
rect 66916 440298 66944 452503
rect 66904 440292 66956 440298
rect 66904 440234 66956 440240
rect 66916 440065 66944 440234
rect 66902 440056 66958 440065
rect 66902 439991 66958 440000
rect 66902 437744 66958 437753
rect 66902 437679 66958 437688
rect 66916 437578 66944 437679
rect 66904 437572 66956 437578
rect 66904 437514 66956 437520
rect 66902 435296 66958 435305
rect 66902 435231 66958 435240
rect 66916 434790 66944 435231
rect 66904 434784 66956 434790
rect 66904 434726 66956 434732
rect 66812 433288 66864 433294
rect 66810 433256 66812 433265
rect 66864 433256 66866 433265
rect 66810 433191 66866 433200
rect 66536 431248 66588 431254
rect 66536 431190 66588 431196
rect 66548 431089 66576 431190
rect 66534 431080 66590 431089
rect 66534 431015 66590 431024
rect 66720 429140 66772 429146
rect 66720 429082 66772 429088
rect 66732 428641 66760 429082
rect 66718 428632 66774 428641
rect 66718 428567 66774 428576
rect 66258 426320 66314 426329
rect 66258 426255 66314 426264
rect 66272 425134 66300 426255
rect 66260 425128 66312 425134
rect 66260 425070 66312 425076
rect 66258 421968 66314 421977
rect 66258 421903 66314 421912
rect 66272 421598 66300 421903
rect 66260 421592 66312 421598
rect 66260 421534 66312 421540
rect 66902 417344 66958 417353
rect 66902 417279 66958 417288
rect 66916 416838 66944 417279
rect 66904 416832 66956 416838
rect 66904 416774 66956 416780
rect 66260 416084 66312 416090
rect 66260 416026 66312 416032
rect 66272 415177 66300 416026
rect 66258 415168 66314 415177
rect 66258 415103 66314 415112
rect 66272 414730 66300 415103
rect 66260 414724 66312 414730
rect 66260 414666 66312 414672
rect 66350 408368 66406 408377
rect 66350 408303 66406 408312
rect 66364 407182 66392 408303
rect 66352 407176 66404 407182
rect 66352 407118 66404 407124
rect 66810 406192 66866 406201
rect 66810 406127 66866 406136
rect 66824 405822 66852 406127
rect 66812 405816 66864 405822
rect 66812 405758 66864 405764
rect 66626 403744 66682 403753
rect 66626 403679 66682 403688
rect 66640 403170 66668 403679
rect 66628 403164 66680 403170
rect 66628 403106 66680 403112
rect 66810 401568 66866 401577
rect 66810 401503 66866 401512
rect 66824 400926 66852 401503
rect 66812 400920 66864 400926
rect 66812 400862 66864 400868
rect 66810 399528 66866 399537
rect 66810 399463 66812 399472
rect 66864 399463 66866 399472
rect 66812 399434 66864 399440
rect 66994 396944 67050 396953
rect 66994 396879 67050 396888
rect 67008 396778 67036 396879
rect 66996 396772 67048 396778
rect 66996 396714 67048 396720
rect 67284 396001 67312 541622
rect 67376 539481 67404 541826
rect 67362 539472 67418 539481
rect 67362 539407 67418 539416
rect 67376 410553 67404 539407
rect 67468 412865 67496 552735
rect 67546 551440 67602 551449
rect 67546 551375 67602 551384
rect 67560 541890 67588 551375
rect 67548 541884 67600 541890
rect 67548 541826 67600 541832
rect 67546 540560 67602 540569
rect 67546 540495 67602 540504
rect 67560 539617 67588 540495
rect 67546 539608 67602 539617
rect 67546 539543 67602 539552
rect 67560 537538 67588 539543
rect 67548 537532 67600 537538
rect 67548 537474 67600 537480
rect 67744 459610 67772 584287
rect 88904 582374 88932 596146
rect 89812 594108 89864 594114
rect 89812 594050 89864 594056
rect 89076 590028 89128 590034
rect 89076 589970 89128 589976
rect 88984 588192 89036 588198
rect 88984 588134 89036 588140
rect 88996 586634 89024 588134
rect 88984 586628 89036 586634
rect 88984 586570 89036 586576
rect 89088 582374 89116 589970
rect 89718 586256 89774 586265
rect 89718 586191 89774 586200
rect 88812 582346 88932 582374
rect 88996 582346 89116 582374
rect 67822 577552 67878 577561
rect 67822 577487 67878 577496
rect 67836 467838 67864 577487
rect 88812 576854 88840 582346
rect 88812 576826 88932 576854
rect 88904 560153 88932 576826
rect 88890 560144 88946 560153
rect 88890 560079 88946 560088
rect 88798 540152 88854 540161
rect 88798 540087 88854 540096
rect 88812 539714 88840 540087
rect 88800 539708 88852 539714
rect 88800 539650 88852 539656
rect 70400 539640 70452 539646
rect 81348 539640 81400 539646
rect 70452 539588 70610 539594
rect 70400 539582 70610 539588
rect 81348 539582 81400 539588
rect 69848 539572 69900 539578
rect 69848 539514 69900 539520
rect 70412 539566 70610 539582
rect 68664 539294 68770 539322
rect 69584 539294 69690 539322
rect 68664 536722 68692 539294
rect 69584 536790 69612 539294
rect 69572 536784 69624 536790
rect 69572 536726 69624 536732
rect 68652 536716 68704 536722
rect 68652 536658 68704 536664
rect 67824 467832 67876 467838
rect 67824 467774 67876 467780
rect 67732 459604 67784 459610
rect 67732 459546 67784 459552
rect 67744 458862 67772 459546
rect 67732 458856 67784 458862
rect 67732 458798 67784 458804
rect 67640 454708 67692 454714
rect 67640 454650 67692 454656
rect 67652 445738 67680 454650
rect 68100 450560 68152 450566
rect 68100 450502 68152 450508
rect 68112 449954 68140 450502
rect 68100 449948 68152 449954
rect 68100 449890 68152 449896
rect 68560 449948 68612 449954
rect 68560 449890 68612 449896
rect 67640 445732 67692 445738
rect 67640 445674 67692 445680
rect 67732 442944 67784 442950
rect 67732 442886 67784 442892
rect 67744 442241 67772 442886
rect 67730 442232 67786 442241
rect 67730 442167 67786 442176
rect 67454 412856 67510 412865
rect 67454 412791 67510 412800
rect 67362 410544 67418 410553
rect 67362 410479 67418 410488
rect 67362 396944 67418 396953
rect 67362 396879 67418 396888
rect 67270 395992 67326 396001
rect 67270 395927 67326 395936
rect 66166 387696 66222 387705
rect 66166 387631 66222 387640
rect 67376 376718 67404 396879
rect 66904 376712 66956 376718
rect 65890 376680 65946 376689
rect 66904 376654 66956 376660
rect 67364 376712 67416 376718
rect 67364 376654 67416 376660
rect 65890 376615 65946 376624
rect 66916 375426 66944 376654
rect 66904 375420 66956 375426
rect 66904 375362 66956 375368
rect 65982 351928 66038 351937
rect 65982 351863 66038 351872
rect 64788 322924 64840 322930
rect 64788 322866 64840 322872
rect 65800 322924 65852 322930
rect 65800 322866 65852 322872
rect 65812 322454 65840 322866
rect 65800 322448 65852 322454
rect 65800 322390 65852 322396
rect 64696 303612 64748 303618
rect 64696 303554 64748 303560
rect 64696 300892 64748 300898
rect 64696 300834 64748 300840
rect 64144 289264 64196 289270
rect 64144 289206 64196 289212
rect 63408 285728 63460 285734
rect 63408 285670 63460 285676
rect 63316 269068 63368 269074
rect 63316 269010 63368 269016
rect 63224 263628 63276 263634
rect 63224 263570 63276 263576
rect 63130 242040 63186 242049
rect 63130 241975 63186 241984
rect 63236 231849 63264 263570
rect 63316 253972 63368 253978
rect 63316 253914 63368 253920
rect 63222 231840 63278 231849
rect 63222 231775 63278 231784
rect 63328 208321 63356 253914
rect 63420 209710 63448 285670
rect 64512 256760 64564 256766
rect 64512 256702 64564 256708
rect 64524 228410 64552 256702
rect 64604 245676 64656 245682
rect 64604 245618 64656 245624
rect 64512 228404 64564 228410
rect 64512 228346 64564 228352
rect 64616 212498 64644 245618
rect 64708 237969 64736 300834
rect 64788 269068 64840 269074
rect 64788 269010 64840 269016
rect 64800 267918 64828 269010
rect 64788 267912 64840 267918
rect 64788 267854 64840 267860
rect 64694 237960 64750 237969
rect 64694 237895 64750 237904
rect 64604 212492 64656 212498
rect 64604 212434 64656 212440
rect 63408 209704 63460 209710
rect 63408 209646 63460 209652
rect 63314 208312 63370 208321
rect 63314 208247 63370 208256
rect 64800 197334 64828 267854
rect 65812 240009 65840 322390
rect 65996 305289 66024 351863
rect 66076 346520 66128 346526
rect 66076 346462 66128 346468
rect 65982 305280 66038 305289
rect 65982 305215 66038 305224
rect 66088 294409 66116 346462
rect 66916 346458 66944 375362
rect 67362 347848 67418 347857
rect 67362 347783 67418 347792
rect 66904 346452 66956 346458
rect 66904 346394 66956 346400
rect 67272 346452 67324 346458
rect 67272 346394 67324 346400
rect 67284 345817 67312 346394
rect 67270 345808 67326 345817
rect 67270 345743 67326 345752
rect 66168 333260 66220 333266
rect 66168 333202 66220 333208
rect 66180 312905 66208 333202
rect 67272 329724 67324 329730
rect 67272 329666 67324 329672
rect 66258 326768 66314 326777
rect 66258 326703 66314 326712
rect 66272 325718 66300 326703
rect 66260 325712 66312 325718
rect 66260 325654 66312 325660
rect 67284 324601 67312 329666
rect 67270 324592 67326 324601
rect 67270 324527 67326 324536
rect 66536 322448 66588 322454
rect 66534 322416 66536 322425
rect 66588 322416 66590 322425
rect 66534 322351 66590 322360
rect 66812 321564 66864 321570
rect 66812 321506 66864 321512
rect 66824 320249 66852 321506
rect 66810 320240 66866 320249
rect 66810 320175 66866 320184
rect 66444 319456 66496 319462
rect 66444 319398 66496 319404
rect 66456 319161 66484 319398
rect 66442 319152 66498 319161
rect 66442 319087 66498 319096
rect 66444 318640 66496 318646
rect 66444 318582 66496 318588
rect 66456 318073 66484 318582
rect 66442 318064 66498 318073
rect 66442 317999 66498 318008
rect 66902 316976 66958 316985
rect 66902 316911 66958 316920
rect 66916 316742 66944 316911
rect 66904 316736 66956 316742
rect 66904 316678 66956 316684
rect 66810 314800 66866 314809
rect 66810 314735 66866 314744
rect 66824 314702 66852 314735
rect 66812 314696 66864 314702
rect 66812 314638 66864 314644
rect 66904 314628 66956 314634
rect 66904 314570 66956 314576
rect 66916 313993 66944 314570
rect 66902 313984 66958 313993
rect 66902 313919 66958 313928
rect 66166 312896 66222 312905
rect 66166 312831 66222 312840
rect 66994 311808 67050 311817
rect 66994 311743 67050 311752
rect 66812 309800 66864 309806
rect 66812 309742 66864 309748
rect 66824 309641 66852 309742
rect 66810 309632 66866 309641
rect 66810 309567 66866 309576
rect 66904 307760 66956 307766
rect 66904 307702 66956 307708
rect 66916 307465 66944 307702
rect 66902 307456 66958 307465
rect 66902 307391 66958 307400
rect 66810 306368 66866 306377
rect 66810 306303 66866 306312
rect 66824 305046 66852 306303
rect 66812 305040 66864 305046
rect 66812 304982 66864 304988
rect 66904 303612 66956 303618
rect 66904 303554 66956 303560
rect 66916 303113 66944 303554
rect 66902 303104 66958 303113
rect 66902 303039 66958 303048
rect 66904 302184 66956 302190
rect 66904 302126 66956 302132
rect 66810 302016 66866 302025
rect 66810 301951 66866 301960
rect 66824 300898 66852 301951
rect 66916 300937 66944 302126
rect 66902 300928 66958 300937
rect 66812 300892 66864 300898
rect 66902 300863 66958 300872
rect 66812 300834 66864 300840
rect 66628 299464 66680 299470
rect 66628 299406 66680 299412
rect 66640 298761 66668 299406
rect 66626 298752 66682 298761
rect 66626 298687 66682 298696
rect 66810 297664 66866 297673
rect 66810 297599 66866 297608
rect 66824 297430 66852 297599
rect 66812 297424 66864 297430
rect 66812 297366 66864 297372
rect 67008 296714 67036 311743
rect 67088 311160 67140 311166
rect 67088 311102 67140 311108
rect 67100 310729 67128 311102
rect 67086 310720 67142 310729
rect 67086 310655 67142 310664
rect 66916 296686 67036 296714
rect 66074 294400 66130 294409
rect 66074 294335 66130 294344
rect 66812 293956 66864 293962
rect 66812 293898 66864 293904
rect 66824 293321 66852 293898
rect 66810 293312 66866 293321
rect 66810 293247 66866 293256
rect 66812 292528 66864 292534
rect 66812 292470 66864 292476
rect 66824 292233 66852 292470
rect 66810 292224 66866 292233
rect 66810 292159 66866 292168
rect 66352 291168 66404 291174
rect 66352 291110 66404 291116
rect 66364 290057 66392 291110
rect 66350 290048 66406 290057
rect 66350 289983 66406 289992
rect 66812 289264 66864 289270
rect 66812 289206 66864 289212
rect 66824 288969 66852 289206
rect 66810 288960 66866 288969
rect 66810 288895 66866 288904
rect 66168 287836 66220 287842
rect 66168 287778 66220 287784
rect 66180 277394 66208 287778
rect 66812 287020 66864 287026
rect 66812 286962 66864 286968
rect 66258 286784 66314 286793
rect 66258 286719 66314 286728
rect 66272 285734 66300 286719
rect 66260 285728 66312 285734
rect 66824 285705 66852 286962
rect 66260 285670 66312 285676
rect 66810 285696 66866 285705
rect 66810 285631 66866 285640
rect 66810 284608 66866 284617
rect 66810 284543 66866 284552
rect 66824 284374 66852 284543
rect 66812 284368 66864 284374
rect 66812 284310 66864 284316
rect 66810 283520 66866 283529
rect 66810 283455 66866 283464
rect 66824 282946 66852 283455
rect 66812 282940 66864 282946
rect 66812 282882 66864 282888
rect 66626 279168 66682 279177
rect 66626 279103 66682 279112
rect 66640 278798 66668 279103
rect 66628 278792 66680 278798
rect 66628 278734 66680 278740
rect 66812 278724 66864 278730
rect 66812 278666 66864 278672
rect 66824 278089 66852 278666
rect 66810 278080 66866 278089
rect 66810 278015 66866 278024
rect 66088 277366 66208 277394
rect 65892 274644 65944 274650
rect 65892 274586 65944 274592
rect 65904 274553 65932 274586
rect 65890 274544 65946 274553
rect 65890 274479 65946 274488
rect 65904 274145 65932 274479
rect 65890 274136 65946 274145
rect 65890 274071 65946 274080
rect 65982 259856 66038 259865
rect 65982 259791 66038 259800
rect 65892 251796 65944 251802
rect 65892 251738 65944 251744
rect 65798 240000 65854 240009
rect 65798 239935 65854 239944
rect 65904 231130 65932 251738
rect 65996 232529 66024 259791
rect 65982 232520 66038 232529
rect 65982 232455 66038 232464
rect 65892 231124 65944 231130
rect 65892 231066 65944 231072
rect 66088 226953 66116 277366
rect 66260 277364 66312 277370
rect 66260 277306 66312 277312
rect 66272 276185 66300 277306
rect 66810 277264 66866 277273
rect 66810 277199 66866 277208
rect 66258 276176 66314 276185
rect 66258 276111 66314 276120
rect 66824 276078 66852 277199
rect 66812 276072 66864 276078
rect 66812 276014 66864 276020
rect 66258 272912 66314 272921
rect 66258 272847 66314 272856
rect 66272 271930 66300 272847
rect 66260 271924 66312 271930
rect 66260 271866 66312 271872
rect 66916 271182 66944 296686
rect 67178 296168 67234 296177
rect 67178 296103 67234 296112
rect 67192 295390 67220 296103
rect 67180 295384 67232 295390
rect 67180 295326 67232 295332
rect 67086 291136 67142 291145
rect 67086 291071 67088 291080
rect 67140 291071 67142 291080
rect 67088 291042 67140 291048
rect 67376 287881 67404 347783
rect 67468 311166 67496 412791
rect 67546 395992 67602 396001
rect 67546 395927 67602 395936
rect 67560 394913 67588 395927
rect 67546 394904 67602 394913
rect 67546 394839 67602 394848
rect 67560 380934 67588 394839
rect 67548 380928 67600 380934
rect 67548 380870 67600 380876
rect 67456 311160 67508 311166
rect 67456 311102 67508 311108
rect 67560 299849 67588 380870
rect 67744 367878 67772 442167
rect 68572 390289 68600 449890
rect 68664 390402 68692 536658
rect 69584 535537 69612 536726
rect 69570 535528 69626 535537
rect 69570 535463 69626 535472
rect 69860 456822 69888 539514
rect 69020 456816 69072 456822
rect 69020 456758 69072 456764
rect 69848 456816 69900 456822
rect 69848 456758 69900 456764
rect 68744 445732 68796 445738
rect 68744 445674 68796 445680
rect 68756 444394 68784 445674
rect 68928 444440 68980 444446
rect 68756 444388 68928 444394
rect 68756 444382 68980 444388
rect 69032 444394 69060 456758
rect 70412 446457 70440 539566
rect 70780 539294 71530 539322
rect 72542 539294 72648 539322
rect 70780 528554 70808 539294
rect 72424 539028 72476 539034
rect 72424 538970 72476 538976
rect 70504 528526 70808 528554
rect 70504 526590 70532 528526
rect 70492 526584 70544 526590
rect 70492 526526 70544 526532
rect 71044 526584 71096 526590
rect 71044 526526 71096 526532
rect 71056 525842 71084 526526
rect 71044 525836 71096 525842
rect 71044 525778 71096 525784
rect 71056 447846 71084 525778
rect 72436 453354 72464 538970
rect 72620 536761 72648 539294
rect 73172 539294 73370 539322
rect 73540 539294 74290 539322
rect 75104 539294 75210 539322
rect 75932 539294 76130 539322
rect 76760 539294 77050 539322
rect 78062 539294 78352 539322
rect 72606 536752 72662 536761
rect 72606 536687 72662 536696
rect 72620 454753 72648 536687
rect 73172 536081 73200 539294
rect 73158 536072 73214 536081
rect 73158 536007 73214 536016
rect 73540 528554 73568 539294
rect 75104 538214 75132 539294
rect 75104 538186 75224 538214
rect 75196 536654 75224 538186
rect 75184 536648 75236 536654
rect 75184 536590 75236 536596
rect 73264 528526 73568 528554
rect 72606 454744 72662 454753
rect 72606 454679 72662 454688
rect 72424 453348 72476 453354
rect 72424 453290 72476 453296
rect 72700 452668 72752 452674
rect 72700 452610 72752 452616
rect 72712 449886 72740 452610
rect 72700 449880 72752 449886
rect 72700 449822 72752 449828
rect 72712 448594 72740 449822
rect 72700 448588 72752 448594
rect 72700 448530 72752 448536
rect 73160 448588 73212 448594
rect 73160 448530 73212 448536
rect 71044 447840 71096 447846
rect 71044 447782 71096 447788
rect 70398 446448 70454 446457
rect 70398 446383 70454 446392
rect 71778 445904 71834 445913
rect 71778 445839 71834 445848
rect 68756 444380 68968 444382
rect 68770 444366 68968 444380
rect 69032 444366 70242 444394
rect 71792 444380 71820 445839
rect 73172 444380 73200 448530
rect 73264 446418 73292 528526
rect 74540 467832 74592 467838
rect 74540 467774 74592 467780
rect 74552 450022 74580 467774
rect 75196 451994 75224 536590
rect 75932 453422 75960 539294
rect 76760 538966 76788 539294
rect 76748 538960 76800 538966
rect 76748 538902 76800 538908
rect 76562 535392 76618 535401
rect 76562 535327 76618 535336
rect 76576 461514 76604 535327
rect 78324 534750 78352 539294
rect 78784 539294 78890 539322
rect 79520 539294 79810 539322
rect 80822 539294 81112 539322
rect 78312 534744 78364 534750
rect 78312 534686 78364 534692
rect 78680 533384 78732 533390
rect 78680 533326 78732 533332
rect 77944 525156 77996 525162
rect 77944 525098 77996 525104
rect 76012 461508 76064 461514
rect 76012 461450 76064 461456
rect 76564 461508 76616 461514
rect 76564 461450 76616 461456
rect 75920 453416 75972 453422
rect 75920 453358 75972 453364
rect 75184 451988 75236 451994
rect 75184 451930 75236 451936
rect 74540 450016 74592 450022
rect 74540 449958 74592 449964
rect 74816 450016 74868 450022
rect 74816 449958 74868 449964
rect 73252 446412 73304 446418
rect 73252 446354 73304 446360
rect 74828 444380 74856 449958
rect 76024 444394 76052 461450
rect 76576 460970 76604 461450
rect 76564 460964 76616 460970
rect 76564 460906 76616 460912
rect 77956 455326 77984 525098
rect 78692 456074 78720 533326
rect 78784 461650 78812 539294
rect 79520 533390 79548 539294
rect 80058 535800 80114 535809
rect 80058 535735 80114 535744
rect 79508 533384 79560 533390
rect 79508 533326 79560 533332
rect 80072 531298 80100 535735
rect 81084 532098 81112 539294
rect 81360 536722 81388 539582
rect 85580 539572 85632 539578
rect 85580 539514 85632 539520
rect 81544 539294 81650 539322
rect 81820 539294 82570 539322
rect 82832 539294 83490 539322
rect 84304 539294 84410 539322
rect 84580 539294 85330 539322
rect 81348 536716 81400 536722
rect 81348 536658 81400 536664
rect 81544 535634 81572 539294
rect 81532 535628 81584 535634
rect 81532 535570 81584 535576
rect 81072 532092 81124 532098
rect 81072 532034 81124 532040
rect 79980 531282 80100 531298
rect 79324 531276 79376 531282
rect 79324 531218 79376 531224
rect 79968 531276 80100 531282
rect 80020 531270 80100 531276
rect 79968 531218 80020 531224
rect 79336 530602 79364 531218
rect 79324 530596 79376 530602
rect 79324 530538 79376 530544
rect 78772 461644 78824 461650
rect 78772 461586 78824 461592
rect 79336 460934 79364 530538
rect 81820 528554 81848 539294
rect 81452 528526 81848 528554
rect 79336 460906 79456 460934
rect 78680 456068 78732 456074
rect 78680 456010 78732 456016
rect 77300 455320 77352 455326
rect 77300 455262 77352 455268
rect 77944 455320 77996 455326
rect 77944 455262 77996 455268
rect 77312 454170 77340 455262
rect 77300 454164 77352 454170
rect 77300 454106 77352 454112
rect 77312 444394 77340 454106
rect 79428 444553 79456 460906
rect 81452 458969 81480 528526
rect 81438 458960 81494 458969
rect 81438 458895 81494 458904
rect 81440 458856 81492 458862
rect 81440 458798 81492 458804
rect 80888 449200 80940 449206
rect 80888 449142 80940 449148
rect 79414 444544 79470 444553
rect 79414 444479 79470 444488
rect 76024 444366 76314 444394
rect 77312 444366 77786 444394
rect 79428 444380 79456 444479
rect 80900 444380 80928 449142
rect 81452 444394 81480 458798
rect 82832 456113 82860 539294
rect 84304 536518 84332 539294
rect 84292 536512 84344 536518
rect 84292 536454 84344 536460
rect 83464 535628 83516 535634
rect 83464 535570 83516 535576
rect 83476 469849 83504 535570
rect 84580 528554 84608 539294
rect 85592 536654 85620 539514
rect 86342 539294 86632 539322
rect 86604 538214 86632 539294
rect 86972 539294 87354 539322
rect 88366 539294 88656 539322
rect 86604 538186 86908 538214
rect 86880 536790 86908 538186
rect 86868 536784 86920 536790
rect 86868 536726 86920 536732
rect 85580 536648 85632 536654
rect 85580 536590 85632 536596
rect 84212 528526 84608 528554
rect 83462 469840 83518 469849
rect 83462 469775 83518 469784
rect 82818 456104 82874 456113
rect 82818 456039 82874 456048
rect 84212 447817 84240 528526
rect 85580 468512 85632 468518
rect 85580 468454 85632 468460
rect 82818 447808 82874 447817
rect 82818 447743 82874 447752
rect 84198 447808 84254 447817
rect 84198 447743 84254 447752
rect 82832 444553 82860 447743
rect 82818 444544 82874 444553
rect 82818 444479 82874 444488
rect 83830 444544 83886 444553
rect 85592 444514 85620 468454
rect 86880 465769 86908 536726
rect 86866 465760 86922 465769
rect 86866 465695 86922 465704
rect 86972 457609 87000 539294
rect 88628 538218 88656 539294
rect 88616 538212 88668 538218
rect 88616 538154 88668 538160
rect 86958 457600 87014 457609
rect 86958 457535 87014 457544
rect 87604 457496 87656 457502
rect 87604 457438 87656 457444
rect 87616 444961 87644 457438
rect 88996 455462 89024 582346
rect 89626 560144 89682 560153
rect 89626 560079 89682 560088
rect 89640 558958 89668 560079
rect 89628 558952 89680 558958
rect 89628 558894 89680 558900
rect 89628 543788 89680 543794
rect 89628 543730 89680 543736
rect 89640 538218 89668 543730
rect 89628 538212 89680 538218
rect 89628 538154 89680 538160
rect 89076 536512 89128 536518
rect 89076 536454 89128 536460
rect 88340 455456 88392 455462
rect 88340 455398 88392 455404
rect 88984 455456 89036 455462
rect 88984 455398 89036 455404
rect 87602 444952 87658 444961
rect 87602 444887 87658 444896
rect 83830 444479 83886 444488
rect 85580 444508 85632 444514
rect 81452 444366 82386 444394
rect 83844 444380 83872 444479
rect 85580 444450 85632 444456
rect 85592 444380 85620 444450
rect 87616 444394 87644 444887
rect 87078 444366 87644 444394
rect 88352 444394 88380 455398
rect 89088 449177 89116 536454
rect 89640 535498 89668 538154
rect 89628 535492 89680 535498
rect 89628 535434 89680 535440
rect 89732 532030 89760 586191
rect 89824 567361 89852 594050
rect 90376 593842 90404 605814
rect 92480 596828 92532 596834
rect 92480 596770 92532 596776
rect 90364 593836 90416 593842
rect 90364 593778 90416 593784
rect 91192 593836 91244 593842
rect 91192 593778 91244 593784
rect 90362 589928 90418 589937
rect 90362 589863 90418 589872
rect 89810 567352 89866 567361
rect 89810 567287 89866 567296
rect 89824 567254 89852 567287
rect 89812 567248 89864 567254
rect 89812 567190 89864 567196
rect 89720 532024 89772 532030
rect 89720 531966 89772 531972
rect 89074 449168 89130 449177
rect 89074 449103 89130 449112
rect 90376 444689 90404 589863
rect 91098 587616 91154 587625
rect 91098 587551 91154 587560
rect 91112 557530 91140 587551
rect 91204 576745 91232 593778
rect 91282 584896 91338 584905
rect 91282 584831 91338 584840
rect 91296 584458 91324 584831
rect 91284 584452 91336 584458
rect 91284 584394 91336 584400
rect 91836 583704 91888 583710
rect 91834 583672 91836 583681
rect 91888 583672 91890 583681
rect 91834 583607 91890 583616
rect 91282 582176 91338 582185
rect 91282 582111 91338 582120
rect 91296 581058 91324 582111
rect 91284 581052 91336 581058
rect 91284 580994 91336 581000
rect 91282 578096 91338 578105
rect 91282 578031 91338 578040
rect 91296 576910 91324 578031
rect 91284 576904 91336 576910
rect 91284 576846 91336 576852
rect 91190 576736 91246 576745
rect 91190 576671 91246 576680
rect 91204 576162 91232 576671
rect 91192 576156 91244 576162
rect 91192 576098 91244 576104
rect 91742 575376 91798 575385
rect 91742 575311 91798 575320
rect 91756 574122 91784 575311
rect 91744 574116 91796 574122
rect 91744 574058 91796 574064
rect 91742 574016 91798 574025
rect 91742 573951 91798 573960
rect 91756 572762 91784 573951
rect 91744 572756 91796 572762
rect 91744 572698 91796 572704
rect 91742 572656 91798 572665
rect 91742 572591 91798 572600
rect 91192 571464 91244 571470
rect 91190 571432 91192 571441
rect 91244 571432 91246 571441
rect 91756 571402 91784 572591
rect 91190 571367 91246 571376
rect 91744 571396 91796 571402
rect 91744 571338 91796 571344
rect 91742 568712 91798 568721
rect 91742 568647 91798 568656
rect 91560 565888 91612 565894
rect 91558 565856 91560 565865
rect 91612 565856 91614 565865
rect 91558 565791 91614 565800
rect 91558 564496 91614 564505
rect 91558 564431 91560 564440
rect 91612 564431 91614 564440
rect 91560 564402 91612 564408
rect 91558 563136 91614 563145
rect 91558 563071 91560 563080
rect 91612 563071 91614 563080
rect 91560 563042 91612 563048
rect 91190 561504 91246 561513
rect 91190 561439 91246 561448
rect 91100 557524 91152 557530
rect 91100 557466 91152 557472
rect 91098 557424 91154 557433
rect 91098 557359 91154 557368
rect 91112 556238 91140 557359
rect 91100 556232 91152 556238
rect 91100 556174 91152 556180
rect 91098 556064 91154 556073
rect 91098 555999 91154 556008
rect 91112 554810 91140 555999
rect 91100 554804 91152 554810
rect 91100 554746 91152 554752
rect 91100 552152 91152 552158
rect 91098 552120 91100 552129
rect 91152 552120 91154 552129
rect 91098 552055 91154 552064
rect 91098 550760 91154 550769
rect 91098 550695 91154 550704
rect 91112 550662 91140 550695
rect 91100 550656 91152 550662
rect 91100 550598 91152 550604
rect 91098 549400 91154 549409
rect 91098 549335 91154 549344
rect 91112 549302 91140 549335
rect 91100 549296 91152 549302
rect 91100 549238 91152 549244
rect 90456 549228 90508 549234
rect 90456 549170 90508 549176
rect 90468 460222 90496 549170
rect 91098 547768 91154 547777
rect 91098 547703 91154 547712
rect 91112 538898 91140 547703
rect 91100 538892 91152 538898
rect 91100 538834 91152 538840
rect 91204 537606 91232 561439
rect 91284 557524 91336 557530
rect 91284 557466 91336 557472
rect 91296 549234 91324 557466
rect 91374 553344 91430 553353
rect 91374 553279 91430 553288
rect 91388 552090 91416 553279
rect 91376 552084 91428 552090
rect 91376 552026 91428 552032
rect 91284 549228 91336 549234
rect 91284 549170 91336 549176
rect 91284 547936 91336 547942
rect 91282 547904 91284 547913
rect 91336 547904 91338 547913
rect 91282 547839 91338 547848
rect 91558 545184 91614 545193
rect 91558 545119 91560 545128
rect 91612 545119 91614 545128
rect 91560 545090 91612 545096
rect 91558 542464 91614 542473
rect 91558 542399 91560 542408
rect 91612 542399 91614 542408
rect 91560 542370 91612 542376
rect 91192 537600 91244 537606
rect 91192 537542 91244 537548
rect 90548 535492 90600 535498
rect 90548 535434 90600 535440
rect 90560 468489 90588 535434
rect 90546 468480 90602 468489
rect 90546 468415 90602 468424
rect 91560 463004 91612 463010
rect 91560 462946 91612 462952
rect 90456 460216 90508 460222
rect 90456 460158 90508 460164
rect 91572 459610 91600 462946
rect 91100 459604 91152 459610
rect 91100 459546 91152 459552
rect 91560 459604 91612 459610
rect 91560 459546 91612 459552
rect 90362 444680 90418 444689
rect 90362 444615 90418 444624
rect 90376 444394 90404 444615
rect 88352 444366 88458 444394
rect 90206 444366 90404 444394
rect 91112 444394 91140 459546
rect 91756 458862 91784 568647
rect 92294 558784 92350 558793
rect 92294 558719 92350 558728
rect 92308 556850 92336 558719
rect 92296 556844 92348 556850
rect 92296 556786 92348 556792
rect 91926 541104 91982 541113
rect 91926 541039 91982 541048
rect 91940 541006 91968 541039
rect 91928 541000 91980 541006
rect 91928 540942 91980 540948
rect 92388 541000 92440 541006
rect 92388 540942 92440 540948
rect 92400 538937 92428 540942
rect 92386 538928 92442 538937
rect 92386 538863 92442 538872
rect 91744 458856 91796 458862
rect 91744 458798 91796 458804
rect 92492 447001 92520 596770
rect 93124 590776 93176 590782
rect 93124 590718 93176 590724
rect 93136 574802 93164 590718
rect 93780 583778 93808 702442
rect 94504 588600 94556 588606
rect 94504 588542 94556 588548
rect 93768 583772 93820 583778
rect 93768 583714 93820 583720
rect 93124 574796 93176 574802
rect 93124 574738 93176 574744
rect 93122 570072 93178 570081
rect 93122 570007 93178 570016
rect 93136 565146 93164 570007
rect 93124 565140 93176 565146
rect 93124 565082 93176 565088
rect 93766 543824 93822 543833
rect 93766 543759 93822 543768
rect 93122 539744 93178 539753
rect 93122 539679 93178 539688
rect 93136 462913 93164 539679
rect 93780 538801 93808 543759
rect 93766 538792 93822 538801
rect 93766 538727 93822 538736
rect 93122 462904 93178 462913
rect 93122 462839 93178 462848
rect 94516 448526 94544 588542
rect 95160 584458 95188 702578
rect 105464 700330 105492 703520
rect 130384 702840 130436 702846
rect 130384 702782 130436 702788
rect 105452 700324 105504 700330
rect 105452 700266 105504 700272
rect 124864 700324 124916 700330
rect 124864 700266 124916 700272
rect 111156 597576 111208 597582
rect 111156 597518 111208 597524
rect 100758 593464 100814 593473
rect 100758 593399 100814 593408
rect 96620 592136 96672 592142
rect 95882 592104 95938 592113
rect 96620 592078 96672 592084
rect 95882 592039 95938 592048
rect 95148 584452 95200 584458
rect 95148 584394 95200 584400
rect 94596 571464 94648 571470
rect 94596 571406 94648 571412
rect 94608 566506 94636 571406
rect 94596 566500 94648 566506
rect 94596 566442 94648 566448
rect 95240 547936 95292 547942
rect 95240 547878 95292 547884
rect 95252 547194 95280 547878
rect 95240 547188 95292 547194
rect 95240 547130 95292 547136
rect 94594 541104 94650 541113
rect 94594 541039 94650 541048
rect 94608 534721 94636 541039
rect 94594 534712 94650 534721
rect 94594 534647 94650 534656
rect 94608 467129 94636 534647
rect 94594 467120 94650 467129
rect 94594 467055 94650 467064
rect 95896 451246 95924 592039
rect 95976 542428 96028 542434
rect 95976 542370 96028 542376
rect 95988 471209 96016 542370
rect 95974 471200 96030 471209
rect 95974 471135 96030 471144
rect 95884 451240 95936 451246
rect 95884 451182 95936 451188
rect 94504 448520 94556 448526
rect 94504 448462 94556 448468
rect 92478 446992 92534 447001
rect 92478 446927 92534 446936
rect 93030 446992 93086 447001
rect 93030 446927 93086 446936
rect 93044 445777 93072 446927
rect 93030 445768 93086 445777
rect 93030 445703 93086 445712
rect 91112 444366 91586 444394
rect 93044 444380 93072 445703
rect 94516 444825 94544 448462
rect 94502 444816 94558 444825
rect 94502 444751 94558 444760
rect 94516 444394 94544 444751
rect 95896 444394 95924 451182
rect 96632 445913 96660 592078
rect 97262 590880 97318 590889
rect 97262 590815 97318 590824
rect 97276 558210 97304 590815
rect 100666 589520 100722 589529
rect 100666 589455 100722 589464
rect 98642 589384 98698 589393
rect 98642 589319 98698 589328
rect 97264 558204 97316 558210
rect 97264 558146 97316 558152
rect 97908 549296 97960 549302
rect 97908 549238 97960 549244
rect 97264 545148 97316 545154
rect 97264 545090 97316 545096
rect 97276 465769 97304 545090
rect 97262 465760 97318 465769
rect 97262 465695 97318 465704
rect 97920 457473 97948 549238
rect 97906 457464 97962 457473
rect 97906 457399 97962 457408
rect 96618 445904 96674 445913
rect 96618 445839 96674 445848
rect 97630 445904 97686 445913
rect 98656 445874 98684 589319
rect 98736 586628 98788 586634
rect 98736 586570 98788 586576
rect 98748 449993 98776 586570
rect 98734 449984 98790 449993
rect 98734 449919 98790 449928
rect 97630 445839 97686 445848
rect 98644 445868 98696 445874
rect 94516 444366 94714 444394
rect 95896 444366 96186 444394
rect 97644 444380 97672 445839
rect 98644 445810 98696 445816
rect 98748 444394 98776 449919
rect 100680 449206 100708 589455
rect 100668 449200 100720 449206
rect 100668 449142 100720 449148
rect 100484 445868 100536 445874
rect 100484 445810 100536 445816
rect 100496 445777 100524 445810
rect 100482 445768 100538 445777
rect 100482 445703 100538 445712
rect 100772 444514 100800 593399
rect 104162 591016 104218 591025
rect 104162 590951 104218 590960
rect 103520 574796 103572 574802
rect 103520 574738 103572 574744
rect 101404 552152 101456 552158
rect 101404 552094 101456 552100
rect 101416 468489 101444 552094
rect 101402 468480 101458 468489
rect 101402 468415 101458 468424
rect 103532 449954 103560 574738
rect 104176 574190 104204 590951
rect 106924 589960 106976 589966
rect 106924 589902 106976 589908
rect 105542 588704 105598 588713
rect 105542 588639 105598 588648
rect 104164 574184 104216 574190
rect 104164 574126 104216 574132
rect 103520 449948 103572 449954
rect 103520 449890 103572 449896
rect 103704 449948 103756 449954
rect 103704 449890 103756 449896
rect 102232 445868 102284 445874
rect 102232 445810 102284 445816
rect 100760 444508 100812 444514
rect 100760 444450 100812 444456
rect 98748 444366 99130 444394
rect 100772 444380 100800 444450
rect 102244 444380 102272 445810
rect 103716 444380 103744 449890
rect 105556 447137 105584 588639
rect 106188 563100 106240 563106
rect 106188 563042 106240 563048
rect 106200 562358 106228 563042
rect 106188 562352 106240 562358
rect 106188 562294 106240 562300
rect 106188 554804 106240 554810
rect 106188 554746 106240 554752
rect 106200 464370 106228 554746
rect 106188 464364 106240 464370
rect 106188 464306 106240 464312
rect 106936 449886 106964 589902
rect 108304 581052 108356 581058
rect 108304 580994 108356 581000
rect 107016 564460 107068 564466
rect 107016 564402 107068 564408
rect 107028 463010 107056 564402
rect 107016 463004 107068 463010
rect 107016 462946 107068 462952
rect 108316 456074 108344 580994
rect 111064 576904 111116 576910
rect 111064 576846 111116 576852
rect 109684 574184 109736 574190
rect 109684 574126 109736 574132
rect 108396 552084 108448 552090
rect 108396 552026 108448 552032
rect 108408 469849 108436 552026
rect 108394 469840 108450 469849
rect 108394 469775 108450 469784
rect 108304 456068 108356 456074
rect 108304 456010 108356 456016
rect 106924 449880 106976 449886
rect 106924 449822 106976 449828
rect 105542 447128 105598 447137
rect 105542 447063 105598 447072
rect 105556 444394 105584 447063
rect 105478 444366 105584 444394
rect 106936 444380 106964 449822
rect 108304 449200 108356 449206
rect 108304 449142 108356 449148
rect 108316 444380 108344 449142
rect 109696 447098 109724 574126
rect 111076 449177 111104 576846
rect 111168 560318 111196 597518
rect 113180 593428 113232 593434
rect 113180 593370 113232 593376
rect 111800 592068 111852 592074
rect 111800 592010 111852 592016
rect 111156 560312 111208 560318
rect 111156 560254 111208 560260
rect 111708 560312 111760 560318
rect 111708 560254 111760 560260
rect 111062 449168 111118 449177
rect 111062 449103 111118 449112
rect 109684 447092 109736 447098
rect 109684 447034 109736 447040
rect 109696 444961 109724 447034
rect 111720 444961 111748 560254
rect 111812 455394 111840 592010
rect 112444 572756 112496 572762
rect 112444 572698 112496 572704
rect 111800 455388 111852 455394
rect 111800 455330 111852 455336
rect 111812 454714 111840 455330
rect 111800 454708 111852 454714
rect 111800 454650 111852 454656
rect 109682 444952 109738 444961
rect 109682 444887 109738 444896
rect 111706 444952 111762 444961
rect 111706 444887 111762 444896
rect 109696 444394 109724 444887
rect 111720 444394 111748 444887
rect 109696 444366 109802 444394
rect 111550 444366 111748 444394
rect 111812 444394 111840 454650
rect 112456 453354 112484 572698
rect 112444 453348 112496 453354
rect 112444 453290 112496 453296
rect 113192 445777 113220 593370
rect 115204 587172 115256 587178
rect 115204 587114 115256 587120
rect 115216 457502 115244 587114
rect 118698 585712 118754 585721
rect 118698 585647 118754 585656
rect 116584 583772 116636 583778
rect 116584 583714 116636 583720
rect 115204 457496 115256 457502
rect 115204 457438 115256 457444
rect 116596 448662 116624 583714
rect 116676 565888 116728 565894
rect 116676 565830 116728 565836
rect 116688 451994 116716 565830
rect 118516 558204 118568 558210
rect 118516 558146 118568 558152
rect 118528 553450 118556 558146
rect 118516 553444 118568 553450
rect 118516 553386 118568 553392
rect 116676 451988 116728 451994
rect 116676 451930 116728 451936
rect 116584 448656 116636 448662
rect 116122 448624 116178 448633
rect 116584 448598 116636 448604
rect 116122 448559 116178 448568
rect 113178 445768 113234 445777
rect 113178 445703 113234 445712
rect 114374 445768 114430 445777
rect 114374 445703 114430 445712
rect 111812 444366 112930 444394
rect 114388 444380 114416 445703
rect 116136 444380 116164 448559
rect 118528 445777 118556 553386
rect 118712 445806 118740 585647
rect 122840 576156 122892 576162
rect 122840 576098 122892 576104
rect 122196 571396 122248 571402
rect 122196 571338 122248 571344
rect 122104 556232 122156 556238
rect 122104 556174 122156 556180
rect 120816 464364 120868 464370
rect 120816 464306 120868 464312
rect 120632 458856 120684 458862
rect 120632 458798 120684 458804
rect 118700 445800 118752 445806
rect 117594 445768 117650 445777
rect 117594 445703 117650 445712
rect 118514 445768 118570 445777
rect 118700 445742 118752 445748
rect 118514 445703 118570 445712
rect 117608 444380 117636 445703
rect 118712 444394 118740 445742
rect 119344 444576 119396 444582
rect 119344 444518 119396 444524
rect 119356 444394 119384 444518
rect 118712 444366 119384 444394
rect 120644 411097 120672 458798
rect 120724 448656 120776 448662
rect 120724 448598 120776 448604
rect 120736 435985 120764 448598
rect 120722 435976 120778 435985
rect 120722 435911 120778 435920
rect 120736 434790 120764 435911
rect 120724 434784 120776 434790
rect 120724 434726 120776 434732
rect 120722 417072 120778 417081
rect 120722 417007 120778 417016
rect 120630 411088 120686 411097
rect 120630 411023 120686 411032
rect 120736 393990 120764 417007
rect 120724 393984 120776 393990
rect 120724 393926 120776 393932
rect 85854 391096 85910 391105
rect 85606 391068 85854 391082
rect 73068 391060 73120 391066
rect 73068 391002 73120 391008
rect 85592 391054 85854 391068
rect 73080 390590 73108 391002
rect 80058 390960 80114 390969
rect 80058 390895 80114 390904
rect 80610 390960 80666 390969
rect 80666 390918 80914 390946
rect 80610 390895 80666 390904
rect 72056 390584 72108 390590
rect 71870 390552 71926 390561
rect 71806 390510 71870 390538
rect 71926 390532 72056 390538
rect 71926 390526 72108 390532
rect 73068 390584 73120 390590
rect 73068 390526 73120 390532
rect 71926 390510 72096 390526
rect 71870 390487 71926 390496
rect 71884 390427 71912 390487
rect 69938 390416 69994 390425
rect 68664 390388 68770 390402
rect 68664 390374 68784 390388
rect 68558 390280 68614 390289
rect 68558 390215 68614 390224
rect 68756 387122 68784 390374
rect 69994 390388 70334 390402
rect 69994 390374 70348 390388
rect 69938 390351 69994 390360
rect 68744 387116 68796 387122
rect 68744 387058 68796 387064
rect 69662 380216 69718 380225
rect 69662 380151 69718 380160
rect 67732 367872 67784 367878
rect 67732 367814 67784 367820
rect 67824 339516 67876 339522
rect 67824 339458 67876 339464
rect 67638 337240 67694 337249
rect 67638 337175 67694 337184
rect 67652 304201 67680 337175
rect 67732 336728 67784 336734
rect 67732 336670 67784 336676
rect 67744 308553 67772 336670
rect 67836 323513 67864 339458
rect 69676 335354 69704 380151
rect 70320 377534 70348 390374
rect 70308 377528 70360 377534
rect 70308 377470 70360 377476
rect 71688 376032 71740 376038
rect 71688 375974 71740 375980
rect 71700 375465 71728 375974
rect 71686 375456 71742 375465
rect 71686 375391 71742 375400
rect 71596 369164 71648 369170
rect 71596 369106 71648 369112
rect 71042 368520 71098 368529
rect 71042 368455 71098 368464
rect 70582 358864 70638 358873
rect 70582 358799 70638 358808
rect 70596 345014 70624 358799
rect 70596 344986 70808 345014
rect 69756 341556 69808 341562
rect 69756 341498 69808 341504
rect 69400 335326 69704 335354
rect 69400 331362 69428 335326
rect 69388 331356 69440 331362
rect 69388 331298 69440 331304
rect 69400 329474 69428 331298
rect 69768 329730 69796 341498
rect 70676 331832 70728 331838
rect 69846 331800 69902 331809
rect 70676 331774 70728 331780
rect 69846 331735 69902 331744
rect 69756 329724 69808 329730
rect 69756 329666 69808 329672
rect 69860 329474 69888 331735
rect 70032 329792 70084 329798
rect 70032 329734 70084 329740
rect 69000 329446 69428 329474
rect 69736 329446 69888 329474
rect 70044 329361 70072 329734
rect 70688 329474 70716 331774
rect 70472 329446 70716 329474
rect 70780 329474 70808 344986
rect 71056 329798 71084 368455
rect 71608 358873 71636 369106
rect 71594 358864 71650 358873
rect 71594 358799 71650 358808
rect 71700 342990 71728 375391
rect 72424 364472 72476 364478
rect 72424 364414 72476 364420
rect 71688 342984 71740 342990
rect 71688 342926 71740 342932
rect 71778 340912 71834 340921
rect 71778 340847 71834 340856
rect 71792 336734 71820 340847
rect 72238 336832 72294 336841
rect 72238 336767 72294 336776
rect 71780 336728 71832 336734
rect 71780 336670 71832 336676
rect 71044 329792 71096 329798
rect 71044 329734 71096 329740
rect 72252 329474 72280 336767
rect 72436 331838 72464 364414
rect 73080 340921 73108 390526
rect 73172 389162 73200 390388
rect 74552 390374 74842 390402
rect 75932 390374 76314 390402
rect 73160 389156 73212 389162
rect 73160 389098 73212 389104
rect 73172 369170 73200 389098
rect 74552 388929 74580 390374
rect 74538 388920 74594 388929
rect 74538 388855 74594 388864
rect 73160 369164 73212 369170
rect 73160 369106 73212 369112
rect 73804 367804 73856 367810
rect 73804 367746 73856 367752
rect 73158 345672 73214 345681
rect 73158 345607 73214 345616
rect 73066 340912 73122 340921
rect 73066 340847 73122 340856
rect 72976 332172 73028 332178
rect 72976 332114 73028 332120
rect 72424 331832 72476 331838
rect 72424 331774 72476 331780
rect 72988 329474 73016 332114
rect 70780 329446 71208 329474
rect 71944 329446 72280 329474
rect 72680 329446 73016 329474
rect 73172 329474 73200 345607
rect 73250 333296 73306 333305
rect 73250 333231 73306 333240
rect 73264 332625 73292 333231
rect 73250 332616 73306 332625
rect 73250 332551 73306 332560
rect 73816 332178 73844 367746
rect 74552 365022 74580 388855
rect 75932 380866 75960 390374
rect 77864 389230 77892 390388
rect 79336 390374 79442 390402
rect 77852 389224 77904 389230
rect 77852 389166 77904 389172
rect 79336 387705 79364 390374
rect 79322 387696 79378 387705
rect 79322 387631 79378 387640
rect 77944 382968 77996 382974
rect 77944 382910 77996 382916
rect 75920 380860 75972 380866
rect 75920 380802 75972 380808
rect 76564 380860 76616 380866
rect 76564 380802 76616 380808
rect 75184 380248 75236 380254
rect 75184 380190 75236 380196
rect 74540 365016 74592 365022
rect 74540 364958 74592 364964
rect 75196 333305 75224 380190
rect 76576 369170 76604 380802
rect 76564 369164 76616 369170
rect 76564 369106 76616 369112
rect 75826 366344 75882 366353
rect 75826 366279 75882 366288
rect 73986 333296 74042 333305
rect 73986 333231 74042 333240
rect 75182 333296 75238 333305
rect 75182 333231 75238 333240
rect 73804 332172 73856 332178
rect 73804 332114 73856 332120
rect 73172 329446 73416 329474
rect 70030 329352 70086 329361
rect 74000 329338 74028 333231
rect 75840 332353 75868 366279
rect 77208 362976 77260 362982
rect 77208 362918 77260 362924
rect 76562 349752 76618 349761
rect 76562 349687 76618 349696
rect 75182 332344 75238 332353
rect 75182 332279 75238 332288
rect 75826 332344 75882 332353
rect 75826 332279 75882 332288
rect 75196 329497 75224 332279
rect 76576 332178 76604 349687
rect 76656 336116 76708 336122
rect 76656 336058 76708 336064
rect 75828 332172 75880 332178
rect 75828 332114 75880 332120
rect 76564 332172 76616 332178
rect 76564 332114 76616 332120
rect 75182 329488 75238 329497
rect 74888 329446 75182 329474
rect 75840 329474 75868 332114
rect 76668 329474 76696 336058
rect 77220 329474 77248 362918
rect 77392 352640 77444 352646
rect 77392 352582 77444 352588
rect 77404 345014 77432 352582
rect 77404 344986 77892 345014
rect 77668 331832 77720 331838
rect 77668 331774 77720 331780
rect 77680 331294 77708 331774
rect 77668 331288 77720 331294
rect 77668 331230 77720 331236
rect 75624 329446 75868 329474
rect 76360 329446 76696 329474
rect 77096 329446 77248 329474
rect 75182 329423 75238 329432
rect 75196 329363 75224 329423
rect 77680 329338 77708 331230
rect 77864 330426 77892 344986
rect 77956 331838 77984 382910
rect 79336 347177 79364 387631
rect 80072 381585 80100 390895
rect 82096 390374 82386 390402
rect 82096 385014 82124 390374
rect 83936 388793 83964 390388
rect 83922 388784 83978 388793
rect 83922 388719 83978 388728
rect 82084 385008 82136 385014
rect 82084 384950 82136 384956
rect 80058 381576 80114 381585
rect 80058 381511 80114 381520
rect 82096 356726 82124 384950
rect 84108 373312 84160 373318
rect 84108 373254 84160 373260
rect 84120 357649 84148 373254
rect 85592 368393 85620 391054
rect 85854 391031 85910 391040
rect 105082 391096 105138 391105
rect 120828 391082 120856 464306
rect 121460 451920 121512 451926
rect 121460 451862 121512 451868
rect 120908 444576 120960 444582
rect 120908 444518 120960 444524
rect 120920 442921 120948 444518
rect 120906 442912 120962 442921
rect 120906 442847 120962 442856
rect 121472 440230 121500 451862
rect 121550 444816 121606 444825
rect 121550 444751 121606 444760
rect 121564 444417 121592 444751
rect 121550 444408 121606 444417
rect 121550 444343 121606 444352
rect 121460 440224 121512 440230
rect 121460 440166 121512 440172
rect 121472 440065 121500 440166
rect 121458 440056 121514 440065
rect 121458 439991 121514 440000
rect 121460 429140 121512 429146
rect 121460 429082 121512 429088
rect 121472 428505 121500 429082
rect 121458 428496 121514 428505
rect 121458 428431 121514 428440
rect 121182 410544 121238 410553
rect 121182 410479 121238 410488
rect 121196 409902 121224 410479
rect 121184 409896 121236 409902
rect 121184 409838 121236 409844
rect 120908 393984 120960 393990
rect 120908 393926 120960 393932
rect 105138 391054 105584 391082
rect 120474 391068 120856 391082
rect 105082 391031 105138 391040
rect 89810 390416 89866 390425
rect 86972 386374 87000 390388
rect 88536 387870 88564 390388
rect 91282 390416 91338 390425
rect 89866 390374 90114 390402
rect 89810 390351 89866 390360
rect 92754 390416 92810 390425
rect 91338 390388 91678 390402
rect 91338 390374 91692 390388
rect 91282 390351 91338 390360
rect 88524 387864 88576 387870
rect 88524 387806 88576 387812
rect 90364 387864 90416 387870
rect 90364 387806 90416 387812
rect 86960 386368 87012 386374
rect 86960 386310 87012 386316
rect 86868 384396 86920 384402
rect 86868 384338 86920 384344
rect 85578 368384 85634 368393
rect 85578 368319 85634 368328
rect 86222 368384 86278 368393
rect 86222 368319 86278 368328
rect 86236 367169 86264 368319
rect 86222 367160 86278 367169
rect 86222 367095 86278 367104
rect 85488 366376 85540 366382
rect 85488 366318 85540 366324
rect 85500 365809 85528 366318
rect 85486 365800 85542 365809
rect 85486 365735 85542 365744
rect 85394 360224 85450 360233
rect 85394 360159 85450 360168
rect 82910 357640 82966 357649
rect 82910 357575 82966 357584
rect 84106 357640 84162 357649
rect 84106 357575 84162 357584
rect 81624 356720 81676 356726
rect 81624 356662 81676 356668
rect 82084 356720 82136 356726
rect 82084 356662 82136 356668
rect 81348 352572 81400 352578
rect 81348 352514 81400 352520
rect 79968 348424 80020 348430
rect 79968 348366 80020 348372
rect 79322 347168 79378 347177
rect 79322 347103 79378 347112
rect 79980 335354 80008 348366
rect 81072 336048 81124 336054
rect 81072 335990 81124 335996
rect 79704 335326 80008 335354
rect 77944 331832 77996 331838
rect 77944 331774 77996 331780
rect 77864 330398 78168 330426
rect 78140 329474 78168 330398
rect 79704 329474 79732 335326
rect 80336 331560 80388 331566
rect 80336 331502 80388 331508
rect 80348 329474 80376 331502
rect 81084 329474 81112 335990
rect 81360 331566 81388 352514
rect 81636 345014 81664 356662
rect 82924 345014 82952 357575
rect 85408 350606 85436 360159
rect 85500 351218 85528 365735
rect 86236 360913 86264 367095
rect 86222 360904 86278 360913
rect 86222 360839 86278 360848
rect 85488 351212 85540 351218
rect 85488 351154 85540 351160
rect 84384 350600 84436 350606
rect 84384 350542 84436 350548
rect 85396 350600 85448 350606
rect 85396 350542 85448 350548
rect 84396 345014 84424 350542
rect 81636 344986 81848 345014
rect 82924 344986 83136 345014
rect 84396 344986 84608 345014
rect 81438 342272 81494 342281
rect 81438 342207 81494 342216
rect 81348 331560 81400 331566
rect 81348 331502 81400 331508
rect 81452 329746 81480 342207
rect 81452 329718 81526 329746
rect 78140 329446 78568 329474
rect 79304 329446 79732 329474
rect 80040 329446 80376 329474
rect 80776 329446 81112 329474
rect 81498 329460 81526 329718
rect 81820 329474 81848 344986
rect 83002 333296 83058 333305
rect 83002 333231 83058 333240
rect 83016 329474 83044 333231
rect 81820 329446 82248 329474
rect 82800 329446 83044 329474
rect 83108 329474 83136 344986
rect 84108 338768 84160 338774
rect 84108 338710 84160 338716
rect 84120 331945 84148 338710
rect 84106 331936 84162 331945
rect 84106 331871 84162 331880
rect 84120 331242 84148 331871
rect 84120 331214 84240 331242
rect 84212 329746 84240 331214
rect 84212 329718 84286 329746
rect 83108 329446 83536 329474
rect 84258 329460 84286 329718
rect 84580 329474 84608 344986
rect 85580 340944 85632 340950
rect 85580 340886 85632 340892
rect 85592 329474 85620 340886
rect 86880 329474 86908 384338
rect 86972 340202 87000 386310
rect 90376 378049 90404 387806
rect 91664 385801 91692 390374
rect 94226 390416 94282 390425
rect 92810 390374 93532 390402
rect 92754 390351 92810 390360
rect 91650 385792 91706 385801
rect 91650 385727 91706 385736
rect 91098 384296 91154 384305
rect 91098 384231 91154 384240
rect 90362 378040 90418 378049
rect 90362 377975 90418 377984
rect 89628 371884 89680 371890
rect 89628 371826 89680 371832
rect 87604 355360 87656 355366
rect 87604 355302 87656 355308
rect 87144 342984 87196 342990
rect 87144 342926 87196 342932
rect 86960 340196 87012 340202
rect 86960 340138 87012 340144
rect 87156 329746 87184 342926
rect 87616 336122 87644 355302
rect 89536 349172 89588 349178
rect 89536 349114 89588 349120
rect 87604 336116 87656 336122
rect 87604 336058 87656 336064
rect 88248 331628 88300 331634
rect 88248 331570 88300 331576
rect 87156 329718 87230 329746
rect 84580 329446 85008 329474
rect 85592 329446 85744 329474
rect 86480 329446 86908 329474
rect 87202 329460 87230 329718
rect 88260 329474 88288 331570
rect 88984 331492 89036 331498
rect 88984 331434 89036 331440
rect 88996 329474 89024 331434
rect 89548 329474 89576 349114
rect 89640 331498 89668 371826
rect 91008 360936 91060 360942
rect 91008 360878 91060 360884
rect 90364 357536 90416 357542
rect 90364 357478 90416 357484
rect 90376 331634 90404 357478
rect 90914 339552 90970 339561
rect 90914 339487 90970 339496
rect 90928 332178 90956 339487
rect 90456 332172 90508 332178
rect 90456 332114 90508 332120
rect 90916 332172 90968 332178
rect 90916 332114 90968 332120
rect 90364 331628 90416 331634
rect 90364 331570 90416 331576
rect 89628 331492 89680 331498
rect 89628 331434 89680 331440
rect 90468 329474 90496 332114
rect 91020 329474 91048 360878
rect 91112 345014 91140 384231
rect 93504 383654 93532 390374
rect 95882 390416 95938 390425
rect 94282 390374 95004 390402
rect 94226 390351 94282 390360
rect 94976 383654 95004 390374
rect 97354 390416 97410 390425
rect 95938 390388 96278 390402
rect 95938 390374 96292 390388
rect 95882 390351 95938 390360
rect 96264 388550 96292 390374
rect 98826 390416 98882 390425
rect 97410 390388 97750 390402
rect 97410 390374 97764 390388
rect 97354 390351 97410 390360
rect 96252 388544 96304 388550
rect 96252 388486 96304 388492
rect 96264 387841 96292 388486
rect 96250 387832 96306 387841
rect 96250 387767 96306 387776
rect 97736 387025 97764 390374
rect 100666 390416 100722 390425
rect 98882 390374 99328 390402
rect 98826 390351 98882 390360
rect 97722 387016 97778 387025
rect 97722 386951 97778 386960
rect 97264 385076 97316 385082
rect 97264 385018 97316 385024
rect 93504 383626 93716 383654
rect 94976 383626 95096 383654
rect 93688 356153 93716 383626
rect 95068 361729 95096 383626
rect 94502 361720 94558 361729
rect 94502 361655 94558 361664
rect 95054 361720 95110 361729
rect 95054 361655 95110 361664
rect 92478 356144 92534 356153
rect 92478 356079 92534 356088
rect 93674 356144 93730 356153
rect 93674 356079 93730 356088
rect 92492 355434 92520 356079
rect 92480 355428 92532 355434
rect 92480 355370 92532 355376
rect 93768 354748 93820 354754
rect 93768 354690 93820 354696
rect 93122 353424 93178 353433
rect 93122 353359 93178 353368
rect 91112 344986 91968 345014
rect 91836 332172 91888 332178
rect 91836 332114 91888 332120
rect 91848 329474 91876 332114
rect 87952 329446 88288 329474
rect 88688 329446 89024 329474
rect 89424 329446 89576 329474
rect 90160 329446 90496 329474
rect 90896 329446 91048 329474
rect 91632 329446 91876 329474
rect 91940 329474 91968 344986
rect 93136 336054 93164 353359
rect 93214 340096 93270 340105
rect 93214 340031 93270 340040
rect 93124 336048 93176 336054
rect 93124 335990 93176 335996
rect 93228 332178 93256 340031
rect 93780 335354 93808 354690
rect 94516 352646 94544 361655
rect 96526 353968 96582 353977
rect 96526 353903 96582 353912
rect 94504 352640 94556 352646
rect 94504 352582 94556 352588
rect 94044 351212 94096 351218
rect 94044 351154 94096 351160
rect 94056 345014 94084 351154
rect 94056 344986 94268 345014
rect 93504 335326 93808 335354
rect 94136 335368 94188 335374
rect 93216 332172 93268 332178
rect 93216 332114 93268 332120
rect 93504 329474 93532 335326
rect 94136 335310 94188 335316
rect 94148 329474 94176 335310
rect 91940 329446 92368 329474
rect 93104 329446 93532 329474
rect 93840 329446 94176 329474
rect 94240 329474 94268 344986
rect 96436 342984 96488 342990
rect 96436 342926 96488 342932
rect 95608 331560 95660 331566
rect 95608 331502 95660 331508
rect 95620 329474 95648 331502
rect 96448 329474 96476 342926
rect 96540 331566 96568 353903
rect 97276 342922 97304 385018
rect 99194 356688 99250 356697
rect 99194 356623 99250 356632
rect 97908 349852 97960 349858
rect 97908 349794 97960 349800
rect 97264 342916 97316 342922
rect 97264 342858 97316 342864
rect 97814 336152 97870 336161
rect 97814 336087 97870 336096
rect 97080 331764 97132 331770
rect 97080 331706 97132 331712
rect 96528 331560 96580 331566
rect 96528 331502 96580 331508
rect 97092 329474 97120 331706
rect 97828 329474 97856 336087
rect 97920 331770 97948 349794
rect 99104 346452 99156 346458
rect 99104 346394 99156 346400
rect 97908 331764 97960 331770
rect 97908 331706 97960 331712
rect 98552 331492 98604 331498
rect 98552 331434 98604 331440
rect 98564 329474 98592 331434
rect 99116 329474 99144 346394
rect 99208 331498 99236 356623
rect 99300 345710 99328 390374
rect 102138 390416 102194 390425
rect 100722 390388 100878 390402
rect 100722 390374 100892 390388
rect 100666 390351 100722 390360
rect 100864 389065 100892 390374
rect 102194 390388 102350 390402
rect 102194 390374 102364 390388
rect 102138 390351 102194 390360
rect 102336 389065 102364 390374
rect 100850 389056 100906 389065
rect 100850 388991 100906 389000
rect 101862 389056 101918 389065
rect 101862 388991 101918 389000
rect 102322 389056 102378 389065
rect 102322 388991 102378 389000
rect 103334 389056 103390 389065
rect 103334 388991 103390 389000
rect 100482 387832 100538 387841
rect 100482 387767 100538 387776
rect 100496 384402 100524 387767
rect 100484 384396 100536 384402
rect 100484 384338 100536 384344
rect 100666 363080 100722 363089
rect 100666 363015 100722 363024
rect 100680 354674 100708 363015
rect 100680 354657 100800 354674
rect 100666 354648 100800 354657
rect 100722 354646 100800 354648
rect 100666 354583 100722 354592
rect 100666 351248 100722 351257
rect 100666 351183 100722 351192
rect 99288 345704 99340 345710
rect 99288 345646 99340 345652
rect 100576 338224 100628 338230
rect 100576 338166 100628 338172
rect 100588 332178 100616 338166
rect 100024 332172 100076 332178
rect 100024 332114 100076 332120
rect 100576 332172 100628 332178
rect 100576 332114 100628 332120
rect 99196 331492 99248 331498
rect 99196 331434 99248 331440
rect 100036 329474 100064 332114
rect 100680 329474 100708 351183
rect 94240 329446 94576 329474
rect 95312 329446 95648 329474
rect 96048 329446 96476 329474
rect 96784 329446 97120 329474
rect 97520 329446 97856 329474
rect 98256 329446 98592 329474
rect 98992 329446 99144 329474
rect 99728 329446 100064 329474
rect 100464 329446 100708 329474
rect 100772 329474 100800 354646
rect 101876 353394 101904 388991
rect 103348 380186 103376 388991
rect 103716 388929 103744 390388
rect 103702 388920 103758 388929
rect 103702 388855 103758 388864
rect 105556 386481 105584 391054
rect 120460 391054 120856 391068
rect 115754 390688 115810 390697
rect 115754 390623 115810 390632
rect 109682 390552 109738 390561
rect 109738 390524 109802 390538
rect 109738 390510 109816 390524
rect 109682 390487 109738 390496
rect 106554 390416 106610 390425
rect 108026 390416 108082 390425
rect 106610 390374 107332 390402
rect 106554 390351 106610 390360
rect 105542 386472 105598 386481
rect 105542 386407 105598 386416
rect 104162 385656 104218 385665
rect 104162 385591 104218 385600
rect 103426 383072 103482 383081
rect 103426 383007 103482 383016
rect 103336 380180 103388 380186
rect 103336 380122 103388 380128
rect 101954 360360 102010 360369
rect 101954 360295 102010 360304
rect 101864 353388 101916 353394
rect 101864 353330 101916 353336
rect 101876 349761 101904 353330
rect 101862 349752 101918 349761
rect 101862 349687 101918 349696
rect 101968 329746 101996 360295
rect 103440 354793 103468 383007
rect 102138 354784 102194 354793
rect 102138 354719 102194 354728
rect 103426 354784 103482 354793
rect 103426 354719 103482 354728
rect 102152 345014 102180 354719
rect 102152 344986 102272 345014
rect 101922 329718 101996 329746
rect 100772 329446 101200 329474
rect 101922 329460 101950 329718
rect 102244 329474 102272 344986
rect 104176 338774 104204 385591
rect 105556 381546 105584 386407
rect 107304 383654 107332 390374
rect 108082 390374 108804 390402
rect 108026 390351 108082 390360
rect 108776 383654 108804 390374
rect 109788 389201 109816 390510
rect 109774 389192 109830 389201
rect 109774 389127 109830 389136
rect 110328 388476 110380 388482
rect 110328 388418 110380 388424
rect 110340 387870 110368 388418
rect 111444 387870 111472 390388
rect 112916 389065 112944 390388
rect 112902 389056 112958 389065
rect 112902 388991 112958 389000
rect 110328 387864 110380 387870
rect 110328 387806 110380 387812
rect 111432 387864 111484 387870
rect 111432 387806 111484 387812
rect 107304 383626 107516 383654
rect 108776 383626 108988 383654
rect 105544 381540 105596 381546
rect 105544 381482 105596 381488
rect 104900 358828 104952 358834
rect 104900 358770 104952 358776
rect 104164 338768 104216 338774
rect 104164 338710 104216 338716
rect 103704 338156 103756 338162
rect 103704 338098 103756 338104
rect 103244 331900 103296 331906
rect 103244 331842 103296 331848
rect 102244 329446 102672 329474
rect 74000 329310 74152 329338
rect 77680 329310 77832 329338
rect 70030 329287 70086 329296
rect 94240 329118 94268 329446
rect 103256 329202 103284 331842
rect 103716 329474 103744 338098
rect 104912 329746 104940 358770
rect 106186 349888 106242 349897
rect 106186 349823 106242 349832
rect 106200 335354 106228 349823
rect 106924 347812 106976 347818
rect 106924 347754 106976 347760
rect 104866 329718 104940 329746
rect 106016 335326 106228 335354
rect 103716 329446 104144 329474
rect 104866 329460 104894 329718
rect 106016 329474 106044 335326
rect 106936 334626 106964 347754
rect 107488 343097 107516 383626
rect 108960 363633 108988 383626
rect 110340 381546 110368 387806
rect 113088 387116 113140 387122
rect 113088 387058 113140 387064
rect 110328 381540 110380 381546
rect 110328 381482 110380 381488
rect 112444 374740 112496 374746
rect 112444 374682 112496 374688
rect 111062 369880 111118 369889
rect 111062 369815 111118 369824
rect 108946 363624 109002 363633
rect 108946 363559 109002 363568
rect 108304 356788 108356 356794
rect 108304 356730 108356 356736
rect 108316 346361 108344 356730
rect 111076 354674 111104 369815
rect 112456 360874 112484 374682
rect 112444 360868 112496 360874
rect 112444 360810 112496 360816
rect 113100 360262 113128 387058
rect 114388 386345 114416 390388
rect 115204 389156 115256 389162
rect 115204 389098 115256 389104
rect 113178 386336 113234 386345
rect 113178 386271 113234 386280
rect 114374 386336 114430 386345
rect 114374 386271 114430 386280
rect 113192 380254 113220 386271
rect 113180 380248 113232 380254
rect 113180 380190 113232 380196
rect 114558 373416 114614 373425
rect 114558 373351 114614 373360
rect 114466 367704 114522 367713
rect 114466 367639 114522 367648
rect 111800 360256 111852 360262
rect 111800 360198 111852 360204
rect 113088 360256 113140 360262
rect 114480 360233 114508 367639
rect 113088 360198 113140 360204
rect 113178 360224 113234 360233
rect 110984 354646 111104 354674
rect 110328 351960 110380 351966
rect 110328 351902 110380 351908
rect 107750 346352 107806 346361
rect 107750 346287 107806 346296
rect 108302 346352 108358 346361
rect 108302 346287 108358 346296
rect 107764 345137 107792 346287
rect 107750 345128 107806 345137
rect 107750 345063 107806 345072
rect 107764 345014 107792 345063
rect 107764 344986 107976 345014
rect 107474 343088 107530 343097
rect 107474 343023 107530 343032
rect 107476 340196 107528 340202
rect 107476 340138 107528 340144
rect 106924 334620 106976 334626
rect 106924 334562 106976 334568
rect 106646 334112 106702 334121
rect 106646 334047 106702 334056
rect 106660 329474 106688 334047
rect 107488 329474 107516 340138
rect 107842 333024 107898 333033
rect 107842 332959 107898 332968
rect 107856 329474 107884 332959
rect 105616 329446 106044 329474
rect 106352 329446 106688 329474
rect 107088 329446 107516 329474
rect 107640 329446 107884 329474
rect 107948 329474 107976 344986
rect 109682 338464 109738 338473
rect 109682 338399 109738 338408
rect 109696 333305 109724 338399
rect 109682 333296 109738 333305
rect 109682 333231 109738 333240
rect 110142 333296 110198 333305
rect 110142 333231 110198 333240
rect 109408 331356 109460 331362
rect 109408 331298 109460 331304
rect 109420 329474 109448 331298
rect 110156 329474 110184 333231
rect 110340 331362 110368 351902
rect 110420 349104 110472 349110
rect 110420 349046 110472 349052
rect 110432 347857 110460 349046
rect 110984 348430 111012 354646
rect 111156 351212 111208 351218
rect 111156 351154 111208 351160
rect 110972 348424 111024 348430
rect 110972 348366 111024 348372
rect 110418 347848 110474 347857
rect 110418 347783 110474 347792
rect 111168 342990 111196 351154
rect 111156 342984 111208 342990
rect 111156 342926 111208 342932
rect 111708 342304 111760 342310
rect 111708 342246 111760 342252
rect 111614 341456 111670 341465
rect 111614 341391 111670 341400
rect 111628 332178 111656 341391
rect 110880 332172 110932 332178
rect 110880 332114 110932 332120
rect 111616 332172 111668 332178
rect 111616 332114 111668 332120
rect 110328 331356 110380 331362
rect 110328 331298 110380 331304
rect 110892 329474 110920 332114
rect 111720 329474 111748 342246
rect 107948 329446 108376 329474
rect 109112 329446 109448 329474
rect 109848 329446 110184 329474
rect 110584 329446 110920 329474
rect 111320 329446 111748 329474
rect 111812 329474 111840 360198
rect 113178 360159 113234 360168
rect 114466 360224 114522 360233
rect 114466 360159 114522 360168
rect 113088 335436 113140 335442
rect 113088 335378 113140 335384
rect 113100 329474 113128 335378
rect 111812 329446 112056 329474
rect 112792 329446 113128 329474
rect 113192 329474 113220 360159
rect 114468 336864 114520 336870
rect 114468 336806 114520 336812
rect 114480 329474 114508 336806
rect 113192 329446 113528 329474
rect 114264 329446 114508 329474
rect 114572 329474 114600 373351
rect 115216 373318 115244 389098
rect 115768 383654 115796 390623
rect 115938 390416 115994 390425
rect 117870 390416 117926 390425
rect 115994 390388 116150 390402
rect 117622 390388 117870 390402
rect 115994 390374 116164 390388
rect 115938 390351 115994 390360
rect 116136 389065 116164 390374
rect 117608 390374 117870 390388
rect 116122 389056 116178 389065
rect 116122 388991 116178 389000
rect 117134 389056 117190 389065
rect 117134 388991 117190 389000
rect 115768 383626 115888 383654
rect 115204 373312 115256 373318
rect 115204 373254 115256 373260
rect 114652 365832 114704 365838
rect 114652 365774 114704 365780
rect 114664 360942 114692 365774
rect 114652 360936 114704 360942
rect 114652 360878 114704 360884
rect 115860 345014 115888 383626
rect 117148 377913 117176 388991
rect 117318 388920 117374 388929
rect 117318 388855 117374 388864
rect 117332 386442 117360 388855
rect 117320 386436 117372 386442
rect 117320 386378 117372 386384
rect 117608 385694 117636 390374
rect 117870 390351 117926 390360
rect 118988 388929 119016 390388
rect 120460 389162 120488 391054
rect 120448 389156 120500 389162
rect 120448 389098 120500 389104
rect 118974 388920 119030 388929
rect 118974 388855 119030 388864
rect 120920 387122 120948 393926
rect 120908 387116 120960 387122
rect 120908 387058 120960 387064
rect 117964 386436 118016 386442
rect 117964 386378 118016 386384
rect 117596 385688 117648 385694
rect 117596 385630 117648 385636
rect 117976 378826 118004 386378
rect 119986 385792 120042 385801
rect 119986 385727 120042 385736
rect 120000 382294 120028 385727
rect 119988 382288 120040 382294
rect 119988 382230 120040 382236
rect 117964 378820 118016 378826
rect 117964 378762 118016 378768
rect 116582 377904 116638 377913
rect 116582 377839 116638 377848
rect 117134 377904 117190 377913
rect 117134 377839 117190 377848
rect 116596 376961 116624 377839
rect 116582 376952 116638 376961
rect 116582 376887 116638 376896
rect 115768 344986 115888 345014
rect 115768 342378 115796 344986
rect 116596 344321 116624 376887
rect 118516 365764 118568 365770
rect 118516 365706 118568 365712
rect 118528 364313 118556 365706
rect 118606 365664 118662 365673
rect 118606 365599 118662 365608
rect 118620 364449 118648 365599
rect 118606 364440 118662 364449
rect 118606 364375 118662 364384
rect 118514 364304 118570 364313
rect 118514 364239 118570 364248
rect 116582 344312 116638 344321
rect 116582 344247 116638 344256
rect 118330 343768 118386 343777
rect 118330 343703 118386 343712
rect 115848 343664 115900 343670
rect 115846 343632 115848 343641
rect 115900 343632 115902 343641
rect 115846 343567 115902 343576
rect 115846 342952 115902 342961
rect 115846 342887 115902 342896
rect 115756 342372 115808 342378
rect 115756 342314 115808 342320
rect 115768 335354 115796 342314
rect 115860 342310 115888 342887
rect 115848 342304 115900 342310
rect 115848 342246 115900 342252
rect 117226 337104 117282 337113
rect 117226 337039 117282 337048
rect 115768 335326 115888 335354
rect 115860 329474 115888 335326
rect 116768 334008 116820 334014
rect 116768 333950 116820 333956
rect 116780 329474 116808 333950
rect 117240 329746 117268 337039
rect 114572 329446 115000 329474
rect 115400 329446 115888 329474
rect 116472 329446 116808 329474
rect 117194 329718 117268 329746
rect 117194 329460 117222 329718
rect 118344 329474 118372 343703
rect 118620 332602 118648 364375
rect 119894 344312 119950 344321
rect 119894 344247 119950 344256
rect 118620 332574 119016 332602
rect 118884 332036 118936 332042
rect 118884 331978 118936 331984
rect 118896 329474 118924 331978
rect 117944 329446 118372 329474
rect 118680 329446 118924 329474
rect 118988 329474 119016 332574
rect 119908 332042 119936 344247
rect 119896 332036 119948 332042
rect 119896 331978 119948 331984
rect 120000 329882 120028 382230
rect 120264 365764 120316 365770
rect 120264 365706 120316 365712
rect 120276 345014 120304 365706
rect 121472 347818 121500 428431
rect 122116 401674 122144 556174
rect 122208 418033 122236 571338
rect 122286 444408 122342 444417
rect 122286 444343 122342 444352
rect 122194 418024 122250 418033
rect 122194 417959 122250 417968
rect 122104 401668 122156 401674
rect 122104 401610 122156 401616
rect 122300 355366 122328 444343
rect 122852 423745 122880 576098
rect 124220 550656 124272 550662
rect 124220 550598 124272 550604
rect 122932 463004 122984 463010
rect 122932 462946 122984 462952
rect 122838 423736 122894 423745
rect 122838 423671 122894 423680
rect 122840 413296 122892 413302
rect 122840 413238 122892 413244
rect 122852 412865 122880 413238
rect 122838 412856 122894 412865
rect 122838 412791 122894 412800
rect 122852 408626 122880 412791
rect 122760 408598 122880 408626
rect 122760 408354 122788 408598
rect 122760 408326 122880 408354
rect 122852 377466 122880 408326
rect 122944 403753 122972 462946
rect 123024 453348 123076 453354
rect 123024 453290 123076 453296
rect 123036 420918 123064 453290
rect 124126 444272 124182 444281
rect 124126 444207 124182 444216
rect 124140 443698 124168 444207
rect 124128 443692 124180 443698
rect 124128 443634 124180 443640
rect 124126 442096 124182 442105
rect 124126 442031 124182 442040
rect 124140 441658 124168 442031
rect 124128 441652 124180 441658
rect 124128 441594 124180 441600
rect 124126 437880 124182 437889
rect 124126 437815 124182 437824
rect 124140 437510 124168 437815
rect 124128 437504 124180 437510
rect 124128 437446 124180 437452
rect 124128 433288 124180 433294
rect 124126 433256 124128 433265
rect 124180 433256 124182 433265
rect 124126 433191 124182 433200
rect 124126 430672 124182 430681
rect 124126 430607 124128 430616
rect 124180 430607 124182 430616
rect 124128 430578 124180 430584
rect 123482 423736 123538 423745
rect 123482 423671 123538 423680
rect 123024 420912 123076 420918
rect 123024 420854 123076 420860
rect 123036 419665 123064 420854
rect 123022 419656 123078 419665
rect 123022 419591 123078 419600
rect 122930 403744 122986 403753
rect 122930 403679 122986 403688
rect 122944 403578 122972 403679
rect 122932 403572 122984 403578
rect 122932 403514 122984 403520
rect 122932 401668 122984 401674
rect 122932 401610 122984 401616
rect 122944 392601 122972 401610
rect 122930 392592 122986 392601
rect 122930 392527 122986 392536
rect 123496 387870 123524 423671
rect 124128 422272 124180 422278
rect 124128 422214 124180 422220
rect 124140 422113 124168 422214
rect 124126 422104 124182 422113
rect 124126 422039 124182 422048
rect 124126 415168 124182 415177
rect 124126 415103 124182 415112
rect 124140 414730 124168 415103
rect 124128 414724 124180 414730
rect 124128 414666 124180 414672
rect 124126 408504 124182 408513
rect 124126 408439 124128 408448
rect 124180 408439 124182 408448
rect 124128 408410 124180 408416
rect 123942 401568 123998 401577
rect 123942 401503 123998 401512
rect 123956 400926 123984 401503
rect 123944 400920 123996 400926
rect 123944 400862 123996 400868
rect 124126 399528 124182 399537
rect 124126 399463 124128 399472
rect 124180 399463 124182 399472
rect 124128 399434 124180 399440
rect 124128 396976 124180 396982
rect 124126 396944 124128 396953
rect 124180 396944 124182 396953
rect 124126 396879 124182 396888
rect 123758 392592 123814 392601
rect 123758 392527 123814 392536
rect 123772 392426 123800 392527
rect 123760 392420 123812 392426
rect 123760 392362 123812 392368
rect 123484 387864 123536 387870
rect 123484 387806 123536 387812
rect 122840 377460 122892 377466
rect 122840 377402 122892 377408
rect 123496 370569 123524 387806
rect 124232 386345 124260 550598
rect 124876 541006 124904 700266
rect 128360 584452 128412 584458
rect 128360 584394 128412 584400
rect 126886 546544 126942 546553
rect 126886 546479 126942 546488
rect 124864 541000 124916 541006
rect 124864 540942 124916 540948
rect 125600 455456 125652 455462
rect 125600 455398 125652 455404
rect 125508 453348 125560 453354
rect 125508 453290 125560 453296
rect 125520 452674 125548 453290
rect 125508 452668 125560 452674
rect 125508 452610 125560 452616
rect 124312 451988 124364 451994
rect 124312 451930 124364 451936
rect 124324 406337 124352 451930
rect 124310 406328 124366 406337
rect 124310 406263 124366 406272
rect 124324 406026 124352 406263
rect 124312 406020 124364 406026
rect 124312 405962 124364 405968
rect 124864 406020 124916 406026
rect 124864 405962 124916 405968
rect 124218 386336 124274 386345
rect 124218 386271 124274 386280
rect 123482 370560 123538 370569
rect 123482 370495 123538 370504
rect 124128 364404 124180 364410
rect 124128 364346 124180 364352
rect 123482 362400 123538 362409
rect 123482 362335 123538 362344
rect 122288 355360 122340 355366
rect 122288 355302 122340 355308
rect 121734 349752 121790 349761
rect 121734 349687 121790 349696
rect 121460 347812 121512 347818
rect 121460 347754 121512 347760
rect 121472 347041 121500 347754
rect 121458 347032 121514 347041
rect 121458 346967 121514 346976
rect 120722 346488 120778 346497
rect 120722 346423 120778 346432
rect 120276 344986 120488 345014
rect 120000 329854 120120 329882
rect 120092 329746 120120 329854
rect 120092 329718 120166 329746
rect 118988 329446 119416 329474
rect 120138 329460 120166 329718
rect 120460 329474 120488 344986
rect 120736 333305 120764 346423
rect 121748 345014 121776 349687
rect 123496 345098 123524 362335
rect 122840 345092 122892 345098
rect 122840 345034 122892 345040
rect 123484 345092 123536 345098
rect 123484 345034 123536 345040
rect 121748 344986 121960 345014
rect 120722 333296 120778 333305
rect 120722 333231 120778 333240
rect 121826 332752 121882 332761
rect 121826 332687 121882 332696
rect 121840 329474 121868 332687
rect 120460 329446 120888 329474
rect 121624 329446 121868 329474
rect 121932 329474 121960 344986
rect 122852 335354 122880 345034
rect 122852 335326 123432 335354
rect 123300 331492 123352 331498
rect 123300 331434 123352 331440
rect 123312 329474 123340 331434
rect 121932 329446 122360 329474
rect 123096 329446 123340 329474
rect 123404 329474 123432 335326
rect 124140 331498 124168 364346
rect 124876 353326 124904 405962
rect 125048 403572 125100 403578
rect 125048 403514 125100 403520
rect 124954 378720 125010 378729
rect 124954 378655 125010 378664
rect 124968 372706 124996 378655
rect 124956 372700 125008 372706
rect 124956 372642 125008 372648
rect 124864 353320 124916 353326
rect 124864 353262 124916 353268
rect 124862 347168 124918 347177
rect 124862 347103 124918 347112
rect 124218 335608 124274 335617
rect 124218 335543 124274 335552
rect 124232 333266 124260 335543
rect 124220 333260 124272 333266
rect 124220 333202 124272 333208
rect 124876 332897 124904 347103
rect 124968 335481 124996 372642
rect 125060 371210 125088 403514
rect 125520 395350 125548 452610
rect 125508 395344 125560 395350
rect 125508 395286 125560 395292
rect 125048 371204 125100 371210
rect 125048 371146 125100 371152
rect 125612 353258 125640 455398
rect 125692 447160 125744 447166
rect 125692 447102 125744 447108
rect 125704 399498 125732 447102
rect 125692 399492 125744 399498
rect 125692 399434 125744 399440
rect 126244 367872 126296 367878
rect 126244 367814 126296 367820
rect 125600 353252 125652 353258
rect 125600 353194 125652 353200
rect 125612 352578 125640 353194
rect 125600 352572 125652 352578
rect 125600 352514 125652 352520
rect 126256 348129 126284 367814
rect 126242 348120 126298 348129
rect 126242 348055 126298 348064
rect 125048 343664 125100 343670
rect 125048 343606 125100 343612
rect 124954 335472 125010 335481
rect 124954 335407 125010 335416
rect 124862 332888 124918 332897
rect 124862 332823 124918 332832
rect 124128 331492 124180 331498
rect 124128 331434 124180 331440
rect 124968 329474 124996 335407
rect 125060 335306 125088 343606
rect 125048 335300 125100 335306
rect 125048 335242 125100 335248
rect 125508 334076 125560 334082
rect 125508 334018 125560 334024
rect 125414 332888 125470 332897
rect 125414 332823 125470 332832
rect 125428 330041 125456 332823
rect 125520 330546 125548 334018
rect 125508 330540 125560 330546
rect 125508 330482 125560 330488
rect 125414 330032 125470 330041
rect 125414 329967 125470 329976
rect 123404 329446 123832 329474
rect 124568 329446 124996 329474
rect 103256 329174 103408 329202
rect 115400 329118 115428 329446
rect 125428 329202 125456 329967
rect 126256 329905 126284 348055
rect 126900 331294 126928 546479
rect 127624 477556 127676 477562
rect 127624 477498 127676 477504
rect 126980 457496 127032 457502
rect 126980 457438 127032 457444
rect 126992 443698 127020 457438
rect 127636 451246 127664 477498
rect 127716 456068 127768 456074
rect 127716 456010 127768 456016
rect 127624 451240 127676 451246
rect 127624 451182 127676 451188
rect 127624 444508 127676 444514
rect 127624 444450 127676 444456
rect 126980 443692 127032 443698
rect 126980 443634 127032 443640
rect 127636 359514 127664 444450
rect 127728 434042 127756 456010
rect 128372 437510 128400 584394
rect 129740 558952 129792 558958
rect 129740 558894 129792 558900
rect 129648 542428 129700 542434
rect 129648 542370 129700 542376
rect 129002 458280 129058 458289
rect 129002 458215 129058 458224
rect 129016 449886 129044 458215
rect 129004 449880 129056 449886
rect 129004 449822 129056 449828
rect 128360 437504 128412 437510
rect 128360 437446 128412 437452
rect 129004 437504 129056 437510
rect 129004 437446 129056 437452
rect 128360 434784 128412 434790
rect 128360 434726 128412 434732
rect 127716 434036 127768 434042
rect 127716 433978 127768 433984
rect 127728 433294 127756 433978
rect 127716 433288 127768 433294
rect 127716 433230 127768 433236
rect 126980 359508 127032 359514
rect 126980 359450 127032 359456
rect 127624 359508 127676 359514
rect 127624 359450 127676 359456
rect 126992 335354 127020 359450
rect 127072 353320 127124 353326
rect 127072 353262 127124 353268
rect 128176 353320 128228 353326
rect 128176 353262 128228 353268
rect 127084 345014 127112 353262
rect 128188 352073 128216 353262
rect 128174 352064 128230 352073
rect 128174 351999 128230 352008
rect 128372 349897 128400 434726
rect 129016 370569 129044 437446
rect 129660 376825 129688 542370
rect 129752 396982 129780 558894
rect 130396 536790 130424 702782
rect 137848 700330 137876 703520
rect 154132 702545 154160 703520
rect 170324 702982 170352 703520
rect 169760 702976 169812 702982
rect 169760 702918 169812 702924
rect 170312 702976 170364 702982
rect 170312 702918 170364 702924
rect 169772 702710 169800 702918
rect 202800 702914 202828 703520
rect 202788 702908 202840 702914
rect 202788 702850 202840 702856
rect 218992 702846 219020 703520
rect 218980 702840 219032 702846
rect 218980 702782 219032 702788
rect 233884 702772 233936 702778
rect 233884 702714 233936 702720
rect 169760 702704 169812 702710
rect 169760 702646 169812 702652
rect 197268 702704 197320 702710
rect 197268 702646 197320 702652
rect 154118 702536 154174 702545
rect 154118 702471 154174 702480
rect 137836 700324 137888 700330
rect 137836 700266 137888 700272
rect 155224 594856 155276 594862
rect 155224 594798 155276 594804
rect 155236 576854 155264 594798
rect 155236 576826 155356 576854
rect 136640 574116 136692 574122
rect 136640 574058 136692 574064
rect 133144 567248 133196 567254
rect 133144 567190 133196 567196
rect 133156 560250 133184 567190
rect 133880 565140 133932 565146
rect 133880 565082 133932 565088
rect 135168 565140 135220 565146
rect 135168 565082 135220 565088
rect 133144 560244 133196 560250
rect 133144 560186 133196 560192
rect 133788 560244 133840 560250
rect 133788 560186 133840 560192
rect 133800 559026 133828 560186
rect 133788 559020 133840 559026
rect 133788 558962 133840 558968
rect 130474 536888 130530 536897
rect 130474 536823 130530 536832
rect 130384 536784 130436 536790
rect 130384 536726 130436 536732
rect 130488 447001 130516 536823
rect 132500 532092 132552 532098
rect 132500 532034 132552 532040
rect 133696 532092 133748 532098
rect 133696 532034 133748 532040
rect 132408 480276 132460 480282
rect 132408 480218 132460 480224
rect 130568 465112 130620 465118
rect 130568 465054 130620 465060
rect 130474 446992 130530 447001
rect 130474 446927 130530 446936
rect 130382 444408 130438 444417
rect 130382 444343 130438 444352
rect 130396 409834 130424 444343
rect 130580 440230 130608 465054
rect 130568 440224 130620 440230
rect 130568 440166 130620 440172
rect 130384 409828 130436 409834
rect 130384 409770 130436 409776
rect 129740 396976 129792 396982
rect 129740 396918 129792 396924
rect 129752 393990 129780 396918
rect 129740 393984 129792 393990
rect 129740 393926 129792 393932
rect 131764 392420 131816 392426
rect 131764 392362 131816 392368
rect 130384 392012 130436 392018
rect 130384 391954 130436 391960
rect 129832 379636 129884 379642
rect 129832 379578 129884 379584
rect 129094 376816 129150 376825
rect 129094 376751 129150 376760
rect 129646 376816 129702 376825
rect 129646 376751 129702 376760
rect 129002 370560 129058 370569
rect 129002 370495 129058 370504
rect 128358 349888 128414 349897
rect 128358 349823 128414 349832
rect 127084 344986 127848 345014
rect 126992 335326 127112 335354
rect 126888 331288 126940 331294
rect 126888 331230 126940 331236
rect 126242 329896 126298 329905
rect 126242 329831 126298 329840
rect 126256 329474 126284 329831
rect 126900 329474 126928 331230
rect 126040 329446 126284 329474
rect 126776 329446 126928 329474
rect 127084 329474 127112 335326
rect 127820 329474 127848 344986
rect 129108 331906 129136 376751
rect 129740 371204 129792 371210
rect 129740 371146 129792 371152
rect 129188 369912 129240 369918
rect 129188 369854 129240 369860
rect 129200 334665 129228 369854
rect 129752 369073 129780 371146
rect 129738 369064 129794 369073
rect 129738 368999 129794 369008
rect 129844 345014 129872 379578
rect 130396 374746 130424 391954
rect 131120 390584 131172 390590
rect 131120 390526 131172 390532
rect 131132 389230 131160 390526
rect 131120 389224 131172 389230
rect 131120 389166 131172 389172
rect 130384 374740 130436 374746
rect 130384 374682 130436 374688
rect 131776 374066 131804 392362
rect 132420 390590 132448 480218
rect 132408 390584 132460 390590
rect 132408 390526 132460 390532
rect 132512 377913 132540 532034
rect 133708 531350 133736 532034
rect 133696 531344 133748 531350
rect 133696 531286 133748 531292
rect 132592 454096 132644 454102
rect 132592 454038 132644 454044
rect 132498 377904 132554 377913
rect 132498 377839 132554 377848
rect 131764 374060 131816 374066
rect 131764 374002 131816 374008
rect 131776 369850 131804 374002
rect 131764 369844 131816 369850
rect 131764 369786 131816 369792
rect 132512 369730 132540 377839
rect 132420 369702 132540 369730
rect 132420 369209 132448 369702
rect 132406 369200 132462 369209
rect 132406 369135 132462 369144
rect 131028 362228 131080 362234
rect 131028 362170 131080 362176
rect 131040 357490 131068 362170
rect 131040 357474 131160 357490
rect 130384 357468 130436 357474
rect 131040 357468 131172 357474
rect 131040 357462 131120 357468
rect 130384 357410 130436 357416
rect 131120 357410 131172 357416
rect 129844 344986 130056 345014
rect 129186 334656 129242 334665
rect 129186 334591 129242 334600
rect 129280 331968 129332 331974
rect 129280 331910 129332 331916
rect 129096 331900 129148 331906
rect 129096 331842 129148 331848
rect 129292 329474 129320 331910
rect 129924 331492 129976 331498
rect 129924 331434 129976 331440
rect 129740 331288 129792 331294
rect 129740 331230 129792 331236
rect 129752 331129 129780 331230
rect 129738 331120 129794 331129
rect 129738 331055 129794 331064
rect 129936 329474 129964 331434
rect 127084 329446 127512 329474
rect 127820 329446 128248 329474
rect 128984 329446 129320 329474
rect 129720 329446 129964 329474
rect 130028 329474 130056 344986
rect 130396 331498 130424 357410
rect 132420 331498 132448 369135
rect 132604 349858 132632 454038
rect 133800 408474 133828 558962
rect 133892 413302 133920 565082
rect 135180 564466 135208 565082
rect 135168 564460 135220 564466
rect 135168 564402 135220 564408
rect 135260 534744 135312 534750
rect 135260 534686 135312 534692
rect 136180 534744 136232 534750
rect 136180 534686 136232 534692
rect 134524 507136 134576 507142
rect 134524 507078 134576 507084
rect 133880 413296 133932 413302
rect 133880 413238 133932 413244
rect 133788 408468 133840 408474
rect 133788 408410 133840 408416
rect 133144 405748 133196 405754
rect 133144 405690 133196 405696
rect 133156 370705 133184 405690
rect 134536 385665 134564 507078
rect 134616 408468 134668 408474
rect 134616 408410 134668 408416
rect 134522 385656 134578 385665
rect 134522 385591 134578 385600
rect 133142 370696 133198 370705
rect 133142 370631 133198 370640
rect 133880 363656 133932 363662
rect 133880 363598 133932 363604
rect 133786 360496 133842 360505
rect 133786 360431 133842 360440
rect 133144 353320 133196 353326
rect 133144 353262 133196 353268
rect 132592 349852 132644 349858
rect 132592 349794 132644 349800
rect 133156 340202 133184 353262
rect 133694 347848 133750 347857
rect 133694 347783 133750 347792
rect 133144 340196 133196 340202
rect 133144 340138 133196 340144
rect 133708 331498 133736 347783
rect 130384 331492 130436 331498
rect 130384 331434 130436 331440
rect 131488 331492 131540 331498
rect 131488 331434 131540 331440
rect 132408 331492 132460 331498
rect 132408 331434 132460 331440
rect 132776 331492 132828 331498
rect 132776 331434 132828 331440
rect 133696 331492 133748 331498
rect 133696 331434 133748 331440
rect 131500 329474 131528 331434
rect 132788 329474 132816 331434
rect 133800 329474 133828 360431
rect 133892 329746 133920 363598
rect 134628 339697 134656 408410
rect 135272 388793 135300 534686
rect 136192 534138 136220 534686
rect 136180 534132 136232 534138
rect 136180 534074 136232 534080
rect 136652 422278 136680 574058
rect 138020 566500 138072 566506
rect 138020 566442 138072 566448
rect 138032 565894 138060 566442
rect 138020 565888 138072 565894
rect 138020 565830 138072 565836
rect 137928 545148 137980 545154
rect 137928 545090 137980 545096
rect 137284 426488 137336 426494
rect 137284 426430 137336 426436
rect 136640 422272 136692 422278
rect 136640 422214 136692 422220
rect 136652 421598 136680 422214
rect 136640 421592 136692 421598
rect 136640 421534 136692 421540
rect 135258 388784 135314 388793
rect 135258 388719 135314 388728
rect 136638 378176 136694 378185
rect 136638 378111 136694 378120
rect 136548 361616 136600 361622
rect 136548 361558 136600 361564
rect 134614 339688 134670 339697
rect 134614 339623 134670 339632
rect 134248 339584 134300 339590
rect 134248 339526 134300 339532
rect 133892 329718 133966 329746
rect 130028 329446 130456 329474
rect 131192 329446 131528 329474
rect 132480 329446 132816 329474
rect 133216 329446 133828 329474
rect 133938 329460 133966 329718
rect 134260 329474 134288 339526
rect 135720 331492 135772 331498
rect 135720 331434 135772 331440
rect 135732 329474 135760 331434
rect 136560 331226 136588 361558
rect 136652 345014 136680 378111
rect 137296 349110 137324 426430
rect 137940 378185 137968 545090
rect 138032 414730 138060 565830
rect 148416 556844 148468 556850
rect 148416 556786 148468 556792
rect 142066 542600 142122 542609
rect 142066 542535 142122 542544
rect 141422 444680 141478 444689
rect 141422 444615 141478 444624
rect 140044 441652 140096 441658
rect 140044 441594 140096 441600
rect 138020 414724 138072 414730
rect 138020 414666 138072 414672
rect 137926 378176 137982 378185
rect 137926 378111 137982 378120
rect 138032 351218 138060 414666
rect 140056 396778 140084 441594
rect 140044 396772 140096 396778
rect 140044 396714 140096 396720
rect 139306 355464 139362 355473
rect 139306 355399 139362 355408
rect 138020 351212 138072 351218
rect 138020 351154 138072 351160
rect 138032 351121 138060 351154
rect 138018 351112 138074 351121
rect 138018 351047 138074 351056
rect 137284 349104 137336 349110
rect 137284 349046 137336 349052
rect 136652 344986 137232 345014
rect 136548 331220 136600 331226
rect 136548 331162 136600 331168
rect 136454 329896 136510 329905
rect 136560 329882 136588 331162
rect 136560 329854 136680 329882
rect 136454 329831 136510 329840
rect 136468 329474 136496 329831
rect 134260 329446 134688 329474
rect 135424 329446 135760 329474
rect 136160 329446 136496 329474
rect 136652 329474 136680 329854
rect 137204 329474 137232 344986
rect 137284 343664 137336 343670
rect 137284 343606 137336 343612
rect 137296 336161 137324 343606
rect 137282 336152 137338 336161
rect 137282 336087 137338 336096
rect 139214 335472 139270 335481
rect 139214 335407 139270 335416
rect 138664 331356 138716 331362
rect 138664 331298 138716 331304
rect 138676 329474 138704 331298
rect 139228 329474 139256 335407
rect 139320 331362 139348 355399
rect 140688 348424 140740 348430
rect 140688 348366 140740 348372
rect 139398 339688 139454 339697
rect 139398 339623 139454 339632
rect 139308 331356 139360 331362
rect 139308 331298 139360 331304
rect 136652 329446 136896 329474
rect 137204 329446 137632 329474
rect 138368 329446 138704 329474
rect 139104 329446 139256 329474
rect 139412 329474 139440 339623
rect 140700 329474 140728 348366
rect 141436 346633 141464 444615
rect 141516 356108 141568 356114
rect 141516 356050 141568 356056
rect 140778 346624 140834 346633
rect 140778 346559 140834 346568
rect 141422 346624 141478 346633
rect 141422 346559 141478 346568
rect 140792 345014 140820 346559
rect 140792 344986 140912 345014
rect 140780 332648 140832 332654
rect 140780 332590 140832 332596
rect 140792 331906 140820 332590
rect 140780 331900 140832 331906
rect 140780 331842 140832 331848
rect 139412 329446 139840 329474
rect 140576 329446 140728 329474
rect 140884 329474 140912 344986
rect 141528 341562 141556 356050
rect 141516 341556 141568 341562
rect 141516 341498 141568 341504
rect 142080 341057 142108 542535
rect 146944 535492 146996 535498
rect 146944 535434 146996 535440
rect 143448 534132 143500 534138
rect 143448 534074 143500 534080
rect 143460 532710 143488 534074
rect 143448 532704 143500 532710
rect 143448 532646 143500 532652
rect 144184 531344 144236 531350
rect 144184 531286 144236 531292
rect 144196 500954 144224 531286
rect 144184 500948 144236 500954
rect 144184 500890 144236 500896
rect 145564 474768 145616 474774
rect 145564 474710 145616 474716
rect 142804 473408 142856 473414
rect 142804 473350 142856 473356
rect 142816 391241 142844 473350
rect 145576 391270 145604 474710
rect 146956 447098 146984 535434
rect 148324 492720 148376 492726
rect 148324 492662 148376 492668
rect 146944 447092 146996 447098
rect 146944 447034 146996 447040
rect 146944 444440 146996 444446
rect 146944 444382 146996 444388
rect 145564 391264 145616 391270
rect 142802 391232 142858 391241
rect 145564 391206 145616 391212
rect 142802 391167 142858 391176
rect 146208 370592 146260 370598
rect 146208 370534 146260 370540
rect 144828 368552 144880 368558
rect 144828 368494 144880 368500
rect 144734 363216 144790 363225
rect 144734 363151 144790 363160
rect 144184 342304 144236 342310
rect 144184 342246 144236 342252
rect 141422 341048 141478 341057
rect 141422 340983 141478 340992
rect 142066 341048 142122 341057
rect 142066 340983 142122 340992
rect 142344 341012 142396 341018
rect 141436 331498 141464 340983
rect 142344 340954 142396 340960
rect 142066 331936 142122 331945
rect 142066 331871 142122 331880
rect 141424 331492 141476 331498
rect 141424 331434 141476 331440
rect 142080 329746 142108 331871
rect 142034 329718 142108 329746
rect 140884 329446 141312 329474
rect 142034 329460 142062 329718
rect 142356 329474 142384 340954
rect 144196 335306 144224 342246
rect 144748 335354 144776 363151
rect 144656 335326 144776 335354
rect 144184 335300 144236 335306
rect 144184 335242 144236 335248
rect 143816 331356 143868 331362
rect 143816 331298 143868 331304
rect 143828 329474 143856 331298
rect 144656 329474 144684 335326
rect 144840 331362 144868 368494
rect 146220 335354 146248 370534
rect 146956 351150 146984 444382
rect 148336 382974 148364 492662
rect 148428 487830 148456 556786
rect 155328 556238 155356 576826
rect 174544 569968 174596 569974
rect 174544 569910 174596 569916
rect 155868 567248 155920 567254
rect 155868 567190 155920 567196
rect 155316 556232 155368 556238
rect 155316 556174 155368 556180
rect 154764 537532 154816 537538
rect 154764 537474 154816 537480
rect 151084 534744 151136 534750
rect 151084 534686 151136 534692
rect 148416 487824 148468 487830
rect 148416 487766 148468 487772
rect 151096 453354 151124 534686
rect 153108 530596 153160 530602
rect 153108 530538 153160 530544
rect 151084 453348 151136 453354
rect 151084 453290 151136 453296
rect 151084 409896 151136 409902
rect 151084 409838 151136 409844
rect 148416 395344 148468 395350
rect 148416 395286 148468 395292
rect 148324 382968 148376 382974
rect 148324 382910 148376 382916
rect 147680 382356 147732 382362
rect 147680 382298 147732 382304
rect 146944 351144 146996 351150
rect 146944 351086 146996 351092
rect 147588 351144 147640 351150
rect 147588 351086 147640 351092
rect 146128 335326 146248 335354
rect 145288 334076 145340 334082
rect 145288 334018 145340 334024
rect 145300 331974 145328 334018
rect 145288 331968 145340 331974
rect 145288 331910 145340 331916
rect 144828 331356 144880 331362
rect 144828 331298 144880 331304
rect 145286 330440 145342 330449
rect 145286 330375 145342 330384
rect 145300 329474 145328 330375
rect 145378 329896 145434 329905
rect 145378 329831 145434 329840
rect 142356 329446 142784 329474
rect 143520 329446 143856 329474
rect 144256 329446 144684 329474
rect 144992 329446 145328 329474
rect 125304 329174 125456 329202
rect 145392 329118 145420 329831
rect 146128 329474 146156 335326
rect 146206 334248 146262 334257
rect 146206 334183 146262 334192
rect 146220 331945 146248 334183
rect 146206 331936 146262 331945
rect 146206 331871 146262 331880
rect 146760 331288 146812 331294
rect 146760 331230 146812 331236
rect 146772 329474 146800 331230
rect 147600 329474 147628 351086
rect 145728 329446 146156 329474
rect 146464 329446 146800 329474
rect 147200 329446 147628 329474
rect 147692 329474 147720 382298
rect 148428 368354 148456 395286
rect 147772 368348 147824 368354
rect 147772 368290 147824 368296
rect 148416 368348 148468 368354
rect 148416 368290 148468 368296
rect 147784 367130 147812 368290
rect 147772 367124 147824 367130
rect 147772 367066 147824 367072
rect 147784 345014 147812 367066
rect 151096 362409 151124 409838
rect 152464 380180 152516 380186
rect 152464 380122 152516 380128
rect 151082 362400 151138 362409
rect 151082 362335 151138 362344
rect 150346 359544 150402 359553
rect 150346 359479 150402 359488
rect 149058 346488 149114 346497
rect 149058 346423 149114 346432
rect 149072 345681 149100 346423
rect 149058 345672 149114 345681
rect 149058 345607 149114 345616
rect 147784 344986 148272 345014
rect 148244 329474 148272 344986
rect 150360 335354 150388 359479
rect 151082 356144 151138 356153
rect 151082 356079 151138 356088
rect 151096 347818 151124 356079
rect 151084 347812 151136 347818
rect 151084 347754 151136 347760
rect 150440 346520 150492 346526
rect 150440 346462 150492 346468
rect 150452 345030 150480 346462
rect 150440 345024 150492 345030
rect 150440 344966 150492 344972
rect 151096 338094 151124 347754
rect 151726 346488 151782 346497
rect 151726 346423 151782 346432
rect 151084 338088 151136 338094
rect 151084 338030 151136 338036
rect 150530 337240 150586 337249
rect 150530 337175 150586 337184
rect 150438 336968 150494 336977
rect 150438 336903 150494 336912
rect 150452 336025 150480 336903
rect 150544 336054 150572 337175
rect 150532 336048 150584 336054
rect 150438 336016 150494 336025
rect 150532 335990 150584 335996
rect 150438 335951 150494 335960
rect 150440 335436 150492 335442
rect 150440 335378 150492 335384
rect 150268 335326 150388 335354
rect 150268 331265 150296 335326
rect 150452 334529 150480 335378
rect 150438 334520 150494 334529
rect 150438 334455 150494 334464
rect 150438 334112 150494 334121
rect 150438 334047 150494 334056
rect 150452 333266 150480 334047
rect 150440 333260 150492 333266
rect 150440 333202 150492 333208
rect 150348 332648 150400 332654
rect 150348 332590 150400 332596
rect 149702 331256 149758 331265
rect 149702 331191 149758 331200
rect 150254 331256 150310 331265
rect 150254 331191 150310 331200
rect 149716 329474 149744 331191
rect 150360 329474 150388 332590
rect 151176 329860 151228 329866
rect 151176 329802 151228 329808
rect 151188 329474 151216 329802
rect 151740 329474 151768 346423
rect 151910 335744 151966 335753
rect 151910 335679 151966 335688
rect 151924 331809 151952 335679
rect 152476 332489 152504 380122
rect 152648 338088 152700 338094
rect 152648 338030 152700 338036
rect 152462 332480 152518 332489
rect 152462 332415 152518 332424
rect 151910 331800 151966 331809
rect 151910 331735 151966 331744
rect 147692 329446 147936 329474
rect 148244 329446 148672 329474
rect 149408 329446 149744 329474
rect 150144 329446 150388 329474
rect 150880 329446 151216 329474
rect 151616 329446 151768 329474
rect 152660 329474 152688 338030
rect 153120 335753 153148 530538
rect 154776 529854 154804 537474
rect 154764 529848 154816 529854
rect 154764 529790 154816 529796
rect 155224 521688 155276 521694
rect 155224 521630 155276 521636
rect 155236 383081 155264 521630
rect 155328 448633 155356 556174
rect 155314 448624 155370 448633
rect 155314 448559 155370 448568
rect 155328 436082 155356 448559
rect 155776 437436 155828 437442
rect 155776 437378 155828 437384
rect 155316 436076 155368 436082
rect 155316 436018 155368 436024
rect 155222 383072 155278 383081
rect 155222 383007 155278 383016
rect 153844 376780 153896 376786
rect 153844 376722 153896 376728
rect 153856 367810 153884 376722
rect 155224 369164 155276 369170
rect 155224 369106 155276 369112
rect 153844 367804 153896 367810
rect 153844 367746 153896 367752
rect 155236 356833 155264 369106
rect 155222 356824 155278 356833
rect 155222 356759 155278 356768
rect 153842 347984 153898 347993
rect 153842 347919 153898 347928
rect 153856 341562 153884 347919
rect 155222 345672 155278 345681
rect 155222 345607 155278 345616
rect 153844 341556 153896 341562
rect 153844 341498 153896 341504
rect 154028 341012 154080 341018
rect 154028 340954 154080 340960
rect 153842 338600 153898 338609
rect 153842 338535 153898 338544
rect 153198 337104 153254 337113
rect 153198 337039 153254 337048
rect 153106 335744 153162 335753
rect 153106 335679 153162 335688
rect 153212 334665 153240 337039
rect 153198 334656 153254 334665
rect 153198 334591 153254 334600
rect 153106 332888 153162 332897
rect 153106 332823 153162 332832
rect 153120 331945 153148 332823
rect 153106 331936 153162 331945
rect 153106 331871 153162 331880
rect 153198 331120 153254 331129
rect 153198 331055 153254 331064
rect 153212 330614 153240 331055
rect 153200 330608 153252 330614
rect 153856 330585 153884 338535
rect 154040 338065 154068 340954
rect 154486 338464 154542 338473
rect 154486 338399 154542 338408
rect 154500 338230 154528 338399
rect 154488 338224 154540 338230
rect 154488 338166 154540 338172
rect 154026 338056 154082 338065
rect 154026 337991 154082 338000
rect 155236 333305 155264 345607
rect 155316 338224 155368 338230
rect 155316 338166 155368 338172
rect 155222 333296 155278 333305
rect 155222 333231 155278 333240
rect 155328 332489 155356 338166
rect 155314 332480 155370 332489
rect 155314 332415 155370 332424
rect 154854 331800 154910 331809
rect 154854 331735 154910 331744
rect 153200 330550 153252 330556
rect 153842 330576 153898 330585
rect 153842 330511 153898 330520
rect 153200 330472 153252 330478
rect 153200 330414 153252 330420
rect 153212 329798 153240 330414
rect 154118 330032 154174 330041
rect 154118 329967 154174 329976
rect 153200 329792 153252 329798
rect 153200 329734 153252 329740
rect 154132 329474 154160 329967
rect 154868 329474 154896 331735
rect 155328 329746 155356 332415
rect 155788 331809 155816 437378
rect 155774 331800 155830 331809
rect 155774 331735 155830 331744
rect 155788 331401 155816 331735
rect 155774 331392 155830 331401
rect 155774 331327 155830 331336
rect 152660 329446 153088 329474
rect 153824 329446 154160 329474
rect 154560 329446 154896 329474
rect 155282 329718 155356 329746
rect 155282 329460 155310 329718
rect 155880 329118 155908 567190
rect 169114 552120 169170 552129
rect 169114 552055 169170 552064
rect 169128 539481 169156 552055
rect 169114 539472 169170 539481
rect 169114 539407 169170 539416
rect 171784 538960 171836 538966
rect 171784 538902 171836 538908
rect 169024 538892 169076 538898
rect 169024 538834 169076 538840
rect 162216 525836 162268 525842
rect 162216 525778 162268 525784
rect 162124 516180 162176 516186
rect 162124 516122 162176 516128
rect 156604 465724 156656 465730
rect 156604 465666 156656 465672
rect 156616 465225 156644 465666
rect 156602 465216 156658 465225
rect 156602 465151 156658 465160
rect 156616 465118 156644 465151
rect 156604 465112 156656 465118
rect 156604 465054 156656 465060
rect 159364 459604 159416 459610
rect 159364 459546 159416 459552
rect 157984 456816 158036 456822
rect 157984 456758 158036 456764
rect 156604 436076 156656 436082
rect 156604 436018 156656 436024
rect 156616 343913 156644 436018
rect 157996 382974 158024 456758
rect 158074 387016 158130 387025
rect 158074 386951 158130 386960
rect 157984 382968 158036 382974
rect 157984 382910 158036 382916
rect 157340 382356 157392 382362
rect 157340 382298 157392 382304
rect 157352 381002 157380 382298
rect 157984 381540 158036 381546
rect 157984 381482 158036 381488
rect 157340 380996 157392 381002
rect 157340 380938 157392 380944
rect 157340 350600 157392 350606
rect 157340 350542 157392 350548
rect 157352 346390 157380 350542
rect 157340 346384 157392 346390
rect 157340 346326 157392 346332
rect 156602 343904 156658 343913
rect 156602 343839 156658 343848
rect 156878 343768 156934 343777
rect 156878 343703 156934 343712
rect 156788 343664 156840 343670
rect 156788 343606 156840 343612
rect 155960 330608 156012 330614
rect 155960 330550 156012 330556
rect 155972 329905 156000 330550
rect 155958 329896 156014 329905
rect 155958 329831 156014 329840
rect 94228 329112 94280 329118
rect 94228 329054 94280 329060
rect 115388 329112 115440 329118
rect 132224 329112 132276 329118
rect 115388 329054 115440 329060
rect 131928 329060 132224 329066
rect 131928 329054 132276 329060
rect 145380 329112 145432 329118
rect 145380 329054 145432 329060
rect 152188 329112 152240 329118
rect 155868 329112 155920 329118
rect 152240 329060 152352 329066
rect 152188 329054 152352 329060
rect 156328 329112 156380 329118
rect 155868 329054 155920 329060
rect 156032 329060 156328 329066
rect 156032 329054 156380 329060
rect 131928 329038 132264 329054
rect 152200 329038 152352 329054
rect 156032 329038 156368 329054
rect 156584 328902 156736 328930
rect 156708 328506 156736 328902
rect 156696 328500 156748 328506
rect 156696 328442 156748 328448
rect 156696 328296 156748 328302
rect 156696 328238 156748 328244
rect 156708 327146 156736 328238
rect 156696 327140 156748 327146
rect 156696 327082 156748 327088
rect 67822 323504 67878 323513
rect 67822 323439 67878 323448
rect 156800 318102 156828 343606
rect 156892 329769 156920 343703
rect 157996 343670 158024 381482
rect 158088 351898 158116 386951
rect 158076 351892 158128 351898
rect 158076 351834 158128 351840
rect 158628 351892 158680 351898
rect 158628 351834 158680 351840
rect 158076 345704 158128 345710
rect 158076 345646 158128 345652
rect 157984 343664 158036 343670
rect 157984 343606 158036 343612
rect 157338 341048 157394 341057
rect 157338 340983 157394 340992
rect 157352 337385 157380 340983
rect 157982 338056 158038 338065
rect 157982 337991 158038 338000
rect 157338 337376 157394 337385
rect 157338 337311 157394 337320
rect 157996 333441 158024 337991
rect 157982 333432 158038 333441
rect 157982 333367 158038 333376
rect 157340 331900 157392 331906
rect 157340 331842 157392 331848
rect 157352 330614 157380 331842
rect 157340 330608 157392 330614
rect 157340 330550 157392 330556
rect 157984 329860 158036 329866
rect 157984 329802 158036 329808
rect 156878 329760 156934 329769
rect 156878 329695 156934 329704
rect 157064 329112 157116 329118
rect 157064 329054 157116 329060
rect 156880 328636 156932 328642
rect 156880 328578 156932 328584
rect 156892 328545 156920 328578
rect 156878 328536 156934 328545
rect 156878 328471 156934 328480
rect 156880 328364 156932 328370
rect 156880 328306 156932 328312
rect 156892 327729 156920 328306
rect 156878 327720 156934 327729
rect 156878 327655 156934 327664
rect 157076 326398 157104 329054
rect 157064 326392 157116 326398
rect 157064 326334 157116 326340
rect 156788 318096 156840 318102
rect 156788 318038 156840 318044
rect 67730 308544 67786 308553
rect 67730 308479 67786 308488
rect 67638 304192 67694 304201
rect 67638 304127 67694 304136
rect 67546 299840 67602 299849
rect 67546 299775 67602 299784
rect 67638 295488 67694 295497
rect 67638 295423 67694 295432
rect 67454 291136 67510 291145
rect 67454 291071 67510 291080
rect 67362 287872 67418 287881
rect 67362 287807 67364 287816
rect 67416 287807 67418 287816
rect 67364 287778 67416 287784
rect 67376 287747 67404 287778
rect 67362 281344 67418 281353
rect 67362 281279 67418 281288
rect 66994 274000 67050 274009
rect 66994 273935 67050 273944
rect 66904 271176 66956 271182
rect 66904 271118 66956 271124
rect 66902 270736 66958 270745
rect 66902 270671 66958 270680
rect 66916 270570 66944 270671
rect 66904 270564 66956 270570
rect 66904 270506 66956 270512
rect 66810 268560 66866 268569
rect 66810 268495 66866 268504
rect 66824 267918 66852 268495
rect 66812 267912 66864 267918
rect 66812 267854 66864 267860
rect 66810 265296 66866 265305
rect 66810 265231 66866 265240
rect 66824 264994 66852 265231
rect 66812 264988 66864 264994
rect 66812 264930 66864 264936
rect 66902 264208 66958 264217
rect 66902 264143 66958 264152
rect 66916 263634 66944 264143
rect 66904 263628 66956 263634
rect 66904 263570 66956 263576
rect 66810 263120 66866 263129
rect 66810 263055 66866 263064
rect 66824 262274 66852 263055
rect 66812 262268 66864 262274
rect 66812 262210 66864 262216
rect 66258 262032 66314 262041
rect 66258 261967 66314 261976
rect 66272 260914 66300 261967
rect 66812 260976 66864 260982
rect 66810 260944 66812 260953
rect 66864 260944 66866 260953
rect 66260 260908 66312 260914
rect 66810 260879 66866 260888
rect 66260 260850 66312 260856
rect 66260 258120 66312 258126
rect 66258 258088 66260 258097
rect 66312 258088 66314 258097
rect 66258 258023 66314 258032
rect 66902 257680 66958 257689
rect 66902 257615 66958 257624
rect 66916 256766 66944 257615
rect 66904 256760 66956 256766
rect 66904 256702 66956 256708
rect 66810 255504 66866 255513
rect 66810 255439 66866 255448
rect 66824 255338 66852 255439
rect 66812 255332 66864 255338
rect 66812 255274 66864 255280
rect 66810 254416 66866 254425
rect 66810 254351 66866 254360
rect 66824 253978 66852 254351
rect 66812 253972 66864 253978
rect 66812 253914 66864 253920
rect 66810 253328 66866 253337
rect 66810 253263 66866 253272
rect 66824 252618 66852 253263
rect 66812 252612 66864 252618
rect 66812 252554 66864 252560
rect 67008 251802 67036 273935
rect 66996 251796 67048 251802
rect 66996 251738 67048 251744
rect 67178 248976 67234 248985
rect 67178 248911 67234 248920
rect 66812 247036 66864 247042
rect 66812 246978 66864 246984
rect 66824 246809 66852 246978
rect 66810 246800 66866 246809
rect 66810 246735 66866 246744
rect 66810 245712 66866 245721
rect 66810 245647 66812 245656
rect 66864 245647 66866 245656
rect 66812 245618 66864 245624
rect 66904 245608 66956 245614
rect 66904 245550 66956 245556
rect 66916 244633 66944 245550
rect 66902 244624 66958 244633
rect 66902 244559 66958 244568
rect 67088 244452 67140 244458
rect 67088 244394 67140 244400
rect 67100 241398 67128 244394
rect 67088 241392 67140 241398
rect 67088 241334 67140 241340
rect 66074 226944 66130 226953
rect 66074 226879 66130 226888
rect 64788 197328 64840 197334
rect 64788 197270 64840 197276
rect 66166 129296 66222 129305
rect 66166 129231 66222 129240
rect 66180 128382 66208 129231
rect 66168 128376 66220 128382
rect 66168 128318 66220 128324
rect 66166 128072 66222 128081
rect 66166 128007 66222 128016
rect 66180 127129 66208 128007
rect 64786 127120 64842 127129
rect 64786 127055 64842 127064
rect 66166 127120 66222 127129
rect 66166 127055 66222 127064
rect 64694 121544 64750 121553
rect 64694 121479 64750 121488
rect 64708 89010 64736 121479
rect 64800 93158 64828 127055
rect 66166 126304 66222 126313
rect 66166 126239 66222 126248
rect 66074 122632 66130 122641
rect 66074 122567 66130 122576
rect 66088 121553 66116 122567
rect 66074 121544 66130 121553
rect 66074 121479 66130 121488
rect 66074 120864 66130 120873
rect 66074 120799 66130 120808
rect 66088 94518 66116 120799
rect 66076 94512 66128 94518
rect 66180 94489 66208 126239
rect 66076 94454 66128 94460
rect 66166 94480 66222 94489
rect 66166 94415 66222 94424
rect 64788 93152 64840 93158
rect 64788 93094 64840 93100
rect 64696 89004 64748 89010
rect 64696 88946 64748 88952
rect 66166 48920 66222 48929
rect 66166 48855 66222 48864
rect 64786 44840 64842 44849
rect 64786 44775 64842 44784
rect 62028 32428 62080 32434
rect 62028 32370 62080 32376
rect 62028 6180 62080 6186
rect 62028 6122 62080 6128
rect 60832 3528 60884 3534
rect 60832 3470 60884 3476
rect 61936 3528 61988 3534
rect 61936 3470 61988 3476
rect 60004 2168 60056 2174
rect 60004 2110 60056 2116
rect 60844 480 60872 3470
rect 62040 480 62068 6122
rect 64800 3602 64828 44775
rect 64328 3596 64380 3602
rect 64328 3538 64380 3544
rect 64788 3596 64840 3602
rect 64788 3538 64840 3544
rect 63224 3528 63276 3534
rect 63224 3470 63276 3476
rect 63236 480 63264 3470
rect 64340 480 64368 3538
rect 66180 3534 66208 48855
rect 67192 22846 67220 248911
rect 67376 244458 67404 281279
rect 67364 244452 67416 244458
rect 67364 244394 67416 244400
rect 67468 244338 67496 291071
rect 67546 280256 67602 280265
rect 67546 280191 67548 280200
rect 67600 280191 67602 280200
rect 67548 280162 67600 280168
rect 67546 251152 67602 251161
rect 67546 251087 67602 251096
rect 67560 248470 67588 251087
rect 67548 248464 67600 248470
rect 67548 248406 67600 248412
rect 67548 248328 67600 248334
rect 67548 248270 67600 248276
rect 67376 244310 67496 244338
rect 67270 243536 67326 243545
rect 67270 243471 67326 243480
rect 67284 222873 67312 243471
rect 67376 240038 67404 244310
rect 67456 244248 67508 244254
rect 67456 244190 67508 244196
rect 67468 243545 67496 244190
rect 67454 243536 67510 243545
rect 67454 243471 67510 243480
rect 67560 243409 67588 248270
rect 67546 243400 67602 243409
rect 67546 243335 67602 243344
rect 67364 240032 67416 240038
rect 67364 239974 67416 239980
rect 67270 222864 67326 222873
rect 67270 222799 67326 222808
rect 67652 214606 67680 295423
rect 67730 282432 67786 282441
rect 67730 282367 67786 282376
rect 67744 236706 67772 282367
rect 156788 262200 156840 262206
rect 156788 262142 156840 262148
rect 67822 250064 67878 250073
rect 67822 249999 67878 250008
rect 67732 236700 67784 236706
rect 67732 236642 67784 236648
rect 67836 224262 67864 249999
rect 67916 248464 67968 248470
rect 67916 248406 67968 248412
rect 67928 248334 67956 248406
rect 67916 248328 67968 248334
rect 67916 248270 67968 248276
rect 156694 242856 156750 242865
rect 156694 242791 156750 242800
rect 80978 242040 81034 242049
rect 69584 241998 70104 242026
rect 68816 241590 68968 241618
rect 69368 241590 69520 241618
rect 68940 239426 68968 241590
rect 69492 240106 69520 241590
rect 69480 240100 69532 240106
rect 69480 240042 69532 240048
rect 68928 239420 68980 239426
rect 68928 239362 68980 239368
rect 69584 238754 69612 241998
rect 154670 242040 154726 242049
rect 81034 241998 81388 242026
rect 80978 241975 81034 241984
rect 69754 241904 69810 241913
rect 69754 241839 69810 241848
rect 69664 240032 69716 240038
rect 69664 239974 69716 239980
rect 69032 238726 69612 238754
rect 69032 238377 69060 238726
rect 69018 238368 69074 238377
rect 69018 238303 69074 238312
rect 67824 224256 67876 224262
rect 67824 224198 67876 224204
rect 67640 214600 67692 214606
rect 67640 214542 67692 214548
rect 69676 206961 69704 239974
rect 69768 216646 69796 241839
rect 69938 241768 69994 241777
rect 69938 241703 69994 241712
rect 69952 236609 69980 241703
rect 70412 241590 70840 241618
rect 71576 241590 71728 241618
rect 72312 241590 72648 241618
rect 69938 236600 69994 236609
rect 69938 236535 69994 236544
rect 69756 216640 69808 216646
rect 69756 216582 69808 216588
rect 69662 206952 69718 206961
rect 69662 206887 69718 206896
rect 70412 204270 70440 241590
rect 71042 240000 71098 240009
rect 71042 239935 71098 239944
rect 71056 215257 71084 239935
rect 71700 239465 71728 241590
rect 72422 240136 72478 240145
rect 72620 240106 72648 241590
rect 72712 241590 73048 241618
rect 73784 241590 74120 241618
rect 74520 241590 74580 241618
rect 75256 241590 75592 241618
rect 72712 240145 72740 241590
rect 73804 241392 73856 241398
rect 73804 241334 73856 241340
rect 72698 240136 72754 240145
rect 72422 240071 72478 240080
rect 72516 240100 72568 240106
rect 71686 239456 71742 239465
rect 71686 239391 71742 239400
rect 71042 215248 71098 215257
rect 71042 215183 71098 215192
rect 70400 204264 70452 204270
rect 70400 204206 70452 204212
rect 72436 195265 72464 240071
rect 72516 240042 72568 240048
rect 72608 240100 72660 240106
rect 72698 240071 72754 240080
rect 73068 240100 73120 240106
rect 72608 240042 72660 240048
rect 73068 240042 73120 240048
rect 72528 210458 72556 240042
rect 73080 224913 73108 240042
rect 73066 224904 73122 224913
rect 73066 224839 73122 224848
rect 73816 219434 73844 241334
rect 74092 239737 74120 241590
rect 74078 239728 74134 239737
rect 74078 239663 74134 239672
rect 74552 226302 74580 241590
rect 75564 240009 75592 241590
rect 75932 241590 75992 241618
rect 76728 241590 77248 241618
rect 75550 240000 75606 240009
rect 75550 239935 75606 239944
rect 75932 238678 75960 241590
rect 75920 238672 75972 238678
rect 75920 238614 75972 238620
rect 75932 237454 75960 238614
rect 75920 237448 75972 237454
rect 75920 237390 75972 237396
rect 76564 237448 76616 237454
rect 76564 237390 76616 237396
rect 74540 226296 74592 226302
rect 74540 226238 74592 226244
rect 76576 220697 76604 237390
rect 77220 227730 77248 241590
rect 77404 241590 77464 241618
rect 77864 241590 78200 241618
rect 78692 241590 78936 241618
rect 79672 241590 80008 241618
rect 80408 241590 80744 241618
rect 77300 240168 77352 240174
rect 77300 240110 77352 240116
rect 77208 227724 77260 227730
rect 77208 227666 77260 227672
rect 77312 225622 77340 240110
rect 77404 237386 77432 241590
rect 77864 240174 77892 241590
rect 77942 240816 77998 240825
rect 77942 240751 77998 240760
rect 77852 240168 77904 240174
rect 77852 240110 77904 240116
rect 77392 237380 77444 237386
rect 77392 237322 77444 237328
rect 77300 225616 77352 225622
rect 77300 225558 77352 225564
rect 76562 220688 76618 220697
rect 76562 220623 76618 220632
rect 73804 219428 73856 219434
rect 73804 219370 73856 219376
rect 77956 217433 77984 240751
rect 77942 217424 77998 217433
rect 77942 217359 77998 217368
rect 72516 210452 72568 210458
rect 72516 210394 72568 210400
rect 72422 195256 72478 195265
rect 72422 195191 72478 195200
rect 78692 193089 78720 241590
rect 79980 200122 80008 241590
rect 80716 239970 80744 241590
rect 80704 239964 80756 239970
rect 80704 239906 80756 239912
rect 81256 239964 81308 239970
rect 81256 239906 81308 239912
rect 81268 229770 81296 239906
rect 81256 229764 81308 229770
rect 81256 229706 81308 229712
rect 81360 200705 81388 241998
rect 154726 241998 154928 242026
rect 154670 241975 154726 241984
rect 81880 241590 81940 241618
rect 81912 240106 81940 241590
rect 82004 241590 82616 241618
rect 83352 241604 83504 241618
rect 83338 241590 83504 241604
rect 84088 241590 84148 241618
rect 81900 240100 81952 240106
rect 81900 240042 81952 240048
rect 82004 238754 82032 241590
rect 83338 241466 83366 241590
rect 83326 241460 83378 241466
rect 83326 241402 83378 241408
rect 82728 240100 82780 240106
rect 82728 240042 82780 240048
rect 81452 238726 82032 238754
rect 81452 213926 81480 238726
rect 82740 217326 82768 240042
rect 82818 237960 82874 237969
rect 82818 237895 82874 237904
rect 82832 234569 82860 237895
rect 82818 234560 82874 234569
rect 82818 234495 82874 234504
rect 82728 217320 82780 217326
rect 82728 217262 82780 217268
rect 81440 213920 81492 213926
rect 81440 213862 81492 213868
rect 83476 205601 83504 241590
rect 84120 239494 84148 241590
rect 84212 241590 84824 241618
rect 85560 241590 85620 241618
rect 84108 239488 84160 239494
rect 83554 239456 83610 239465
rect 84108 239430 84160 239436
rect 83554 239391 83610 239400
rect 83568 218006 83596 239391
rect 84212 238241 84240 241590
rect 85592 240106 85620 241590
rect 85684 241590 86296 241618
rect 86972 241590 87032 241618
rect 87156 241590 87768 241618
rect 88504 241590 88840 241618
rect 89240 241590 89668 241618
rect 85580 240100 85632 240106
rect 85580 240042 85632 240048
rect 84198 238232 84254 238241
rect 84198 238167 84254 238176
rect 83556 218000 83608 218006
rect 83556 217942 83608 217948
rect 85684 212537 85712 241590
rect 86868 240100 86920 240106
rect 86868 240042 86920 240048
rect 86880 215937 86908 240042
rect 86972 229838 87000 241590
rect 86960 229832 87012 229838
rect 86960 229774 87012 229780
rect 86866 215928 86922 215937
rect 86866 215863 86922 215872
rect 85670 212528 85726 212537
rect 85670 212463 85726 212472
rect 86866 212528 86922 212537
rect 86866 212463 86922 212472
rect 83462 205592 83518 205601
rect 83462 205527 83518 205536
rect 81346 200696 81402 200705
rect 81346 200631 81402 200640
rect 79968 200116 80020 200122
rect 79968 200058 80020 200064
rect 86880 198257 86908 212463
rect 87156 204950 87184 241590
rect 88812 239970 88840 241590
rect 88800 239964 88852 239970
rect 88800 239906 88852 239912
rect 89536 239964 89588 239970
rect 89536 239906 89588 239912
rect 87602 228304 87658 228313
rect 87602 228239 87658 228248
rect 87144 204944 87196 204950
rect 87144 204886 87196 204892
rect 86866 198248 86922 198257
rect 86866 198183 86922 198192
rect 87616 196625 87644 228239
rect 89548 224777 89576 239906
rect 89534 224768 89590 224777
rect 89534 224703 89590 224712
rect 87602 196616 87658 196625
rect 87602 196551 87658 196560
rect 89640 195294 89668 241590
rect 89824 241590 89976 241618
rect 90376 241590 90712 241618
rect 91204 241590 91448 241618
rect 91848 241590 92184 241618
rect 92920 241590 93072 241618
rect 89720 240168 89772 240174
rect 89720 240110 89772 240116
rect 89732 209409 89760 240110
rect 89824 235929 89852 241590
rect 90376 240174 90404 241590
rect 90364 240168 90416 240174
rect 90364 240110 90416 240116
rect 91100 240168 91152 240174
rect 91100 240110 91152 240116
rect 89810 235920 89866 235929
rect 89810 235855 89866 235864
rect 89824 234705 89852 235855
rect 89810 234696 89866 234705
rect 89810 234631 89866 234640
rect 90362 234696 90418 234705
rect 90362 234631 90418 234640
rect 89718 209400 89774 209409
rect 89718 209335 89774 209344
rect 89628 195288 89680 195294
rect 89628 195230 89680 195236
rect 90376 194177 90404 234631
rect 91006 209400 91062 209409
rect 91006 209335 91062 209344
rect 91020 202337 91048 209335
rect 91112 206281 91140 240110
rect 91204 227769 91232 241590
rect 91848 240174 91876 241590
rect 91836 240168 91888 240174
rect 91836 240110 91888 240116
rect 93044 240106 93072 241590
rect 93136 241590 93472 241618
rect 93964 241590 94208 241618
rect 93032 240100 93084 240106
rect 93032 240042 93084 240048
rect 93136 239290 93164 241590
rect 93858 241360 93914 241369
rect 93858 241295 93914 241304
rect 93768 240100 93820 240106
rect 93768 240042 93820 240048
rect 92572 239284 92624 239290
rect 92572 239226 92624 239232
rect 93124 239284 93176 239290
rect 93124 239226 93176 239232
rect 92584 238746 92612 239226
rect 92572 238740 92624 238746
rect 92572 238682 92624 238688
rect 92584 237454 92612 238682
rect 92572 237448 92624 237454
rect 92572 237390 92624 237396
rect 93124 237448 93176 237454
rect 93124 237390 93176 237396
rect 92386 228848 92442 228857
rect 92386 228783 92442 228792
rect 92400 227769 92428 228783
rect 91190 227760 91246 227769
rect 91190 227695 91246 227704
rect 92386 227760 92442 227769
rect 92386 227695 92442 227704
rect 91098 206272 91154 206281
rect 91098 206207 91154 206216
rect 92400 203561 92428 227695
rect 92386 203552 92442 203561
rect 92386 203487 92442 203496
rect 91006 202328 91062 202337
rect 91006 202263 91062 202272
rect 90362 194168 90418 194177
rect 90362 194103 90418 194112
rect 93136 193118 93164 237390
rect 93124 193112 93176 193118
rect 78678 193080 78734 193089
rect 93124 193054 93176 193060
rect 78678 193015 78734 193024
rect 93780 182073 93808 240042
rect 93872 229129 93900 241295
rect 93858 229120 93914 229129
rect 93858 229055 93914 229064
rect 93964 207670 93992 241590
rect 94930 241369 94958 241604
rect 95252 241590 95680 241618
rect 95804 241590 96416 241618
rect 97152 241590 97488 241618
rect 97888 241590 97948 241618
rect 98624 241590 99144 241618
rect 99360 241590 99696 241618
rect 100096 241590 100708 241618
rect 94916 241360 94972 241369
rect 94916 241295 94972 241304
rect 94502 229120 94558 229129
rect 94502 229055 94558 229064
rect 94516 221921 94544 229055
rect 95252 225049 95280 241590
rect 95804 238754 95832 241590
rect 97356 239488 97408 239494
rect 97460 239465 97488 241590
rect 97356 239430 97408 239436
rect 97446 239456 97502 239465
rect 95344 238726 95832 238754
rect 95344 229090 95372 238726
rect 97368 229809 97396 239430
rect 97446 239391 97502 239400
rect 97354 229800 97410 229809
rect 97264 229764 97316 229770
rect 97354 229735 97410 229744
rect 97264 229706 97316 229712
rect 95332 229084 95384 229090
rect 95332 229026 95384 229032
rect 96526 225584 96582 225593
rect 96526 225519 96582 225528
rect 96540 225049 96568 225519
rect 95238 225040 95294 225049
rect 95238 224975 95294 224984
rect 96526 225040 96582 225049
rect 96526 224975 96582 224984
rect 94502 221912 94558 221921
rect 94502 221847 94558 221856
rect 95148 208344 95200 208350
rect 95148 208286 95200 208292
rect 95160 207670 95188 208286
rect 93952 207664 94004 207670
rect 93952 207606 94004 207612
rect 95148 207664 95200 207670
rect 95148 207606 95200 207612
rect 95160 186969 95188 207606
rect 96540 189689 96568 224975
rect 97276 205630 97304 229706
rect 97264 205624 97316 205630
rect 97264 205566 97316 205572
rect 97920 201482 97948 241590
rect 98368 240780 98420 240786
rect 98368 240722 98420 240728
rect 98380 240009 98408 240722
rect 98366 240000 98422 240009
rect 98366 239935 98422 239944
rect 99116 238754 99144 241590
rect 99668 239834 99696 241590
rect 99656 239828 99708 239834
rect 99656 239770 99708 239776
rect 100576 239828 100628 239834
rect 100576 239770 100628 239776
rect 99116 238726 99328 238754
rect 99300 208185 99328 238726
rect 100588 231198 100616 239770
rect 100576 231192 100628 231198
rect 100576 231134 100628 231140
rect 100680 212401 100708 241590
rect 100772 241590 100832 241618
rect 100956 241590 101568 241618
rect 102152 241590 102304 241618
rect 102428 241590 103040 241618
rect 103776 241590 103836 241618
rect 100772 229770 100800 241590
rect 100760 229764 100812 229770
rect 100760 229706 100812 229712
rect 100956 215121 100984 241590
rect 102152 228313 102180 241590
rect 102428 237289 102456 241590
rect 103808 240106 103836 241590
rect 103900 241590 104512 241618
rect 105248 241590 105584 241618
rect 103796 240100 103848 240106
rect 103796 240042 103848 240048
rect 103900 238754 103928 241590
rect 104808 240100 104860 240106
rect 104808 240042 104860 240048
rect 103532 238726 103928 238754
rect 102414 237280 102470 237289
rect 102414 237215 102470 237224
rect 103532 235890 103560 238726
rect 103520 235884 103572 235890
rect 103520 235826 103572 235832
rect 104716 235884 104768 235890
rect 104716 235826 104768 235832
rect 104728 235521 104756 235826
rect 104714 235512 104770 235521
rect 104714 235447 104770 235456
rect 102138 228304 102194 228313
rect 102138 228239 102194 228248
rect 103426 228304 103482 228313
rect 103426 228239 103482 228248
rect 100942 215112 100998 215121
rect 100942 215047 100998 215056
rect 102046 215112 102102 215121
rect 102046 215047 102102 215056
rect 100666 212392 100722 212401
rect 100666 212327 100722 212336
rect 99286 208176 99342 208185
rect 99286 208111 99342 208120
rect 102060 203590 102088 215047
rect 102048 203584 102100 203590
rect 102048 203526 102100 203532
rect 97908 201476 97960 201482
rect 97908 201418 97960 201424
rect 103440 199481 103468 228239
rect 103426 199472 103482 199481
rect 103426 199407 103482 199416
rect 104820 193905 104848 240042
rect 105556 239290 105584 241590
rect 105648 241590 105984 241618
rect 106292 241590 106720 241618
rect 107456 241590 107608 241618
rect 105544 239284 105596 239290
rect 105544 239226 105596 239232
rect 105648 238754 105676 241590
rect 106188 239284 106240 239290
rect 106188 239226 106240 239232
rect 104912 238726 105676 238754
rect 104912 233238 104940 238726
rect 104900 233232 104952 233238
rect 104900 233174 104952 233180
rect 105544 229832 105596 229838
rect 105544 229774 105596 229780
rect 105556 206922 105584 229774
rect 106200 209778 106228 239226
rect 106292 234433 106320 241590
rect 106278 234424 106334 234433
rect 106278 234359 106334 234368
rect 106188 209772 106240 209778
rect 106188 209714 106240 209720
rect 105544 206916 105596 206922
rect 105544 206858 105596 206864
rect 104806 193896 104862 193905
rect 104806 193831 104862 193840
rect 107580 191049 107608 241590
rect 108178 241369 108206 241604
rect 108928 241590 108988 241618
rect 108164 241360 108220 241369
rect 108164 241295 108220 241304
rect 108960 239494 108988 241590
rect 109052 241590 109664 241618
rect 110400 241590 110736 241618
rect 108948 239488 109000 239494
rect 108948 239430 109000 239436
rect 109052 236745 109080 241590
rect 110708 239970 110736 241590
rect 111122 241466 111150 241604
rect 111812 241590 111872 241618
rect 112608 241590 113036 241618
rect 111110 241460 111162 241466
rect 111110 241402 111162 241408
rect 110696 239964 110748 239970
rect 110696 239906 110748 239912
rect 111708 239964 111760 239970
rect 111708 239906 111760 239912
rect 109038 236736 109094 236745
rect 109038 236671 109094 236680
rect 108304 231192 108356 231198
rect 108304 231134 108356 231140
rect 108316 213761 108344 231134
rect 109682 229800 109738 229809
rect 109682 229735 109738 229744
rect 109696 216481 109724 229735
rect 111720 227662 111748 239906
rect 111812 230353 111840 241590
rect 111798 230344 111854 230353
rect 111798 230279 111854 230288
rect 111708 227656 111760 227662
rect 111708 227598 111760 227604
rect 113008 217297 113036 241590
rect 113192 241590 113344 241618
rect 114080 241590 114508 241618
rect 114816 241590 115152 241618
rect 113192 238610 113220 241590
rect 113180 238604 113232 238610
rect 113180 238546 113232 238552
rect 114282 232656 114338 232665
rect 114282 232591 114338 232600
rect 114296 231810 114324 232591
rect 114284 231804 114336 231810
rect 114284 231746 114336 231752
rect 113086 230344 113142 230353
rect 113086 230279 113142 230288
rect 112994 217288 113050 217297
rect 112994 217223 113050 217232
rect 109682 216472 109738 216481
rect 109682 216407 109738 216416
rect 108302 213752 108358 213761
rect 108302 213687 108358 213696
rect 113100 196761 113128 230279
rect 114480 206990 114508 241590
rect 114652 240100 114704 240106
rect 114652 240042 114704 240048
rect 114664 233209 114692 240042
rect 115124 239154 115152 241590
rect 115216 241590 115552 241618
rect 115952 241590 116288 241618
rect 117024 241590 117268 241618
rect 115216 240106 115244 241590
rect 115204 240100 115256 240106
rect 115204 240042 115256 240048
rect 115112 239148 115164 239154
rect 115112 239090 115164 239096
rect 115848 239148 115900 239154
rect 115848 239090 115900 239096
rect 114650 233200 114706 233209
rect 114650 233135 114706 233144
rect 115860 228410 115888 239090
rect 115020 228404 115072 228410
rect 115020 228346 115072 228352
rect 115848 228404 115900 228410
rect 115848 228346 115900 228352
rect 115032 223553 115060 228346
rect 115952 226273 115980 241590
rect 115938 226264 115994 226273
rect 115938 226199 115994 226208
rect 115952 225049 115980 226199
rect 115938 225040 115994 225049
rect 115938 224975 115994 224984
rect 117134 225040 117190 225049
rect 117134 224975 117190 224984
rect 115018 223544 115074 223553
rect 115018 223479 115074 223488
rect 114468 206984 114520 206990
rect 114468 206926 114520 206932
rect 113086 196752 113142 196761
rect 113086 196687 113142 196696
rect 107566 191040 107622 191049
rect 107566 190975 107622 190984
rect 96526 189680 96582 189689
rect 96526 189615 96582 189624
rect 95146 186960 95202 186969
rect 95146 186895 95202 186904
rect 110328 186380 110380 186386
rect 110328 186322 110380 186328
rect 106186 185192 106242 185201
rect 106186 185127 106242 185136
rect 100666 185056 100722 185065
rect 100666 184991 100722 185000
rect 98826 182200 98882 182209
rect 98826 182135 98882 182144
rect 93766 182064 93822 182073
rect 93766 181999 93822 182008
rect 97262 179480 97318 179489
rect 97262 179415 97318 179424
rect 97276 176905 97304 179415
rect 98840 177585 98868 182135
rect 98826 177576 98882 177585
rect 98826 177511 98882 177520
rect 97262 176896 97318 176905
rect 97262 176831 97318 176840
rect 100680 176769 100708 184991
rect 102046 183696 102102 183705
rect 102046 183631 102102 183640
rect 102060 177585 102088 183631
rect 103336 182232 103388 182238
rect 103336 182174 103388 182180
rect 102046 177576 102102 177585
rect 102046 177511 102102 177520
rect 103348 176769 103376 182174
rect 106200 177585 106228 185127
rect 108118 180840 108174 180849
rect 108118 180775 108174 180784
rect 108132 177585 108160 180775
rect 110340 177585 110368 186322
rect 117148 184249 117176 224975
rect 117240 195945 117268 241590
rect 117424 241590 117760 241618
rect 117976 241590 118312 241618
rect 119048 241590 119384 241618
rect 119784 241590 119936 241618
rect 120520 241590 120856 241618
rect 117320 239216 117372 239222
rect 117320 239158 117372 239164
rect 117332 210361 117360 239158
rect 117424 219201 117452 241590
rect 117976 239222 118004 241590
rect 119356 240106 119384 241590
rect 119344 240100 119396 240106
rect 119344 240042 119396 240048
rect 117964 239216 118016 239222
rect 117964 239158 118016 239164
rect 119908 231169 119936 241590
rect 119988 240100 120040 240106
rect 119988 240042 120040 240048
rect 119894 231160 119950 231169
rect 119894 231095 119950 231104
rect 117410 219192 117466 219201
rect 117410 219127 117466 219136
rect 117318 210352 117374 210361
rect 117318 210287 117374 210296
rect 120000 198121 120028 240042
rect 120828 239290 120856 241590
rect 120920 241590 121256 241618
rect 121992 241590 122328 241618
rect 122728 241590 122788 241618
rect 120816 239284 120868 239290
rect 120816 239226 120868 239232
rect 120920 238754 120948 241590
rect 121642 239728 121698 239737
rect 121642 239663 121698 239672
rect 121368 239284 121420 239290
rect 121368 239226 121420 239232
rect 120092 238726 120948 238754
rect 120092 202881 120120 238726
rect 120078 202872 120134 202881
rect 120078 202807 120134 202816
rect 121380 200025 121408 239226
rect 121656 238678 121684 239663
rect 122300 239601 122328 241590
rect 122286 239592 122342 239601
rect 122286 239527 122342 239536
rect 121644 238672 121696 238678
rect 121644 238614 121696 238620
rect 122102 236872 122158 236881
rect 122102 236807 122158 236816
rect 122116 220833 122144 236807
rect 122102 220824 122158 220833
rect 122102 220759 122158 220768
rect 122760 200802 122788 241590
rect 122852 241590 123464 241618
rect 124200 241590 124260 241618
rect 122852 209545 122880 241590
rect 123484 232552 123536 232558
rect 123484 232494 123536 232500
rect 123496 209681 123524 232494
rect 124232 215286 124260 241590
rect 124324 241590 124936 241618
rect 125612 241590 125672 241618
rect 126408 241590 126928 241618
rect 127144 241590 127204 241618
rect 124220 215280 124272 215286
rect 124220 215222 124272 215228
rect 124324 210526 124352 241590
rect 125612 235890 125640 241590
rect 125600 235884 125652 235890
rect 125600 235826 125652 235832
rect 124312 210520 124364 210526
rect 124312 210462 124364 210468
rect 123482 209672 123538 209681
rect 123482 209607 123538 209616
rect 122838 209536 122894 209545
rect 122838 209471 122894 209480
rect 126900 202774 126928 241590
rect 127176 240106 127204 241590
rect 127268 241590 127880 241618
rect 128616 241590 128952 241618
rect 129352 241590 129688 241618
rect 127164 240100 127216 240106
rect 127164 240042 127216 240048
rect 127268 238754 127296 241590
rect 128268 240100 128320 240106
rect 128268 240042 128320 240048
rect 126992 238726 127296 238754
rect 126992 219366 127020 238726
rect 126980 219360 127032 219366
rect 126980 219302 127032 219308
rect 128280 215121 128308 240042
rect 128924 239290 128952 241590
rect 128912 239284 128964 239290
rect 128912 239226 128964 239232
rect 129556 239284 129608 239290
rect 129556 239226 129608 239232
rect 129004 236768 129056 236774
rect 129004 236710 129056 236716
rect 128266 215112 128322 215121
rect 128266 215047 128322 215056
rect 129016 202842 129044 236710
rect 129568 231266 129596 239226
rect 129556 231260 129608 231266
rect 129556 231202 129608 231208
rect 129660 213625 129688 241590
rect 129752 241590 130088 241618
rect 130824 241590 130976 241618
rect 131560 241590 131896 241618
rect 132296 241590 132448 241618
rect 133032 241590 133368 241618
rect 129752 224641 129780 241590
rect 129738 224632 129794 224641
rect 129738 224567 129794 224576
rect 130948 222154 130976 241590
rect 131868 240106 131896 241590
rect 131856 240100 131908 240106
rect 131856 240042 131908 240048
rect 132316 240100 132368 240106
rect 132316 240042 132368 240048
rect 131026 224632 131082 224641
rect 131026 224567 131082 224576
rect 130936 222148 130988 222154
rect 130936 222090 130988 222096
rect 129646 213616 129702 213625
rect 129646 213551 129702 213560
rect 129004 202836 129056 202842
rect 129004 202778 129056 202784
rect 126888 202768 126940 202774
rect 126888 202710 126940 202716
rect 122748 200796 122800 200802
rect 122748 200738 122800 200744
rect 121366 200016 121422 200025
rect 121366 199951 121422 199960
rect 119986 198112 120042 198121
rect 119986 198047 120042 198056
rect 117226 195936 117282 195945
rect 117226 195871 117282 195880
rect 118608 190528 118660 190534
rect 118608 190470 118660 190476
rect 117134 184240 117190 184249
rect 117134 184175 117190 184184
rect 114376 182300 114428 182306
rect 114376 182242 114428 182248
rect 110694 179616 110750 179625
rect 110694 179551 110750 179560
rect 106186 177576 106242 177585
rect 106186 177511 106242 177520
rect 108118 177576 108174 177585
rect 108118 177511 108174 177520
rect 110326 177576 110382 177585
rect 110326 177511 110382 177520
rect 110708 177177 110736 179551
rect 113732 178084 113784 178090
rect 113732 178026 113784 178032
rect 110694 177168 110750 177177
rect 110694 177103 110750 177112
rect 113744 176769 113772 178026
rect 114388 177585 114416 182242
rect 115848 178152 115900 178158
rect 115848 178094 115900 178100
rect 114374 177576 114430 177585
rect 114374 177511 114430 177520
rect 115860 176769 115888 178094
rect 118620 177449 118648 190470
rect 122748 189100 122800 189106
rect 122748 189042 122800 189048
rect 119528 179512 119580 179518
rect 119528 179454 119580 179460
rect 118606 177440 118662 177449
rect 118606 177375 118662 177384
rect 119540 176769 119568 179454
rect 120816 178016 120868 178022
rect 120816 177958 120868 177964
rect 120828 176769 120856 177958
rect 122760 177585 122788 189042
rect 125508 187740 125560 187746
rect 125508 187682 125560 187688
rect 124864 183592 124916 183598
rect 124864 183534 124916 183540
rect 124036 180940 124088 180946
rect 124036 180882 124088 180888
rect 124048 177585 124076 180882
rect 124876 178022 124904 183534
rect 124864 178016 124916 178022
rect 124864 177958 124916 177964
rect 125520 177585 125548 187682
rect 126888 186448 126940 186454
rect 126888 186390 126940 186396
rect 126900 177585 126928 186390
rect 130936 185020 130988 185026
rect 130936 184962 130988 184968
rect 129464 179444 129516 179450
rect 129464 179386 129516 179392
rect 122746 177576 122802 177585
rect 122746 177511 122802 177520
rect 124034 177576 124090 177585
rect 124034 177511 124090 177520
rect 125506 177576 125562 177585
rect 125506 177511 125562 177520
rect 126886 177576 126942 177585
rect 126886 177511 126942 177520
rect 129476 176769 129504 179386
rect 130948 177585 130976 184962
rect 131040 183161 131068 224567
rect 132328 223514 132356 240042
rect 132316 223508 132368 223514
rect 132316 223450 132368 223456
rect 132420 216578 132448 241590
rect 133340 239766 133368 241590
rect 133708 241590 133768 241618
rect 134504 241590 135116 241618
rect 135240 241590 135300 241618
rect 133328 239760 133380 239766
rect 133328 239702 133380 239708
rect 132408 216572 132460 216578
rect 132408 216514 132460 216520
rect 133144 214600 133196 214606
rect 133144 214542 133196 214548
rect 133156 205465 133184 214542
rect 133708 211041 133736 241590
rect 133788 239760 133840 239766
rect 133788 239702 133840 239708
rect 133694 211032 133750 211041
rect 133694 210967 133750 210976
rect 133800 207670 133828 239702
rect 135088 238754 135116 241590
rect 135088 238726 135208 238754
rect 133788 207664 133840 207670
rect 133788 207606 133840 207612
rect 133142 205456 133198 205465
rect 133142 205391 133198 205400
rect 135180 196654 135208 238726
rect 135272 230217 135300 241590
rect 135364 241590 135976 241618
rect 136652 241590 136712 241618
rect 136836 241590 137448 241618
rect 138032 241590 138184 241618
rect 138676 241604 138920 241618
rect 138676 241590 138934 241604
rect 135364 235793 135392 241590
rect 135350 235784 135406 235793
rect 135350 235719 135406 235728
rect 135258 230208 135314 230217
rect 135258 230143 135314 230152
rect 136546 230208 136602 230217
rect 136546 230143 136602 230152
rect 136560 200841 136588 230143
rect 136652 212430 136680 241590
rect 136836 237153 136864 241590
rect 136822 237144 136878 237153
rect 136822 237079 136878 237088
rect 136836 236774 136864 237079
rect 136824 236768 136876 236774
rect 136824 236710 136876 236716
rect 137282 236736 137338 236745
rect 137282 236671 137338 236680
rect 137296 235657 137324 236671
rect 137282 235648 137338 235657
rect 137282 235583 137338 235592
rect 138032 233986 138060 241590
rect 138020 233980 138072 233986
rect 138020 233922 138072 233928
rect 138018 232656 138074 232665
rect 138018 232591 138074 232600
rect 138032 230489 138060 232591
rect 138018 230480 138074 230489
rect 138018 230415 138074 230424
rect 138676 220561 138704 241590
rect 138906 241505 138934 241590
rect 139596 241590 139656 241618
rect 140056 241590 140392 241618
rect 141128 241590 141464 241618
rect 141864 241590 142108 241618
rect 142600 241590 142936 241618
rect 143152 241590 143488 241618
rect 143888 241590 144224 241618
rect 138892 241496 138948 241505
rect 138892 241431 138948 241440
rect 139400 240168 139452 240174
rect 139400 240110 139452 240116
rect 139124 231192 139176 231198
rect 139124 231134 139176 231140
rect 139136 226302 139164 231134
rect 139216 231124 139268 231130
rect 139216 231066 139268 231072
rect 139228 226302 139256 231066
rect 139124 226296 139176 226302
rect 139124 226238 139176 226244
rect 139216 226296 139268 226302
rect 139216 226238 139268 226244
rect 138662 220552 138718 220561
rect 138662 220487 138718 220496
rect 136640 212424 136692 212430
rect 136640 212366 136692 212372
rect 136546 200832 136602 200841
rect 136546 200767 136602 200776
rect 139412 198626 139440 240110
rect 139492 236768 139544 236774
rect 139492 236710 139544 236716
rect 139504 235890 139532 236710
rect 139492 235884 139544 235890
rect 139492 235826 139544 235832
rect 139596 235278 139624 241590
rect 140056 240174 140084 241590
rect 140044 240168 140096 240174
rect 140044 240110 140096 240116
rect 141436 239290 141464 241590
rect 141424 239284 141476 239290
rect 141424 239226 141476 239232
rect 141976 239284 142028 239290
rect 141976 239226 142028 239232
rect 139584 235272 139636 235278
rect 139584 235214 139636 235220
rect 139492 231872 139544 231878
rect 139492 231814 139544 231820
rect 139504 230382 139532 231814
rect 139492 230376 139544 230382
rect 139492 230318 139544 230324
rect 140780 229764 140832 229770
rect 140780 229706 140832 229712
rect 140792 224330 140820 229706
rect 140780 224324 140832 224330
rect 140780 224266 140832 224272
rect 141422 215928 141478 215937
rect 141422 215863 141478 215872
rect 141436 202201 141464 215863
rect 141988 215218 142016 239226
rect 141976 215212 142028 215218
rect 141976 215154 142028 215160
rect 141422 202192 141478 202201
rect 141422 202127 141478 202136
rect 139400 198620 139452 198626
rect 139400 198562 139452 198568
rect 135168 196648 135220 196654
rect 135168 196590 135220 196596
rect 142080 193225 142108 241590
rect 142908 240106 142936 241590
rect 143460 241097 143488 241590
rect 143446 241088 143502 241097
rect 143446 241023 143502 241032
rect 142896 240100 142948 240106
rect 142896 240042 142948 240048
rect 143448 240100 143500 240106
rect 143448 240042 143500 240048
rect 143632 240100 143684 240106
rect 143632 240042 143684 240048
rect 143356 231260 143408 231266
rect 143356 231202 143408 231208
rect 143368 230450 143396 231202
rect 143356 230444 143408 230450
rect 143356 230386 143408 230392
rect 142158 229120 142214 229129
rect 142158 229055 142214 229064
rect 142172 227662 142200 229055
rect 142160 227656 142212 227662
rect 142160 227598 142212 227604
rect 143460 226273 143488 240042
rect 143644 235958 143672 240042
rect 144196 239290 144224 241590
rect 144288 241590 144624 241618
rect 144932 241590 145360 241618
rect 145576 241590 146096 241618
rect 146832 241590 147168 241618
rect 144288 240106 144316 241590
rect 144276 240100 144328 240106
rect 144276 240042 144328 240048
rect 144184 239284 144236 239290
rect 144184 239226 144236 239232
rect 144828 239284 144880 239290
rect 144828 239226 144880 239232
rect 143632 235952 143684 235958
rect 143632 235894 143684 235900
rect 144184 235952 144236 235958
rect 144184 235894 144236 235900
rect 144196 228721 144224 235894
rect 144182 228712 144238 228721
rect 144182 228647 144238 228656
rect 144736 228404 144788 228410
rect 144736 228346 144788 228352
rect 144092 228336 144144 228342
rect 144748 228313 144776 228346
rect 144092 228278 144144 228284
rect 144734 228304 144790 228313
rect 144104 227633 144132 228278
rect 144734 228239 144790 228248
rect 144090 227624 144146 227633
rect 144090 227559 144146 227568
rect 143446 226264 143502 226273
rect 143446 226199 143502 226208
rect 142804 224256 142856 224262
rect 142804 224198 142856 224204
rect 142816 216617 142844 224198
rect 142802 216608 142858 216617
rect 142802 216543 142858 216552
rect 144840 193866 144868 239226
rect 144932 204241 144960 241590
rect 145576 238754 145604 241590
rect 147140 239290 147168 241590
rect 147508 241590 147568 241618
rect 148304 241590 148732 241618
rect 149040 241590 149100 241618
rect 147128 239284 147180 239290
rect 147128 239226 147180 239232
rect 145024 238726 145604 238754
rect 145024 228585 145052 238726
rect 145010 228576 145066 228585
rect 145010 228511 145066 228520
rect 147508 213858 147536 241590
rect 147588 239284 147640 239290
rect 147588 239226 147640 239232
rect 147496 213852 147548 213858
rect 147496 213794 147548 213800
rect 147600 205329 147628 239226
rect 148704 238754 148732 241590
rect 148704 238726 149008 238754
rect 148324 233980 148376 233986
rect 148324 233922 148376 233928
rect 147680 233912 147732 233918
rect 147680 233854 147732 233860
rect 147692 231810 147720 233854
rect 147680 231804 147732 231810
rect 147680 231746 147732 231752
rect 147680 227044 147732 227050
rect 147680 226986 147732 226992
rect 147692 226302 147720 226986
rect 147680 226296 147732 226302
rect 147680 226238 147732 226244
rect 147772 226296 147824 226302
rect 147772 226238 147824 226244
rect 147784 225593 147812 226238
rect 147770 225584 147826 225593
rect 147770 225519 147826 225528
rect 148336 223582 148364 233922
rect 148324 223576 148376 223582
rect 148324 223518 148376 223524
rect 147586 205320 147642 205329
rect 147586 205255 147642 205264
rect 144918 204232 144974 204241
rect 144918 204167 144974 204176
rect 144828 193860 144880 193866
rect 144828 193802 144880 193808
rect 142066 193216 142122 193225
rect 142066 193151 142122 193160
rect 148876 184952 148928 184958
rect 148876 184894 148928 184900
rect 133788 183660 133840 183666
rect 133788 183602 133840 183608
rect 131026 183152 131082 183161
rect 131026 183087 131082 183096
rect 132408 180872 132460 180878
rect 132408 180814 132460 180820
rect 132420 177585 132448 180814
rect 133800 177585 133828 183602
rect 148888 177585 148916 184894
rect 148980 179353 149008 238726
rect 149072 236842 149100 241590
rect 149164 241590 149776 241618
rect 150512 241590 150848 241618
rect 151248 241590 151768 241618
rect 151984 241590 152320 241618
rect 152720 241590 153056 241618
rect 153456 241590 153792 241618
rect 149060 236836 149112 236842
rect 149060 236778 149112 236784
rect 149058 236600 149114 236609
rect 149058 236535 149114 236544
rect 149072 235958 149100 236535
rect 149060 235952 149112 235958
rect 149060 235894 149112 235900
rect 149164 226001 149192 241590
rect 150820 240281 150848 241590
rect 150806 240272 150862 240281
rect 150806 240207 150862 240216
rect 149244 236836 149296 236842
rect 149244 236778 149296 236784
rect 149256 234598 149284 236778
rect 149334 236056 149390 236065
rect 149334 235991 149390 236000
rect 149244 234592 149296 234598
rect 149244 234534 149296 234540
rect 149348 232665 149376 235991
rect 150440 235272 150492 235278
rect 150440 235214 150492 235220
rect 149334 232656 149390 232665
rect 149334 232591 149390 232600
rect 150452 232558 150480 235214
rect 150440 232552 150492 232558
rect 150440 232494 150492 232500
rect 149150 225992 149206 226001
rect 149150 225927 149206 225936
rect 151740 224262 151768 241590
rect 152292 240009 152320 241590
rect 153028 241233 153056 241590
rect 153108 241528 153160 241534
rect 153108 241470 153160 241476
rect 153120 241369 153148 241470
rect 153106 241360 153162 241369
rect 153106 241295 153162 241304
rect 153014 241224 153070 241233
rect 153014 241159 153070 241168
rect 153382 240272 153438 240281
rect 153382 240207 153438 240216
rect 153292 240100 153344 240106
rect 153292 240042 153344 240048
rect 152278 240000 152334 240009
rect 152278 239935 152334 239944
rect 153106 240000 153162 240009
rect 153106 239935 153162 239944
rect 153014 237416 153070 237425
rect 153014 237351 153070 237360
rect 152738 231976 152794 231985
rect 152738 231911 152794 231920
rect 152752 230382 152780 231911
rect 152740 230376 152792 230382
rect 152740 230318 152792 230324
rect 153028 227633 153056 237351
rect 153014 227624 153070 227633
rect 153014 227559 153070 227568
rect 151728 224256 151780 224262
rect 151728 224198 151780 224204
rect 150346 217560 150402 217569
rect 150346 217495 150402 217504
rect 150360 213761 150388 217495
rect 150346 213752 150402 213761
rect 150346 213687 150402 213696
rect 151082 213752 151138 213761
rect 151082 213687 151138 213696
rect 151096 187105 151124 213687
rect 153120 199345 153148 239935
rect 153304 237289 153332 240042
rect 153396 238649 153424 240207
rect 153764 239970 153792 241590
rect 153856 241590 154192 241618
rect 153856 240106 153884 241590
rect 153844 240100 153896 240106
rect 153844 240042 153896 240048
rect 153752 239964 153804 239970
rect 153752 239906 153804 239912
rect 154488 239964 154540 239970
rect 154488 239906 154540 239912
rect 153382 238640 153438 238649
rect 153382 238575 153438 238584
rect 153290 237280 153346 237289
rect 153290 237215 153346 237224
rect 153106 199336 153162 199345
rect 153106 199271 153162 199280
rect 154500 189825 154528 239906
rect 154684 237017 154712 241975
rect 155664 241590 155908 241618
rect 155682 240816 155738 240825
rect 155682 240751 155738 240760
rect 154670 237008 154726 237017
rect 154670 236943 154726 236952
rect 155696 235657 155724 240751
rect 155682 235648 155738 235657
rect 155682 235583 155738 235592
rect 155224 234660 155276 234666
rect 155224 234602 155276 234608
rect 155236 227050 155264 234602
rect 155774 232520 155830 232529
rect 155774 232455 155830 232464
rect 155788 231305 155816 232455
rect 155774 231296 155830 231305
rect 155774 231231 155830 231240
rect 155224 227044 155276 227050
rect 155224 226986 155276 226992
rect 154580 226364 154632 226370
rect 154580 226306 154632 226312
rect 154592 223582 154620 226306
rect 154580 223576 154632 223582
rect 154580 223518 154632 223524
rect 155224 223576 155276 223582
rect 155224 223518 155276 223524
rect 155236 195974 155264 223518
rect 155224 195968 155276 195974
rect 155224 195910 155276 195916
rect 154486 189816 154542 189825
rect 154486 189751 154542 189760
rect 151082 187096 151138 187105
rect 151082 187031 151138 187040
rect 155880 181529 155908 241590
rect 156386 241505 156414 241604
rect 156708 241534 156736 242791
rect 156696 241528 156748 241534
rect 156372 241496 156428 241505
rect 156696 241470 156748 241476
rect 156372 241431 156428 241440
rect 155960 237312 156012 237318
rect 155958 237280 155960 237289
rect 156012 237280 156014 237289
rect 155958 237215 156014 237224
rect 156604 231736 156656 231742
rect 156604 231678 156656 231684
rect 156510 220688 156566 220697
rect 156510 220623 156566 220632
rect 156524 220114 156552 220623
rect 156512 220108 156564 220114
rect 156512 220050 156564 220056
rect 156616 202881 156644 231678
rect 156800 226370 156828 262142
rect 157996 260166 158024 329802
rect 158088 300121 158116 345646
rect 158166 332752 158222 332761
rect 158166 332687 158222 332696
rect 158180 320890 158208 332687
rect 158168 320884 158220 320890
rect 158168 320826 158220 320832
rect 158074 300112 158130 300121
rect 158074 300047 158130 300056
rect 157984 260160 158036 260166
rect 157984 260102 158036 260108
rect 157982 254552 158038 254561
rect 157982 254487 158038 254496
rect 156972 242956 157024 242962
rect 156972 242898 157024 242904
rect 156880 242208 156932 242214
rect 156880 242150 156932 242156
rect 156892 231198 156920 242150
rect 156984 236774 157012 242898
rect 157338 240136 157394 240145
rect 157338 240071 157394 240080
rect 156972 236768 157024 236774
rect 156972 236710 157024 236716
rect 156880 231192 156932 231198
rect 156880 231134 156932 231140
rect 157352 228857 157380 240071
rect 157996 231742 158024 254487
rect 158088 242185 158116 300047
rect 158168 284980 158220 284986
rect 158168 284922 158220 284928
rect 158074 242176 158130 242185
rect 158074 242111 158130 242120
rect 158180 240009 158208 284922
rect 158640 277817 158668 351834
rect 159376 341601 159404 459546
rect 162136 437442 162164 516122
rect 162228 510610 162256 525778
rect 167644 521008 167696 521014
rect 167644 520950 167696 520956
rect 162216 510604 162268 510610
rect 162216 510546 162268 510552
rect 165528 467900 165580 467906
rect 165528 467842 165580 467848
rect 162124 437436 162176 437442
rect 162124 437378 162176 437384
rect 162768 436144 162820 436150
rect 162768 436086 162820 436092
rect 162676 421592 162728 421598
rect 162676 421534 162728 421540
rect 161388 411324 161440 411330
rect 161388 411266 161440 411272
rect 159456 378820 159508 378826
rect 159456 378762 159508 378768
rect 159362 341592 159418 341601
rect 159362 341527 159418 341536
rect 159364 332648 159416 332654
rect 159364 332590 159416 332596
rect 158718 326496 158774 326505
rect 158718 326431 158774 326440
rect 158732 325718 158760 326431
rect 158720 325712 158772 325718
rect 158720 325654 158772 325660
rect 158902 324456 158958 324465
rect 158902 324391 158958 324400
rect 158718 324320 158774 324329
rect 158718 324255 158774 324264
rect 158732 323066 158760 324255
rect 158812 324216 158864 324222
rect 158812 324158 158864 324164
rect 158824 323241 158852 324158
rect 158810 323232 158866 323241
rect 158810 323167 158866 323176
rect 158720 323060 158772 323066
rect 158720 323002 158772 323008
rect 158720 322856 158772 322862
rect 158720 322798 158772 322804
rect 158732 322153 158760 322798
rect 158718 322144 158774 322153
rect 158718 322079 158774 322088
rect 158718 321056 158774 321065
rect 158718 320991 158774 321000
rect 158732 320210 158760 320991
rect 158916 320793 158944 324391
rect 158902 320784 158958 320793
rect 158902 320719 158958 320728
rect 158720 320204 158772 320210
rect 158720 320146 158772 320152
rect 158812 320136 158864 320142
rect 158812 320078 158864 320084
rect 158718 319152 158774 319161
rect 158718 319087 158774 319096
rect 158626 277808 158682 277817
rect 158626 277743 158682 277752
rect 158640 277438 158668 277743
rect 158628 277432 158680 277438
rect 158628 277374 158680 277380
rect 158628 262132 158680 262138
rect 158628 262074 158680 262080
rect 158640 261497 158668 262074
rect 158626 261488 158682 261497
rect 158626 261423 158682 261432
rect 158166 240000 158222 240009
rect 158166 239935 158222 239944
rect 158640 234705 158668 261423
rect 158626 234696 158682 234705
rect 158626 234631 158682 234640
rect 158076 234524 158128 234530
rect 158076 234466 158128 234472
rect 157984 231736 158036 231742
rect 157984 231678 158036 231684
rect 157338 228848 157394 228857
rect 157338 228783 157394 228792
rect 156788 226364 156840 226370
rect 156788 226306 156840 226312
rect 156696 220040 156748 220046
rect 156696 219982 156748 219988
rect 156602 202872 156658 202881
rect 156708 202842 156736 219982
rect 158088 216345 158116 234466
rect 158732 233889 158760 319087
rect 158824 318889 158852 320078
rect 158810 318880 158866 318889
rect 158810 318815 158866 318824
rect 158812 315988 158864 315994
rect 158812 315930 158864 315936
rect 158824 315625 158852 315930
rect 158810 315616 158866 315625
rect 158810 315551 158866 315560
rect 158810 313440 158866 313449
rect 158810 313375 158866 313384
rect 158824 313342 158852 313375
rect 158812 313336 158864 313342
rect 158812 313278 158864 313284
rect 158902 311264 158958 311273
rect 158902 311199 158958 311208
rect 158916 310554 158944 311199
rect 158904 310548 158956 310554
rect 158904 310490 158956 310496
rect 158812 310480 158864 310486
rect 158812 310422 158864 310428
rect 158824 310185 158852 310422
rect 158810 310176 158866 310185
rect 158810 310111 158866 310120
rect 158812 308984 158864 308990
rect 158812 308926 158864 308932
rect 158824 308009 158852 308926
rect 158810 308000 158866 308009
rect 158810 307935 158866 307944
rect 158810 306912 158866 306921
rect 158810 306847 158866 306856
rect 158824 306406 158852 306847
rect 158812 306400 158864 306406
rect 158812 306342 158864 306348
rect 158810 305824 158866 305833
rect 158810 305759 158866 305768
rect 158824 305046 158852 305759
rect 158812 305040 158864 305046
rect 158812 304982 158864 304988
rect 158810 304736 158866 304745
rect 158810 304671 158866 304680
rect 158824 304026 158852 304671
rect 158812 304020 158864 304026
rect 158812 303962 158864 303968
rect 158812 303680 158864 303686
rect 158810 303648 158812 303657
rect 158864 303648 158866 303657
rect 158810 303583 158866 303592
rect 158810 301472 158866 301481
rect 158810 301407 158866 301416
rect 158824 300150 158852 301407
rect 158994 300384 159050 300393
rect 158994 300319 158996 300328
rect 159048 300319 159050 300328
rect 158996 300290 159048 300296
rect 158812 300144 158864 300150
rect 158812 300086 158864 300092
rect 158812 299464 158864 299470
rect 158812 299406 158864 299412
rect 158824 298217 158852 299406
rect 158810 298208 158866 298217
rect 158810 298143 158866 298152
rect 158810 297120 158866 297129
rect 158810 297055 158866 297064
rect 158824 296750 158852 297055
rect 158812 296744 158864 296750
rect 158812 296686 158864 296692
rect 158810 296032 158866 296041
rect 158810 295967 158812 295976
rect 158864 295967 158866 295976
rect 158812 295938 158864 295944
rect 158812 295316 158864 295322
rect 158812 295258 158864 295264
rect 158824 294953 158852 295258
rect 158810 294944 158866 294953
rect 158810 294879 158866 294888
rect 158902 293856 158958 293865
rect 158902 293791 158958 293800
rect 158810 293040 158866 293049
rect 158810 292975 158866 292984
rect 158824 292670 158852 292975
rect 158812 292664 158864 292670
rect 158812 292606 158864 292612
rect 158916 292602 158944 293791
rect 158904 292596 158956 292602
rect 158904 292538 158956 292544
rect 158810 291952 158866 291961
rect 158810 291887 158866 291896
rect 158824 291242 158852 291887
rect 158812 291236 158864 291242
rect 158812 291178 158864 291184
rect 158810 290864 158866 290873
rect 158810 290799 158866 290808
rect 158824 289882 158852 290799
rect 158812 289876 158864 289882
rect 158812 289818 158864 289824
rect 158902 289776 158958 289785
rect 158902 289711 158958 289720
rect 158812 289264 158864 289270
rect 158812 289206 158864 289212
rect 158824 288697 158852 289206
rect 158810 288688 158866 288697
rect 158810 288623 158866 288632
rect 158916 288386 158944 289711
rect 158904 288380 158956 288386
rect 158904 288322 158956 288328
rect 158810 287600 158866 287609
rect 158810 287535 158866 287544
rect 158824 287094 158852 287535
rect 158812 287088 158864 287094
rect 158812 287030 158864 287036
rect 158812 286340 158864 286346
rect 158812 286282 158864 286288
rect 158824 285433 158852 286282
rect 158810 285424 158866 285433
rect 158810 285359 158866 285368
rect 158810 284880 158866 284889
rect 158810 284815 158866 284824
rect 158824 282169 158852 284815
rect 158810 282160 158866 282169
rect 158810 282095 158866 282104
rect 158810 281072 158866 281081
rect 158810 281007 158866 281016
rect 158824 280294 158852 281007
rect 158812 280288 158864 280294
rect 158812 280230 158864 280236
rect 159376 279478 159404 332590
rect 159468 330546 159496 378762
rect 160742 355328 160798 355337
rect 160742 355263 160798 355272
rect 159548 343664 159600 343670
rect 159548 343606 159600 343612
rect 159456 330540 159508 330546
rect 159456 330482 159508 330488
rect 159560 328506 159588 343606
rect 160098 336968 160154 336977
rect 160098 336903 160154 336912
rect 160112 334801 160140 336903
rect 160098 334792 160154 334801
rect 160098 334727 160154 334736
rect 159638 334248 159694 334257
rect 159638 334183 159694 334192
rect 159456 328500 159508 328506
rect 159456 328442 159508 328448
rect 159548 328500 159600 328506
rect 159548 328442 159600 328448
rect 159468 322318 159496 328442
rect 159560 327593 159588 328442
rect 159546 327584 159602 327593
rect 159546 327519 159602 327528
rect 159652 325009 159680 334183
rect 160100 330540 160152 330546
rect 160100 330482 160152 330488
rect 159730 328672 159786 328681
rect 159730 328607 159786 328616
rect 159638 325000 159694 325009
rect 159638 324935 159694 324944
rect 159744 323649 159772 328607
rect 159730 323640 159786 323649
rect 159730 323575 159786 323584
rect 159456 322312 159508 322318
rect 159456 322254 159508 322260
rect 160008 316736 160060 316742
rect 160006 316704 160008 316713
rect 160060 316704 160062 316713
rect 160006 316639 160062 316648
rect 160008 301504 160060 301510
rect 160008 301446 160060 301452
rect 159364 279472 159416 279478
rect 159364 279414 159416 279420
rect 159822 278896 159878 278905
rect 159822 278831 159878 278840
rect 158812 277364 158864 277370
rect 158812 277306 158864 277312
rect 158824 276729 158852 277306
rect 158810 276720 158866 276729
rect 158810 276655 158866 276664
rect 158812 275936 158864 275942
rect 158812 275878 158864 275884
rect 158824 275641 158852 275878
rect 158810 275632 158866 275641
rect 158810 275567 158866 275576
rect 159836 275330 159864 278831
rect 159824 275324 159876 275330
rect 159824 275266 159876 275272
rect 159546 274952 159602 274961
rect 159546 274887 159602 274896
rect 158812 274644 158864 274650
rect 158812 274586 158864 274592
rect 158824 274553 158852 274586
rect 158810 274544 158866 274553
rect 158810 274479 158866 274488
rect 158810 273456 158866 273465
rect 158810 273391 158866 273400
rect 158824 273290 158852 273391
rect 158812 273284 158864 273290
rect 158812 273226 158864 273232
rect 158810 271280 158866 271289
rect 158810 271215 158866 271224
rect 158824 270842 158852 271215
rect 158812 270836 158864 270842
rect 158812 270778 158864 270784
rect 158810 269104 158866 269113
rect 158810 269039 158812 269048
rect 158864 269039 158866 269048
rect 158812 269010 158864 269016
rect 159362 268016 159418 268025
rect 159362 267951 159418 267960
rect 158812 266348 158864 266354
rect 158812 266290 158864 266296
rect 158824 265849 158852 266290
rect 158810 265840 158866 265849
rect 158810 265775 158866 265784
rect 158812 264920 158864 264926
rect 158812 264862 158864 264868
rect 158824 264761 158852 264862
rect 158810 264752 158866 264761
rect 158810 264687 158866 264696
rect 158812 263560 158864 263566
rect 158812 263502 158864 263508
rect 158824 262585 158852 263502
rect 158810 262576 158866 262585
rect 158810 262511 158866 262520
rect 158902 260400 158958 260409
rect 158902 260335 158958 260344
rect 158916 259486 158944 260335
rect 158904 259480 158956 259486
rect 158904 259422 158956 259428
rect 158810 258224 158866 258233
rect 158810 258159 158866 258168
rect 158824 258126 158852 258159
rect 158812 258120 158864 258126
rect 158812 258062 158864 258068
rect 159270 257136 159326 257145
rect 159270 257071 159272 257080
rect 159324 257071 159326 257080
rect 159272 257042 159324 257048
rect 158810 256320 158866 256329
rect 158810 256255 158866 256264
rect 158824 255338 158852 256255
rect 158812 255332 158864 255338
rect 158812 255274 158864 255280
rect 158902 255232 158958 255241
rect 158902 255167 158958 255176
rect 158812 254584 158864 254590
rect 158812 254526 158864 254532
rect 158824 254153 158852 254526
rect 158810 254144 158866 254153
rect 158810 254079 158866 254088
rect 158916 253978 158944 255167
rect 158904 253972 158956 253978
rect 158904 253914 158956 253920
rect 158810 253056 158866 253065
rect 158810 252991 158866 253000
rect 158824 252686 158852 252991
rect 158812 252680 158864 252686
rect 158812 252622 158864 252628
rect 158902 251968 158958 251977
rect 159376 251938 159404 267951
rect 159456 262268 159508 262274
rect 159456 262210 159508 262216
rect 158902 251903 158958 251912
rect 159364 251932 159416 251938
rect 158812 251184 158864 251190
rect 158812 251126 158864 251132
rect 158824 250889 158852 251126
rect 158810 250880 158866 250889
rect 158810 250815 158866 250824
rect 158810 249792 158866 249801
rect 158810 249727 158866 249736
rect 158824 248470 158852 249727
rect 158916 249257 158944 251903
rect 159364 251874 159416 251880
rect 158902 249248 158958 249257
rect 158902 249183 158958 249192
rect 159468 248713 159496 262210
rect 159560 262206 159588 274887
rect 160020 270450 160048 301446
rect 160112 300354 160140 330482
rect 160756 324222 160784 355263
rect 160834 334520 160890 334529
rect 160834 334455 160890 334464
rect 160744 324216 160796 324222
rect 160744 324158 160796 324164
rect 160848 318170 160876 334455
rect 160836 318164 160888 318170
rect 160836 318106 160888 318112
rect 161296 316736 161348 316742
rect 161296 316678 161348 316684
rect 160742 309904 160798 309913
rect 160742 309839 160798 309848
rect 160100 300348 160152 300354
rect 160100 300290 160152 300296
rect 160098 284336 160154 284345
rect 160098 284271 160154 284280
rect 160112 282198 160140 284271
rect 160100 282192 160152 282198
rect 160100 282134 160152 282140
rect 160020 270422 160140 270450
rect 159548 262200 159600 262206
rect 159548 262142 159600 262148
rect 159640 252612 159692 252618
rect 159640 252554 159692 252560
rect 159454 248704 159510 248713
rect 159454 248639 159510 248648
rect 158812 248464 158864 248470
rect 158812 248406 158864 248412
rect 159548 247104 159600 247110
rect 159548 247046 159600 247052
rect 158810 246528 158866 246537
rect 158810 246463 158866 246472
rect 158824 246430 158852 246463
rect 158812 246424 158864 246430
rect 158812 246366 158864 246372
rect 158810 245440 158866 245449
rect 158810 245375 158866 245384
rect 158824 244934 158852 245375
rect 158812 244928 158864 244934
rect 158812 244870 158864 244876
rect 158810 244352 158866 244361
rect 158810 244287 158812 244296
rect 158864 244287 158866 244296
rect 158812 244258 158864 244264
rect 158810 243264 158866 243273
rect 158810 243199 158866 243208
rect 158824 243030 158852 243199
rect 158812 243024 158864 243030
rect 158812 242966 158864 242972
rect 159456 240848 159508 240854
rect 159456 240790 159508 240796
rect 159362 234696 159418 234705
rect 159362 234631 159418 234640
rect 158718 233880 158774 233889
rect 158718 233815 158774 233824
rect 158720 217320 158772 217326
rect 158720 217262 158772 217268
rect 158074 216336 158130 216345
rect 158074 216271 158130 216280
rect 158732 210497 158760 217262
rect 158718 210488 158774 210497
rect 158718 210423 158774 210432
rect 156602 202807 156658 202816
rect 156696 202836 156748 202842
rect 156616 191826 156644 202807
rect 156696 202778 156748 202784
rect 156604 191820 156656 191826
rect 156604 191762 156656 191768
rect 159376 190466 159404 234631
rect 159468 224913 159496 240790
rect 159560 235521 159588 247046
rect 159652 241466 159680 252554
rect 160006 247616 160062 247625
rect 160112 247602 160140 270422
rect 160062 247574 160140 247602
rect 160006 247551 160062 247560
rect 159640 241460 159692 241466
rect 159640 241402 159692 241408
rect 160756 237318 160784 309839
rect 160836 304020 160888 304026
rect 160836 303962 160888 303968
rect 160848 294545 160876 303962
rect 160928 300348 160980 300354
rect 160928 300290 160980 300296
rect 160834 294536 160890 294545
rect 160834 294471 160890 294480
rect 160940 292505 160968 300290
rect 160926 292496 160982 292505
rect 160926 292431 160982 292440
rect 160836 280832 160888 280838
rect 160836 280774 160888 280780
rect 160848 257106 160876 280774
rect 160928 280288 160980 280294
rect 160928 280230 160980 280236
rect 160940 276690 160968 280230
rect 160928 276684 160980 276690
rect 160928 276626 160980 276632
rect 161308 268394 161336 316678
rect 161400 313993 161428 411266
rect 162124 387864 162176 387870
rect 162124 387806 162176 387812
rect 161478 363624 161534 363633
rect 161478 363559 161534 363568
rect 161386 313984 161442 313993
rect 161386 313919 161442 313928
rect 161296 268388 161348 268394
rect 161296 268330 161348 268336
rect 160836 257100 160888 257106
rect 160836 257042 160888 257048
rect 160744 237312 160796 237318
rect 160744 237254 160796 237260
rect 159546 235512 159602 235521
rect 159546 235447 159602 235456
rect 160098 230480 160154 230489
rect 160098 230415 160100 230424
rect 160152 230415 160154 230424
rect 160100 230386 160152 230392
rect 159454 224904 159510 224913
rect 159454 224839 159510 224848
rect 160848 194041 160876 257042
rect 160928 250504 160980 250510
rect 160928 250446 160980 250452
rect 160940 240786 160968 250446
rect 161020 242276 161072 242282
rect 161020 242218 161072 242224
rect 160928 240780 160980 240786
rect 160928 240722 160980 240728
rect 161032 238649 161060 242218
rect 161018 238640 161074 238649
rect 161018 238575 161074 238584
rect 161492 237402 161520 363559
rect 161570 343768 161626 343777
rect 161570 343703 161626 343712
rect 161584 322862 161612 343703
rect 162136 330546 162164 387806
rect 162688 362234 162716 421534
rect 162676 362228 162728 362234
rect 162676 362170 162728 362176
rect 162124 330540 162176 330546
rect 162124 330482 162176 330488
rect 162122 329760 162178 329769
rect 162122 329695 162178 329704
rect 162136 324970 162164 329695
rect 162124 324964 162176 324970
rect 162124 324906 162176 324912
rect 161572 322856 161624 322862
rect 161572 322798 161624 322804
rect 161570 317792 161626 317801
rect 161570 317727 161626 317736
rect 161584 312594 161612 317727
rect 161572 312588 161624 312594
rect 161572 312530 161624 312536
rect 162216 290488 162268 290494
rect 162216 290430 162268 290436
rect 162124 287088 162176 287094
rect 162124 287030 162176 287036
rect 162136 246362 162164 287030
rect 162228 275942 162256 290430
rect 162780 289270 162808 436086
rect 164884 396772 164936 396778
rect 164884 396714 164936 396720
rect 163412 380996 163464 381002
rect 163412 380938 163464 380944
rect 163424 374678 163452 380938
rect 162860 374672 162912 374678
rect 162860 374614 162912 374620
rect 163412 374672 163464 374678
rect 163412 374614 163464 374620
rect 162872 308990 162900 374614
rect 163502 369064 163558 369073
rect 163502 368999 163558 369008
rect 163320 334076 163372 334082
rect 163320 334018 163372 334024
rect 162950 328264 163006 328273
rect 162950 328199 163006 328208
rect 162964 322250 162992 328199
rect 163332 327758 163360 334018
rect 163320 327752 163372 327758
rect 163320 327694 163372 327700
rect 162952 322244 163004 322250
rect 162952 322186 163004 322192
rect 162860 308984 162912 308990
rect 162860 308926 162912 308932
rect 162768 289264 162820 289270
rect 162768 289206 162820 289212
rect 162780 289105 162808 289206
rect 162766 289096 162822 289105
rect 162766 289031 162822 289040
rect 162216 275936 162268 275942
rect 162216 275878 162268 275884
rect 162216 270836 162268 270842
rect 162216 270778 162268 270784
rect 162228 257378 162256 270778
rect 162216 257372 162268 257378
rect 162216 257314 162268 257320
rect 162216 256012 162268 256018
rect 162216 255954 162268 255960
rect 162124 246356 162176 246362
rect 162124 246298 162176 246304
rect 161308 237374 161520 237402
rect 161308 230489 161336 237374
rect 162122 233336 162178 233345
rect 162122 233271 162178 233280
rect 161386 230616 161442 230625
rect 161386 230551 161442 230560
rect 161294 230480 161350 230489
rect 161294 230415 161350 230424
rect 160834 194032 160890 194041
rect 160834 193967 160890 193976
rect 159364 190460 159416 190466
rect 159364 190402 159416 190408
rect 159376 188358 159404 190402
rect 161400 188465 161428 230551
rect 162136 190369 162164 233271
rect 162228 231169 162256 255954
rect 162768 253972 162820 253978
rect 162768 253914 162820 253920
rect 162780 251870 162808 253914
rect 162768 251864 162820 251870
rect 162768 251806 162820 251812
rect 162306 245712 162362 245721
rect 162306 245647 162362 245656
rect 162320 234530 162348 245647
rect 162308 234524 162360 234530
rect 162308 234466 162360 234472
rect 162214 231160 162270 231169
rect 162214 231095 162270 231104
rect 163516 222154 163544 368999
rect 164240 362228 164292 362234
rect 164240 362170 164292 362176
rect 163596 341556 163648 341562
rect 163596 341498 163648 341504
rect 163608 331809 163636 341498
rect 163594 331800 163650 331809
rect 163594 331735 163650 331744
rect 163688 320204 163740 320210
rect 163688 320146 163740 320152
rect 163594 301608 163650 301617
rect 163594 301543 163650 301552
rect 163608 235793 163636 301543
rect 163700 300218 163728 320146
rect 164252 310486 164280 362170
rect 164790 331936 164846 331945
rect 164790 331871 164846 331880
rect 164804 329118 164832 331871
rect 164792 329112 164844 329118
rect 164792 329054 164844 329060
rect 164896 318753 164924 396714
rect 164976 328500 165028 328506
rect 164976 328442 165028 328448
rect 164882 318744 164938 318753
rect 164882 318679 164938 318688
rect 164882 317384 164938 317393
rect 164882 317319 164938 317328
rect 164240 310480 164292 310486
rect 164240 310422 164292 310428
rect 163688 300212 163740 300218
rect 163688 300154 163740 300160
rect 164148 270564 164200 270570
rect 164148 270506 164200 270512
rect 163688 269136 163740 269142
rect 163688 269078 163740 269084
rect 163594 235784 163650 235793
rect 163594 235719 163650 235728
rect 163504 222148 163556 222154
rect 163504 222090 163556 222096
rect 163700 211138 163728 269078
rect 164160 242282 164188 270506
rect 164148 242276 164200 242282
rect 164148 242218 164200 242224
rect 164146 235784 164202 235793
rect 164146 235719 164202 235728
rect 163778 231704 163834 231713
rect 163778 231639 163834 231648
rect 162768 211132 162820 211138
rect 162768 211074 162820 211080
rect 163688 211132 163740 211138
rect 163688 211074 163740 211080
rect 162780 210526 162808 211074
rect 163792 211041 163820 231639
rect 164160 231130 164188 235719
rect 164148 231124 164200 231130
rect 164148 231066 164200 231072
rect 164896 226302 164924 317319
rect 164988 301578 165016 328442
rect 165540 316538 165568 467842
rect 166264 460216 166316 460222
rect 166264 460158 166316 460164
rect 166276 434722 166304 460158
rect 166908 443760 166960 443766
rect 166908 443702 166960 443708
rect 165620 434716 165672 434722
rect 165620 434658 165672 434664
rect 166264 434716 166316 434722
rect 166264 434658 166316 434664
rect 165632 434042 165660 434658
rect 165620 434036 165672 434042
rect 165620 433978 165672 433984
rect 165068 316532 165120 316538
rect 165068 316474 165120 316480
rect 165528 316532 165580 316538
rect 165528 316474 165580 316480
rect 165080 316062 165108 316474
rect 165068 316056 165120 316062
rect 165068 315998 165120 316004
rect 164976 301572 165028 301578
rect 164976 301514 165028 301520
rect 164976 287700 165028 287706
rect 164976 287642 165028 287648
rect 164988 240825 165016 287642
rect 165080 286346 165108 315998
rect 165528 310480 165580 310486
rect 165528 310422 165580 310428
rect 165540 309874 165568 310422
rect 165528 309868 165580 309874
rect 165528 309810 165580 309816
rect 165632 301510 165660 433978
rect 166920 400994 166948 443702
rect 166908 400988 166960 400994
rect 166908 400930 166960 400936
rect 166262 389192 166318 389201
rect 166262 389127 166318 389136
rect 166276 302433 166304 389127
rect 167000 377528 167052 377534
rect 167000 377470 167052 377476
rect 166908 369164 166960 369170
rect 166908 369106 166960 369112
rect 166356 360324 166408 360330
rect 166356 360266 166408 360272
rect 166368 316742 166396 360266
rect 166920 320618 166948 369106
rect 167012 361554 167040 377470
rect 167000 361548 167052 361554
rect 167000 361490 167052 361496
rect 167012 360330 167040 361490
rect 167000 360324 167052 360330
rect 167000 360266 167052 360272
rect 167656 338337 167684 520950
rect 169036 445777 169064 538834
rect 170496 535560 170548 535566
rect 170496 535502 170548 535508
rect 170402 527776 170458 527785
rect 170402 527711 170458 527720
rect 168470 445768 168526 445777
rect 168470 445703 168526 445712
rect 169022 445768 169078 445777
rect 169022 445703 169078 445712
rect 168484 444553 168512 445703
rect 168470 444544 168526 444553
rect 168470 444479 168526 444488
rect 167736 423700 167788 423706
rect 167736 423642 167788 423648
rect 167748 364334 167776 423642
rect 168380 390584 168432 390590
rect 168380 390526 168432 390532
rect 167748 364306 167868 364334
rect 167840 351218 167868 364306
rect 167828 351212 167880 351218
rect 167828 351154 167880 351160
rect 167734 341592 167790 341601
rect 167734 341527 167790 341536
rect 167642 338328 167698 338337
rect 167642 338263 167698 338272
rect 166908 320612 166960 320618
rect 166908 320554 166960 320560
rect 166920 320142 166948 320554
rect 166908 320136 166960 320142
rect 166908 320078 166960 320084
rect 167656 319530 167684 338263
rect 167644 319524 167696 319530
rect 167644 319466 167696 319472
rect 166998 318744 167054 318753
rect 166998 318679 167054 318688
rect 166448 318164 166500 318170
rect 166448 318106 166500 318112
rect 166356 316736 166408 316742
rect 166356 316678 166408 316684
rect 166262 302424 166318 302433
rect 166262 302359 166318 302368
rect 165620 301504 165672 301510
rect 166080 301504 166132 301510
rect 165620 301446 165672 301452
rect 166078 301472 166080 301481
rect 166132 301472 166134 301481
rect 166078 301407 166134 301416
rect 165160 297424 165212 297430
rect 165160 297366 165212 297372
rect 165068 286340 165120 286346
rect 165068 286282 165120 286288
rect 165172 277370 165200 297366
rect 165528 279812 165580 279818
rect 165528 279754 165580 279760
rect 165160 277364 165212 277370
rect 165160 277306 165212 277312
rect 165068 258732 165120 258738
rect 165068 258674 165120 258680
rect 165080 246265 165108 258674
rect 165066 246256 165122 246265
rect 165066 246191 165122 246200
rect 165540 243386 165568 279754
rect 166276 263566 166304 302359
rect 166460 286006 166488 318106
rect 166540 308984 166592 308990
rect 166540 308926 166592 308932
rect 166448 286000 166500 286006
rect 166448 285942 166500 285948
rect 166356 285728 166408 285734
rect 166356 285670 166408 285676
rect 166264 263560 166316 263566
rect 166264 263502 166316 263508
rect 166264 259480 166316 259486
rect 166264 259422 166316 259428
rect 165080 243358 165568 243386
rect 164974 240816 165030 240825
rect 164974 240751 165030 240760
rect 164884 226296 164936 226302
rect 164884 226238 164936 226244
rect 164148 222148 164200 222154
rect 164148 222090 164200 222096
rect 164160 221542 164188 222090
rect 164148 221536 164200 221542
rect 164148 221478 164200 221484
rect 163778 211032 163834 211041
rect 163778 210967 163834 210976
rect 162768 210520 162820 210526
rect 162768 210462 162820 210468
rect 162122 190360 162178 190369
rect 162122 190295 162178 190304
rect 161386 188456 161442 188465
rect 161386 188391 161442 188400
rect 162780 188358 162808 210462
rect 163792 200114 163820 210967
rect 165080 201482 165108 243358
rect 165540 243001 165568 243358
rect 165526 242992 165582 243001
rect 165526 242927 165582 242936
rect 165250 242176 165306 242185
rect 165250 242111 165306 242120
rect 165160 240780 165212 240786
rect 165160 240722 165212 240728
rect 165172 227730 165200 240722
rect 165264 237153 165292 242111
rect 165250 237144 165306 237153
rect 165250 237079 165306 237088
rect 165160 227724 165212 227730
rect 165160 227666 165212 227672
rect 165068 201476 165120 201482
rect 165068 201418 165120 201424
rect 163608 200086 163820 200114
rect 163504 195968 163556 195974
rect 163504 195910 163556 195916
rect 159364 188352 159416 188358
rect 159364 188294 159416 188300
rect 162768 188352 162820 188358
rect 162768 188294 162820 188300
rect 162124 183660 162176 183666
rect 162124 183602 162176 183608
rect 155866 181520 155922 181529
rect 155866 181455 155922 181464
rect 148966 179344 149022 179353
rect 148966 179279 149022 179288
rect 130934 177576 130990 177585
rect 130934 177511 130990 177520
rect 132406 177576 132462 177585
rect 132406 177511 132462 177520
rect 133786 177576 133842 177585
rect 133786 177511 133842 177520
rect 148874 177576 148930 177585
rect 148874 177511 148930 177520
rect 158996 176792 159048 176798
rect 100666 176760 100722 176769
rect 100666 176695 100722 176704
rect 103334 176760 103390 176769
rect 103334 176695 103390 176704
rect 113730 176760 113786 176769
rect 113730 176695 113786 176704
rect 115846 176760 115902 176769
rect 115846 176695 115902 176704
rect 119526 176760 119582 176769
rect 119526 176695 119582 176704
rect 120814 176760 120870 176769
rect 120814 176695 120870 176704
rect 127070 176760 127126 176769
rect 127070 176695 127072 176704
rect 127124 176695 127126 176704
rect 129462 176760 129518 176769
rect 129462 176695 129518 176704
rect 158994 176760 158996 176769
rect 159048 176760 159050 176769
rect 158994 176695 159050 176704
rect 127072 176666 127124 176672
rect 135720 176656 135772 176662
rect 135720 176598 135772 176604
rect 134432 175976 134484 175982
rect 134432 175918 134484 175924
rect 134444 175409 134472 175918
rect 135732 175409 135760 176598
rect 134430 175400 134486 175409
rect 134430 175335 134486 175344
rect 135718 175400 135774 175409
rect 135718 175335 135774 175344
rect 162136 175234 162164 183602
rect 163516 176633 163544 195910
rect 163608 195362 163636 200086
rect 166172 198008 166224 198014
rect 166172 197950 166224 197956
rect 163596 195356 163648 195362
rect 163596 195298 163648 195304
rect 163596 193860 163648 193866
rect 163596 193802 163648 193808
rect 163608 187241 163636 193802
rect 166184 193186 166212 197950
rect 166172 193180 166224 193186
rect 166172 193122 166224 193128
rect 163594 187232 163650 187241
rect 163594 187167 163650 187176
rect 164884 186448 164936 186454
rect 164884 186390 164936 186396
rect 163502 176624 163558 176633
rect 163502 176559 163558 176568
rect 162124 175228 162176 175234
rect 162124 175170 162176 175176
rect 164896 171086 164924 186390
rect 164976 182300 165028 182306
rect 164976 182242 165028 182248
rect 164988 173233 165016 182242
rect 166276 180033 166304 259422
rect 166368 251190 166396 285670
rect 166552 281450 166580 308926
rect 166816 296064 166868 296070
rect 166816 296006 166868 296012
rect 166540 281444 166592 281450
rect 166540 281386 166592 281392
rect 166356 251184 166408 251190
rect 166356 251126 166408 251132
rect 166828 224777 166856 296006
rect 166908 276004 166960 276010
rect 166908 275946 166960 275952
rect 166814 224768 166870 224777
rect 166814 224703 166870 224712
rect 166828 224233 166856 224703
rect 166814 224224 166870 224233
rect 166814 224159 166870 224168
rect 166920 198626 166948 275946
rect 166908 198620 166960 198626
rect 166908 198562 166960 198568
rect 166920 197985 166948 198562
rect 166906 197976 166962 197985
rect 166906 197911 166962 197920
rect 166356 195288 166408 195294
rect 166356 195230 166408 195236
rect 166262 180024 166318 180033
rect 166262 179959 166318 179968
rect 166264 176792 166316 176798
rect 166264 176734 166316 176740
rect 165436 176724 165488 176730
rect 165436 176666 165488 176672
rect 165448 174593 165476 176666
rect 165528 175976 165580 175982
rect 165528 175918 165580 175924
rect 165540 175166 165568 175918
rect 165528 175160 165580 175166
rect 165528 175102 165580 175108
rect 165526 174992 165582 175001
rect 165526 174927 165582 174936
rect 165434 174584 165490 174593
rect 165434 174519 165490 174528
rect 164974 173224 165030 173233
rect 164974 173159 165030 173168
rect 164884 171080 164936 171086
rect 164884 171022 164936 171028
rect 165540 161430 165568 174927
rect 165528 161424 165580 161430
rect 165528 161366 165580 161372
rect 166276 149054 166304 176734
rect 166368 172514 166396 195230
rect 166540 180940 166592 180946
rect 166540 180882 166592 180888
rect 166446 179616 166502 179625
rect 166446 179551 166502 179560
rect 166356 172508 166408 172514
rect 166356 172450 166408 172456
rect 166460 162858 166488 179551
rect 166552 169726 166580 180882
rect 166540 169720 166592 169726
rect 166540 169662 166592 169668
rect 166448 162852 166500 162858
rect 166448 162794 166500 162800
rect 166264 149048 166316 149054
rect 166264 148990 166316 148996
rect 67454 125216 67510 125225
rect 67454 125151 67510 125160
rect 67362 123584 67418 123593
rect 67362 123519 67418 123528
rect 67376 93226 67404 123519
rect 67364 93220 67416 93226
rect 67364 93162 67416 93168
rect 67468 82142 67496 125151
rect 166264 124228 166316 124234
rect 166264 124170 166316 124176
rect 164884 113824 164936 113830
rect 164884 113766 164936 113772
rect 67638 102368 67694 102377
rect 67638 102303 67694 102312
rect 67546 100736 67602 100745
rect 67546 100671 67602 100680
rect 67560 90370 67588 100671
rect 67548 90364 67600 90370
rect 67548 90306 67600 90312
rect 67456 82136 67508 82142
rect 67456 82078 67508 82084
rect 67652 74526 67680 102303
rect 100666 94752 100722 94761
rect 100666 94687 100722 94696
rect 120630 94752 120686 94761
rect 120630 94687 120686 94696
rect 100680 93906 100708 94687
rect 111156 94512 111208 94518
rect 106922 94480 106978 94489
rect 111156 94454 111208 94460
rect 106922 94415 106978 94424
rect 100668 93900 100720 93906
rect 100668 93842 100720 93848
rect 103426 93256 103482 93265
rect 97264 93220 97316 93226
rect 103426 93191 103482 93200
rect 97264 93162 97316 93168
rect 85118 92440 85174 92449
rect 85118 92375 85174 92384
rect 75274 91216 75330 91225
rect 75274 91151 75330 91160
rect 75288 87650 75316 91151
rect 85132 91118 85160 92375
rect 86866 91352 86922 91361
rect 86866 91287 86922 91296
rect 86774 91216 86830 91225
rect 86774 91151 86830 91160
rect 85120 91112 85172 91118
rect 85120 91054 85172 91060
rect 75276 87644 75328 87650
rect 75276 87586 75328 87592
rect 86788 82822 86816 91151
rect 86776 82816 86828 82822
rect 86776 82758 86828 82764
rect 70306 76664 70362 76673
rect 70306 76599 70362 76608
rect 67640 74520 67692 74526
rect 67640 74462 67692 74468
rect 68926 71088 68982 71097
rect 68926 71023 68982 71032
rect 67180 22840 67232 22846
rect 67180 22782 67232 22788
rect 66720 7608 66772 7614
rect 66720 7550 66772 7556
rect 65524 3528 65576 3534
rect 65524 3470 65576 3476
rect 66168 3528 66220 3534
rect 66168 3470 66220 3476
rect 65536 480 65564 3470
rect 66732 480 66760 7550
rect 68940 3534 68968 71023
rect 70214 68368 70270 68377
rect 70214 68303 70270 68312
rect 70228 3534 70256 68303
rect 67916 3528 67968 3534
rect 67916 3470 67968 3476
rect 68928 3528 68980 3534
rect 68928 3470 68980 3476
rect 69112 3528 69164 3534
rect 69112 3470 69164 3476
rect 70216 3528 70268 3534
rect 70216 3470 70268 3476
rect 67928 480 67956 3470
rect 69124 480 69152 3470
rect 70320 480 70348 76599
rect 73066 73808 73122 73817
rect 73066 73743 73122 73752
rect 71044 46232 71096 46238
rect 71044 46174 71096 46180
rect 71056 3602 71084 46174
rect 71504 10396 71556 10402
rect 71504 10338 71556 10344
rect 71044 3596 71096 3602
rect 71044 3538 71096 3544
rect 71516 480 71544 10338
rect 73080 3534 73108 73743
rect 75826 69592 75882 69601
rect 75826 69527 75882 69536
rect 74448 32496 74500 32502
rect 74448 32438 74500 32444
rect 74460 3534 74488 32438
rect 75840 3534 75868 69527
rect 77206 67008 77262 67017
rect 77206 66943 77262 66952
rect 77220 3534 77248 66943
rect 79966 65648 80022 65657
rect 79966 65583 80022 65592
rect 78588 31136 78640 31142
rect 78588 31078 78640 31084
rect 78496 3596 78548 3602
rect 78496 3538 78548 3544
rect 72608 3528 72660 3534
rect 72608 3470 72660 3476
rect 73068 3528 73120 3534
rect 73068 3470 73120 3476
rect 73804 3528 73856 3534
rect 73804 3470 73856 3476
rect 74448 3528 74500 3534
rect 74448 3470 74500 3476
rect 75000 3528 75052 3534
rect 75000 3470 75052 3476
rect 75828 3528 75880 3534
rect 75828 3470 75880 3476
rect 76196 3528 76248 3534
rect 76196 3470 76248 3476
rect 77208 3528 77260 3534
rect 77208 3470 77260 3476
rect 77392 3528 77444 3534
rect 77392 3470 77444 3476
rect 72620 480 72648 3470
rect 73816 480 73844 3470
rect 75012 480 75040 3470
rect 76208 480 76236 3470
rect 77404 480 77432 3470
rect 78508 1850 78536 3538
rect 78600 3534 78628 31078
rect 79980 6914 80008 65583
rect 84108 60036 84160 60042
rect 84108 59978 84160 59984
rect 81348 26988 81400 26994
rect 81348 26930 81400 26936
rect 79704 6886 80008 6914
rect 78588 3528 78640 3534
rect 78588 3470 78640 3476
rect 78508 1822 78628 1850
rect 78600 480 78628 1822
rect 79704 480 79732 6886
rect 81360 3602 81388 26930
rect 84120 3602 84148 59978
rect 86880 49706 86908 91287
rect 88062 91216 88118 91225
rect 88062 91151 88118 91160
rect 89626 91216 89682 91225
rect 89626 91151 89682 91160
rect 90730 91216 90786 91225
rect 90730 91151 90786 91160
rect 91926 91216 91982 91225
rect 91926 91151 91982 91160
rect 93030 91216 93086 91225
rect 93030 91151 93086 91160
rect 95146 91216 95202 91225
rect 95146 91151 95202 91160
rect 96342 91216 96398 91225
rect 96342 91151 96398 91160
rect 88076 86970 88104 91151
rect 88064 86964 88116 86970
rect 88064 86906 88116 86912
rect 89640 63510 89668 91151
rect 90744 88233 90772 91151
rect 90730 88224 90786 88233
rect 90730 88159 90786 88168
rect 91940 86873 91968 91151
rect 91926 86864 91982 86873
rect 91926 86799 91982 86808
rect 93044 85377 93072 91151
rect 93030 85368 93086 85377
rect 93030 85303 93086 85312
rect 95160 81433 95188 91151
rect 96356 88097 96384 91151
rect 96342 88088 96398 88097
rect 96342 88023 96398 88032
rect 95146 81424 95202 81433
rect 95146 81359 95202 81368
rect 97276 81297 97304 93162
rect 98644 93152 98696 93158
rect 98644 93094 98696 93100
rect 97814 91352 97870 91361
rect 97814 91287 97870 91296
rect 97262 81288 97318 81297
rect 97262 81223 97318 81232
rect 95146 78024 95202 78033
rect 95146 77959 95202 77968
rect 89628 63504 89680 63510
rect 89628 63446 89680 63452
rect 87602 61432 87658 61441
rect 87602 61367 87658 61376
rect 86868 49700 86920 49706
rect 86868 49642 86920 49648
rect 85488 46300 85540 46306
rect 85488 46242 85540 46248
rect 80888 3596 80940 3602
rect 80888 3538 80940 3544
rect 81348 3596 81400 3602
rect 81348 3538 81400 3544
rect 83280 3596 83332 3602
rect 83280 3538 83332 3544
rect 84108 3596 84160 3602
rect 84108 3538 84160 3544
rect 80900 480 80928 3538
rect 82082 2000 82138 2009
rect 82082 1935 82138 1944
rect 82096 480 82124 1935
rect 83292 480 83320 3538
rect 85500 3534 85528 46242
rect 86868 33856 86920 33862
rect 86868 33798 86920 33804
rect 84476 3528 84528 3534
rect 84476 3470 84528 3476
rect 85488 3528 85540 3534
rect 85488 3470 85540 3476
rect 84488 480 84516 3470
rect 85670 3360 85726 3369
rect 85670 3295 85726 3304
rect 85684 480 85712 3295
rect 86880 480 86908 33798
rect 87616 3602 87644 61367
rect 91008 55888 91060 55894
rect 91008 55830 91060 55836
rect 89628 54528 89680 54534
rect 89628 54470 89680 54476
rect 88248 19984 88300 19990
rect 88248 19926 88300 19932
rect 88260 6914 88288 19926
rect 87984 6886 88288 6914
rect 87604 3596 87656 3602
rect 87604 3538 87656 3544
rect 87984 480 88012 6886
rect 89640 3534 89668 54470
rect 91020 3534 91048 55830
rect 93766 51776 93822 51785
rect 93766 51711 93822 51720
rect 91560 9036 91612 9042
rect 91560 8978 91612 8984
rect 89168 3528 89220 3534
rect 89168 3470 89220 3476
rect 89628 3528 89680 3534
rect 89628 3470 89680 3476
rect 90364 3528 90416 3534
rect 90364 3470 90416 3476
rect 91008 3528 91060 3534
rect 91008 3470 91060 3476
rect 89180 480 89208 3470
rect 90376 480 90404 3470
rect 91572 480 91600 8978
rect 93780 3534 93808 51711
rect 95056 44872 95108 44878
rect 95056 44814 95108 44820
rect 95068 3534 95096 44814
rect 92756 3528 92808 3534
rect 92756 3470 92808 3476
rect 93768 3528 93820 3534
rect 93768 3470 93820 3476
rect 93952 3528 94004 3534
rect 93952 3470 94004 3476
rect 95056 3528 95108 3534
rect 95056 3470 95108 3476
rect 92768 480 92796 3470
rect 93964 480 93992 3470
rect 95160 480 95188 77959
rect 97828 73137 97856 91287
rect 97906 91216 97962 91225
rect 97906 91151 97962 91160
rect 97920 84182 97948 91151
rect 97908 84176 97960 84182
rect 97908 84118 97960 84124
rect 98656 75886 98684 93094
rect 100024 91792 100076 91798
rect 100024 91734 100076 91740
rect 99194 91216 99250 91225
rect 99194 91151 99250 91160
rect 98644 75880 98696 75886
rect 98644 75822 98696 75828
rect 97906 75304 97962 75313
rect 97906 75239 97962 75248
rect 97814 73128 97870 73137
rect 97814 73063 97870 73072
rect 96252 14476 96304 14482
rect 96252 14418 96304 14424
rect 96264 480 96292 14418
rect 97920 3534 97948 75239
rect 99208 70378 99236 91151
rect 100036 71738 100064 91734
rect 101954 91352 102010 91361
rect 101954 91287 102010 91296
rect 100666 91216 100722 91225
rect 100666 91151 100722 91160
rect 100680 74458 100708 91151
rect 101968 78674 101996 91287
rect 102046 91216 102102 91225
rect 102046 91151 102102 91160
rect 103334 91216 103390 91225
rect 103440 91186 103468 93191
rect 104162 91488 104218 91497
rect 104162 91423 104218 91432
rect 103334 91151 103390 91160
rect 103428 91180 103480 91186
rect 101956 78668 102008 78674
rect 101956 78610 102008 78616
rect 100668 74452 100720 74458
rect 100668 74394 100720 74400
rect 100024 71732 100076 71738
rect 100024 71674 100076 71680
rect 99196 70372 99248 70378
rect 99196 70314 99248 70320
rect 102060 64870 102088 91151
rect 103348 67590 103376 91151
rect 103428 91122 103480 91128
rect 103336 67584 103388 67590
rect 103336 67526 103388 67532
rect 102048 64864 102100 64870
rect 102048 64806 102100 64812
rect 102046 62928 102102 62937
rect 102046 62863 102102 62872
rect 99288 40792 99340 40798
rect 99288 40734 99340 40740
rect 99300 3534 99328 40734
rect 100668 24132 100720 24138
rect 100668 24074 100720 24080
rect 100680 3534 100708 24074
rect 102060 3534 102088 62863
rect 104176 62082 104204 91423
rect 106186 91352 106242 91361
rect 106186 91287 106242 91296
rect 104438 91216 104494 91225
rect 104438 91151 104494 91160
rect 106094 91216 106150 91225
rect 106094 91151 106150 91160
rect 104452 85513 104480 91151
rect 105544 91112 105596 91118
rect 105544 91054 105596 91060
rect 104438 85504 104494 85513
rect 104438 85439 104494 85448
rect 105556 82657 105584 91054
rect 105542 82648 105598 82657
rect 105542 82583 105598 82592
rect 106108 68950 106136 91151
rect 106096 68944 106148 68950
rect 106096 68886 106148 68892
rect 104164 62076 104216 62082
rect 104164 62018 104216 62024
rect 104808 57248 104860 57254
rect 104808 57190 104860 57196
rect 103428 18624 103480 18630
rect 103428 18566 103480 18572
rect 103440 6914 103468 18566
rect 104820 6914 104848 57190
rect 106200 51066 106228 91287
rect 106936 84153 106964 94415
rect 110142 93256 110198 93265
rect 110142 93191 110198 93200
rect 108120 92540 108172 92546
rect 108120 92482 108172 92488
rect 108132 92449 108160 92482
rect 108118 92440 108174 92449
rect 110156 92410 110184 93191
rect 108118 92375 108174 92384
rect 110144 92404 110196 92410
rect 110144 92346 110196 92352
rect 107566 91352 107622 91361
rect 107566 91287 107622 91296
rect 107474 91216 107530 91225
rect 107474 91151 107530 91160
rect 106922 84144 106978 84153
rect 106922 84079 106978 84088
rect 107488 57934 107516 91151
rect 107580 79966 107608 91287
rect 108670 91216 108726 91225
rect 108304 91180 108356 91186
rect 108670 91151 108726 91160
rect 109222 91216 109278 91225
rect 109222 91151 109278 91160
rect 110142 91216 110198 91225
rect 110142 91151 110198 91160
rect 108304 91122 108356 91128
rect 107568 79960 107620 79966
rect 107568 79902 107620 79908
rect 107568 72548 107620 72554
rect 107568 72490 107620 72496
rect 107476 57928 107528 57934
rect 107476 57870 107528 57876
rect 106188 51060 106240 51066
rect 106188 51002 106240 51008
rect 105544 42084 105596 42090
rect 105544 42026 105596 42032
rect 103348 6886 103468 6914
rect 104544 6886 104848 6914
rect 97448 3528 97500 3534
rect 97448 3470 97500 3476
rect 97908 3528 97960 3534
rect 97908 3470 97960 3476
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 99288 3528 99340 3534
rect 99288 3470 99340 3476
rect 99840 3528 99892 3534
rect 99840 3470 99892 3476
rect 100668 3528 100720 3534
rect 100668 3470 100720 3476
rect 101036 3528 101088 3534
rect 101036 3470 101088 3476
rect 102048 3528 102100 3534
rect 102048 3470 102100 3476
rect 97460 480 97488 3470
rect 98656 480 98684 3470
rect 99852 480 99880 3470
rect 101048 480 101076 3470
rect 102232 2168 102284 2174
rect 102232 2110 102284 2116
rect 102244 480 102272 2110
rect 103348 480 103376 6886
rect 104544 480 104572 6886
rect 105556 2106 105584 42026
rect 106832 11756 106884 11762
rect 106832 11698 106884 11704
rect 105728 4820 105780 4826
rect 105728 4762 105780 4768
rect 105544 2100 105596 2106
rect 105544 2042 105596 2048
rect 105740 480 105768 4762
rect 106844 3466 106872 11698
rect 107580 3534 107608 72490
rect 108316 59362 108344 91122
rect 108684 85542 108712 91151
rect 109236 88262 109264 91151
rect 109224 88256 109276 88262
rect 109224 88198 109276 88204
rect 108672 85536 108724 85542
rect 108672 85478 108724 85484
rect 108948 77988 109000 77994
rect 108948 77930 109000 77936
rect 108304 59356 108356 59362
rect 108304 59298 108356 59304
rect 108960 3534 108988 77930
rect 110156 66230 110184 91151
rect 111064 89004 111116 89010
rect 111064 88946 111116 88952
rect 111076 74497 111104 88946
rect 111168 80034 111196 94454
rect 120644 93974 120672 94687
rect 160742 94480 160798 94489
rect 160742 94415 160798 94424
rect 120632 93968 120684 93974
rect 120632 93910 120684 93916
rect 118238 93528 118294 93537
rect 118238 93463 118294 93472
rect 124126 93528 124182 93537
rect 124126 93463 124182 93472
rect 118252 93158 118280 93463
rect 124140 93226 124168 93463
rect 124128 93220 124180 93226
rect 124128 93162 124180 93168
rect 118240 93152 118292 93158
rect 118240 93094 118292 93100
rect 122104 92540 122156 92546
rect 122104 92482 122156 92488
rect 111246 92440 111302 92449
rect 115754 92440 115810 92449
rect 111246 92375 111302 92384
rect 112444 92404 112496 92410
rect 111260 91118 111288 92375
rect 115754 92375 115810 92384
rect 116766 92440 116822 92449
rect 116766 92375 116822 92384
rect 112444 92346 112496 92352
rect 111338 91896 111394 91905
rect 111338 91831 111394 91840
rect 111248 91112 111300 91118
rect 111248 91054 111300 91060
rect 111352 89729 111380 91831
rect 112166 91216 112222 91225
rect 112166 91151 112222 91160
rect 111338 89720 111394 89729
rect 111338 89655 111394 89664
rect 112180 87961 112208 91151
rect 112166 87952 112222 87961
rect 112166 87887 112222 87896
rect 111156 80028 111208 80034
rect 111156 79970 111208 79976
rect 111706 76800 111762 76809
rect 111706 76735 111762 76744
rect 111062 74488 111118 74497
rect 111062 74423 111118 74432
rect 110144 66224 110196 66230
rect 110144 66166 110196 66172
rect 111616 21480 111668 21486
rect 111616 21422 111668 21428
rect 111628 16574 111656 21422
rect 111536 16546 111656 16574
rect 106924 3528 106976 3534
rect 106924 3470 106976 3476
rect 107568 3528 107620 3534
rect 107568 3470 107620 3476
rect 108120 3528 108172 3534
rect 108120 3470 108172 3476
rect 108948 3528 109000 3534
rect 108948 3470 109000 3476
rect 109316 3528 109368 3534
rect 109316 3470 109368 3476
rect 106832 3460 106884 3466
rect 106832 3402 106884 3408
rect 106936 480 106964 3470
rect 108132 480 108160 3470
rect 109328 480 109356 3470
rect 111536 3126 111564 16546
rect 111720 6914 111748 76735
rect 112456 55214 112484 92346
rect 115478 92168 115534 92177
rect 115478 92103 115534 92112
rect 113086 91216 113142 91225
rect 113086 91151 113142 91160
rect 114374 91216 114430 91225
rect 114374 91151 114430 91160
rect 112536 87644 112588 87650
rect 112536 87586 112588 87592
rect 112548 64802 112576 87586
rect 113100 81394 113128 91151
rect 114388 86902 114416 91151
rect 115296 91112 115348 91118
rect 115296 91054 115348 91060
rect 115204 90364 115256 90370
rect 115204 90306 115256 90312
rect 114376 86896 114428 86902
rect 114376 86838 114428 86844
rect 113088 81388 113140 81394
rect 113088 81330 113140 81336
rect 115216 69018 115244 90306
rect 115308 75818 115336 91054
rect 115492 90409 115520 92103
rect 115768 91050 115796 92375
rect 116582 91896 116638 91905
rect 116582 91831 116638 91840
rect 115756 91044 115808 91050
rect 115756 90986 115808 90992
rect 115478 90400 115534 90409
rect 115478 90335 115534 90344
rect 115296 75812 115348 75818
rect 115296 75754 115348 75760
rect 115204 69012 115256 69018
rect 115204 68954 115256 68960
rect 112536 64796 112588 64802
rect 112536 64738 112588 64744
rect 116596 60722 116624 91831
rect 116780 91118 116808 92375
rect 120722 91896 120778 91905
rect 120722 91831 120778 91840
rect 119894 91760 119950 91769
rect 119894 91695 119950 91704
rect 117134 91216 117190 91225
rect 117134 91151 117190 91160
rect 118054 91216 118110 91225
rect 118054 91151 118110 91160
rect 116768 91112 116820 91118
rect 116768 91054 116820 91060
rect 116584 60716 116636 60722
rect 116584 60658 116636 60664
rect 115848 58676 115900 58682
rect 115848 58618 115900 58624
rect 112444 55208 112496 55214
rect 112444 55150 112496 55156
rect 114468 49020 114520 49026
rect 114468 48962 114520 48968
rect 112444 29708 112496 29714
rect 112444 29650 112496 29656
rect 112456 7682 112484 29650
rect 112812 13184 112864 13190
rect 112812 13126 112864 13132
rect 112444 7676 112496 7682
rect 112444 7618 112496 7624
rect 111628 6886 111748 6914
rect 110512 3120 110564 3126
rect 110512 3062 110564 3068
rect 111524 3120 111576 3126
rect 111524 3062 111576 3068
rect 110524 480 110552 3062
rect 111628 480 111656 6886
rect 112824 480 112852 13126
rect 114480 3466 114508 48962
rect 115860 3466 115888 58618
rect 117148 52426 117176 91151
rect 118068 85241 118096 91151
rect 119908 89690 119936 91695
rect 119986 91216 120042 91225
rect 119986 91151 120042 91160
rect 119896 89684 119948 89690
rect 119896 89626 119948 89632
rect 118054 85232 118110 85241
rect 118054 85167 118110 85176
rect 117226 83600 117282 83609
rect 117226 83535 117282 83544
rect 117136 52420 117188 52426
rect 117136 52362 117188 52368
rect 117240 3466 117268 83535
rect 120000 82521 120028 91151
rect 120736 82793 120764 91831
rect 120722 82784 120778 82793
rect 120722 82719 120778 82728
rect 119986 82512 120042 82521
rect 119986 82447 120042 82456
rect 122116 77178 122144 92482
rect 125784 92472 125836 92478
rect 125782 92440 125784 92449
rect 125836 92440 125838 92449
rect 125782 92375 125838 92384
rect 133142 92440 133198 92449
rect 133142 92375 133144 92384
rect 133196 92375 133198 92384
rect 133144 92346 133196 92352
rect 130750 91760 130806 91769
rect 130750 91695 130806 91704
rect 151634 91760 151690 91769
rect 151634 91695 151690 91704
rect 124034 91488 124090 91497
rect 124034 91423 124090 91432
rect 122286 91216 122342 91225
rect 122286 91151 122342 91160
rect 122300 88330 122328 91151
rect 122288 88324 122340 88330
rect 122288 88266 122340 88272
rect 123484 82136 123536 82142
rect 123484 82078 123536 82084
rect 122104 77172 122156 77178
rect 122104 77114 122156 77120
rect 119986 73944 120042 73953
rect 119986 73879 120042 73888
rect 117596 7676 117648 7682
rect 117596 7618 117648 7624
rect 114008 3460 114060 3466
rect 114008 3402 114060 3408
rect 114468 3460 114520 3466
rect 114468 3402 114520 3408
rect 115204 3460 115256 3466
rect 115204 3402 115256 3408
rect 115848 3460 115900 3466
rect 115848 3402 115900 3408
rect 116400 3460 116452 3466
rect 116400 3402 116452 3408
rect 117228 3460 117280 3466
rect 117228 3402 117280 3408
rect 114020 480 114048 3402
rect 115216 480 115244 3402
rect 116412 480 116440 3402
rect 117608 480 117636 7618
rect 120000 6914 120028 73879
rect 122748 72480 122800 72486
rect 122748 72422 122800 72428
rect 119908 6886 120028 6914
rect 118792 2100 118844 2106
rect 118792 2042 118844 2048
rect 118804 480 118832 2042
rect 119908 480 119936 6886
rect 121090 3496 121146 3505
rect 122760 3466 122788 72422
rect 123496 56574 123524 82078
rect 124048 67522 124076 91423
rect 126794 91352 126850 91361
rect 126794 91287 126850 91296
rect 124126 91216 124182 91225
rect 124126 91151 124182 91160
rect 125414 91216 125470 91225
rect 125414 91151 125470 91160
rect 124036 67516 124088 67522
rect 124036 67458 124088 67464
rect 124140 63442 124168 91151
rect 125428 77246 125456 91151
rect 126808 84114 126836 91287
rect 126886 91216 126942 91225
rect 126886 91151 126942 91160
rect 129646 91216 129702 91225
rect 129646 91151 129702 91160
rect 126796 84108 126848 84114
rect 126796 84050 126848 84056
rect 125416 77240 125468 77246
rect 125416 77182 125468 77188
rect 126900 71670 126928 91151
rect 126888 71664 126940 71670
rect 126888 71606 126940 71612
rect 126886 69728 126942 69737
rect 126886 69663 126942 69672
rect 124128 63436 124180 63442
rect 124128 63378 124180 63384
rect 123484 56568 123536 56574
rect 123484 56510 123536 56516
rect 125508 25560 125560 25566
rect 125508 25502 125560 25508
rect 125520 3534 125548 25502
rect 126244 15972 126296 15978
rect 126244 15914 126296 15920
rect 126256 3602 126284 15914
rect 126244 3596 126296 3602
rect 126244 3538 126296 3544
rect 126900 3534 126928 69663
rect 129660 48278 129688 91151
rect 130764 89593 130792 91695
rect 151542 91352 151598 91361
rect 151542 91287 151598 91296
rect 132406 91216 132462 91225
rect 132406 91151 132462 91160
rect 135166 91216 135222 91225
rect 135166 91151 135222 91160
rect 136546 91216 136602 91225
rect 136546 91151 136602 91160
rect 130750 89584 130806 89593
rect 130750 89519 130806 89528
rect 132420 78577 132448 91151
rect 132868 91112 132920 91118
rect 132868 91054 132920 91060
rect 132880 86737 132908 91054
rect 132866 86728 132922 86737
rect 132866 86663 132922 86672
rect 135180 81326 135208 91151
rect 135168 81320 135220 81326
rect 135168 81262 135220 81268
rect 132406 78568 132462 78577
rect 132406 78503 132462 78512
rect 136560 50998 136588 91151
rect 151556 66162 151584 91287
rect 151648 89622 151676 91695
rect 151726 91216 151782 91225
rect 151726 91151 151782 91160
rect 153106 91216 153162 91225
rect 153106 91151 153162 91160
rect 151636 89616 151688 89622
rect 151636 89558 151688 89564
rect 151740 85474 151768 91151
rect 151728 85468 151780 85474
rect 151728 85410 151780 85416
rect 153120 82754 153148 91151
rect 153108 82748 153160 82754
rect 153108 82690 153160 82696
rect 160756 81326 160784 94415
rect 162490 93392 162546 93401
rect 162490 93327 162546 93336
rect 162122 93256 162178 93265
rect 162122 93191 162178 93200
rect 160744 81320 160796 81326
rect 160744 81262 160796 81268
rect 151544 66156 151596 66162
rect 151544 66098 151596 66104
rect 147034 64288 147090 64297
rect 147034 64223 147090 64232
rect 146944 53168 146996 53174
rect 146944 53110 146996 53116
rect 136548 50992 136600 50998
rect 136548 50934 136600 50940
rect 135260 50380 135312 50386
rect 135260 50322 135312 50328
rect 129648 48272 129700 48278
rect 129648 48214 129700 48220
rect 133144 47592 133196 47598
rect 133144 47534 133196 47540
rect 133156 20058 133184 47534
rect 133144 20052 133196 20058
rect 133144 19994 133196 20000
rect 130382 19952 130438 19961
rect 130382 19887 130438 19896
rect 130396 3534 130424 19887
rect 135272 11830 135300 50322
rect 144826 40624 144882 40633
rect 144826 40559 144882 40568
rect 141422 28248 141478 28257
rect 141422 28183 141478 28192
rect 135260 11824 135312 11830
rect 135260 11766 135312 11772
rect 136456 11824 136508 11830
rect 136456 11766 136508 11772
rect 132958 6216 133014 6225
rect 132958 6151 133014 6160
rect 124680 3528 124732 3534
rect 124680 3470 124732 3476
rect 125508 3528 125560 3534
rect 125508 3470 125560 3476
rect 125876 3528 125928 3534
rect 125876 3470 125928 3476
rect 126888 3528 126940 3534
rect 126888 3470 126940 3476
rect 129372 3528 129424 3534
rect 129372 3470 129424 3476
rect 130384 3528 130436 3534
rect 130384 3470 130436 3476
rect 121090 3431 121146 3440
rect 122288 3460 122340 3466
rect 121104 480 121132 3431
rect 122288 3402 122340 3408
rect 122748 3460 122800 3466
rect 122748 3402 122800 3408
rect 123484 3460 123536 3466
rect 123484 3402 123536 3408
rect 122300 480 122328 3402
rect 123496 480 123524 3402
rect 124692 480 124720 3470
rect 125888 480 125916 3470
rect 129384 480 129412 3470
rect 132972 480 133000 6151
rect 136468 480 136496 11766
rect 141436 3534 141464 28183
rect 144840 3534 144868 40559
rect 146956 8974 146984 53110
rect 147048 42158 147076 64223
rect 162136 63510 162164 93191
rect 162214 89040 162270 89049
rect 162214 88975 162270 88984
rect 162228 82521 162256 88975
rect 162504 85241 162532 93327
rect 162490 85232 162546 85241
rect 162490 85167 162546 85176
rect 164896 84114 164924 113766
rect 164976 100020 165028 100026
rect 164976 99962 165028 99968
rect 164884 84108 164936 84114
rect 164884 84050 164936 84056
rect 162214 82512 162270 82521
rect 162214 82447 162270 82456
rect 164988 77178 165016 99962
rect 165068 99884 165120 99890
rect 165068 99826 165120 99832
rect 165080 92177 165108 99826
rect 166276 93226 166304 124170
rect 166356 120148 166408 120154
rect 166356 120090 166408 120096
rect 166264 93220 166316 93226
rect 166264 93162 166316 93168
rect 166368 93129 166396 120090
rect 166540 111852 166592 111858
rect 166540 111794 166592 111800
rect 166448 106344 166500 106350
rect 166448 106286 166500 106292
rect 166354 93120 166410 93129
rect 166354 93055 166410 93064
rect 165066 92168 165122 92177
rect 165066 92103 165122 92112
rect 166460 85377 166488 106286
rect 166552 93906 166580 111794
rect 166540 93900 166592 93906
rect 166540 93842 166592 93848
rect 166446 85368 166502 85377
rect 166446 85303 166502 85312
rect 164976 77172 165028 77178
rect 164976 77114 165028 77120
rect 162124 63504 162176 63510
rect 162124 63446 162176 63452
rect 147036 42152 147088 42158
rect 147036 42094 147088 42100
rect 147128 42152 147180 42158
rect 147128 42094 147180 42100
rect 147140 28286 147168 42094
rect 160744 28416 160796 28422
rect 160744 28358 160796 28364
rect 147128 28280 147180 28286
rect 147128 28222 147180 28228
rect 160756 13190 160784 28358
rect 160744 13184 160796 13190
rect 160744 13126 160796 13132
rect 146944 8968 146996 8974
rect 146944 8910 146996 8916
rect 167012 6225 167040 318679
rect 167748 306374 167776 341527
rect 167840 331974 167868 351154
rect 168286 345672 168342 345681
rect 168286 345607 168342 345616
rect 167828 331968 167880 331974
rect 167828 331910 167880 331916
rect 167920 330608 167972 330614
rect 167920 330550 167972 330556
rect 167932 318170 167960 330550
rect 167920 318164 167972 318170
rect 167920 318106 167972 318112
rect 167828 318096 167880 318102
rect 167828 318038 167880 318044
rect 167656 306346 167776 306374
rect 167656 303657 167684 306346
rect 167642 303648 167698 303657
rect 167642 303583 167698 303592
rect 167656 280129 167684 303583
rect 167840 297498 167868 318038
rect 168300 315994 168328 345607
rect 168288 315988 168340 315994
rect 168288 315930 168340 315936
rect 168300 315382 168328 315930
rect 168288 315376 168340 315382
rect 168288 315318 168340 315324
rect 168286 298072 168342 298081
rect 168286 298007 168342 298016
rect 167828 297492 167880 297498
rect 167828 297434 167880 297440
rect 168300 296750 168328 298007
rect 168288 296744 168340 296750
rect 168288 296686 168340 296692
rect 167642 280120 167698 280129
rect 167642 280055 167698 280064
rect 167644 277432 167696 277438
rect 167644 277374 167696 277380
rect 167656 262857 167684 277374
rect 167736 265668 167788 265674
rect 167736 265610 167788 265616
rect 167642 262848 167698 262857
rect 167642 262783 167698 262792
rect 167090 261760 167146 261769
rect 167090 261695 167146 261704
rect 167104 260914 167132 261695
rect 167092 260908 167144 260914
rect 167092 260850 167144 260856
rect 167104 254561 167132 260850
rect 167090 254552 167146 254561
rect 167090 254487 167146 254496
rect 167642 251832 167698 251841
rect 167642 251767 167698 251776
rect 167656 235958 167684 251767
rect 167748 250510 167776 265610
rect 167736 250504 167788 250510
rect 167736 250446 167788 250452
rect 168194 249112 168250 249121
rect 168194 249047 168250 249056
rect 168208 242865 168236 249047
rect 168194 242856 168250 242865
rect 168194 242791 168250 242800
rect 167644 235952 167696 235958
rect 167644 235894 167696 235900
rect 168300 235793 168328 296686
rect 168392 242185 168420 390526
rect 168484 298081 168512 444479
rect 169760 443692 169812 443698
rect 169760 443634 169812 443640
rect 168562 370560 168618 370569
rect 168562 370495 168618 370504
rect 168470 298072 168526 298081
rect 168470 298007 168526 298016
rect 168576 279818 168604 370495
rect 169576 347064 169628 347070
rect 169576 347006 169628 347012
rect 169588 346633 169616 347006
rect 169574 346624 169630 346633
rect 169574 346559 169630 346568
rect 169588 345014 169616 346559
rect 169588 344986 169708 345014
rect 169024 289128 169076 289134
rect 169024 289070 169076 289076
rect 168564 279812 168616 279818
rect 168564 279754 168616 279760
rect 168378 242176 168434 242185
rect 168378 242111 168434 242120
rect 168286 235784 168342 235793
rect 168286 235719 168342 235728
rect 168286 235240 168342 235249
rect 168286 235175 168342 235184
rect 168300 201482 168328 235175
rect 169036 217569 169064 289070
rect 169574 278216 169630 278225
rect 169574 278151 169630 278160
rect 169022 217560 169078 217569
rect 169022 217495 169078 217504
rect 168380 215212 168432 215218
rect 168380 215154 168432 215160
rect 168392 214606 168420 215154
rect 169588 214606 169616 278151
rect 169680 269249 169708 344986
rect 169772 301617 169800 443634
rect 170416 317393 170444 527711
rect 170508 420918 170536 535502
rect 170496 420912 170548 420918
rect 170496 420854 170548 420860
rect 171048 394732 171100 394738
rect 171048 394674 171100 394680
rect 171060 356114 171088 394674
rect 171796 362982 171824 538902
rect 173254 535664 173310 535673
rect 173254 535599 173310 535608
rect 173164 502988 173216 502994
rect 173164 502930 173216 502936
rect 171874 449984 171930 449993
rect 171874 449919 171930 449928
rect 171784 362976 171836 362982
rect 171784 362918 171836 362924
rect 170496 356108 170548 356114
rect 170496 356050 170548 356056
rect 170588 356108 170640 356114
rect 170588 356050 170640 356056
rect 171048 356108 171100 356114
rect 171048 356050 171100 356056
rect 170508 325038 170536 356050
rect 170600 355473 170628 356050
rect 170586 355464 170642 355473
rect 170586 355399 170642 355408
rect 171784 354000 171836 354006
rect 171784 353942 171836 353948
rect 170588 353388 170640 353394
rect 170588 353330 170640 353336
rect 170496 325032 170548 325038
rect 170496 324974 170548 324980
rect 170496 320612 170548 320618
rect 170496 320554 170548 320560
rect 170402 317384 170458 317393
rect 170402 317319 170458 317328
rect 170404 306400 170456 306406
rect 170404 306342 170456 306348
rect 169758 301608 169814 301617
rect 169758 301543 169814 301552
rect 170416 279546 170444 306342
rect 170404 279540 170456 279546
rect 170404 279482 170456 279488
rect 169666 269240 169722 269249
rect 169666 269175 169722 269184
rect 170402 269240 170458 269249
rect 170402 269175 170458 269184
rect 168380 214600 168432 214606
rect 168380 214542 168432 214548
rect 169576 214600 169628 214606
rect 169576 214542 169628 214548
rect 170416 213217 170444 269175
rect 170508 255513 170536 320554
rect 170600 318102 170628 353330
rect 171140 325712 171192 325718
rect 171140 325654 171192 325660
rect 171152 319462 171180 325654
rect 171140 319456 171192 319462
rect 171140 319398 171192 319404
rect 170588 318096 170640 318102
rect 170588 318038 170640 318044
rect 171046 312488 171102 312497
rect 171046 312423 171102 312432
rect 170588 283620 170640 283626
rect 170588 283562 170640 283568
rect 170600 269074 170628 283562
rect 170588 269068 170640 269074
rect 170588 269010 170640 269016
rect 170862 267064 170918 267073
rect 170862 266999 170918 267008
rect 170876 266393 170904 266999
rect 170862 266384 170918 266393
rect 170862 266319 170918 266328
rect 170588 264240 170640 264246
rect 170588 264182 170640 264188
rect 170494 255504 170550 255513
rect 170494 255439 170550 255448
rect 170600 240854 170628 264182
rect 170588 240848 170640 240854
rect 170588 240790 170640 240796
rect 170402 213208 170458 213217
rect 170402 213143 170458 213152
rect 168288 201476 168340 201482
rect 168288 201418 168340 201424
rect 168300 198694 168328 201418
rect 169022 200696 169078 200705
rect 169022 200631 169078 200640
rect 168288 198688 168340 198694
rect 168288 198630 168340 198636
rect 167642 185192 167698 185201
rect 167642 185127 167698 185136
rect 167656 160070 167684 185127
rect 167734 175536 167790 175545
rect 167734 175471 167790 175480
rect 167748 165753 167776 175471
rect 167826 171592 167882 171601
rect 167826 171527 167882 171536
rect 167734 165744 167790 165753
rect 167734 165679 167790 165688
rect 167840 163538 167868 171527
rect 167828 163532 167880 163538
rect 167828 163474 167880 163480
rect 167644 160064 167696 160070
rect 167644 160006 167696 160012
rect 169036 146946 169064 200631
rect 170496 190528 170548 190534
rect 170496 190470 170548 190476
rect 169208 185020 169260 185026
rect 169208 184962 169260 184968
rect 169114 183696 169170 183705
rect 169114 183631 169170 183640
rect 169128 157350 169156 183631
rect 169220 173874 169248 184962
rect 170402 179480 170458 179489
rect 170402 179415 170458 179424
rect 169208 173868 169260 173874
rect 169208 173810 169260 173816
rect 169116 157344 169168 157350
rect 169116 157286 169168 157292
rect 170416 155922 170444 179415
rect 170508 167006 170536 190470
rect 170876 185609 170904 266319
rect 171060 265033 171088 312423
rect 171046 265024 171102 265033
rect 171046 264959 171102 264968
rect 170954 255368 171010 255377
rect 170954 255303 171010 255312
rect 170968 219201 170996 255303
rect 171796 244934 171824 353942
rect 171888 349897 171916 449919
rect 172428 430636 172480 430642
rect 172428 430578 172480 430584
rect 172440 376038 172468 430578
rect 173176 383654 173204 502930
rect 173268 430642 173296 535599
rect 173256 430636 173308 430642
rect 173256 430578 173308 430584
rect 173808 384328 173860 384334
rect 173808 384270 173860 384276
rect 173176 383626 173296 383654
rect 172428 376032 172480 376038
rect 172428 375974 172480 375980
rect 172060 372700 172112 372706
rect 172060 372642 172112 372648
rect 171968 362976 172020 362982
rect 171968 362918 172020 362924
rect 171874 349888 171930 349897
rect 171874 349823 171930 349832
rect 171980 311137 172008 362918
rect 172072 326369 172100 372642
rect 173268 369918 173296 383626
rect 173820 382401 173848 384270
rect 173806 382392 173862 382401
rect 173806 382327 173862 382336
rect 173256 369912 173308 369918
rect 173256 369854 173308 369860
rect 172518 356824 172574 356833
rect 172518 356759 172574 356768
rect 172426 338464 172482 338473
rect 172426 338399 172482 338408
rect 172058 326360 172114 326369
rect 172058 326295 172114 326304
rect 171966 311128 172022 311137
rect 171966 311063 172022 311072
rect 171968 309800 172020 309806
rect 171968 309742 172020 309748
rect 171876 286000 171928 286006
rect 171876 285942 171928 285948
rect 171784 244928 171836 244934
rect 171784 244870 171836 244876
rect 171796 224369 171824 244870
rect 171888 240854 171916 285942
rect 171980 285734 172008 309742
rect 172060 286340 172112 286346
rect 172060 286282 172112 286288
rect 171968 285728 172020 285734
rect 171968 285670 172020 285676
rect 171966 268424 172022 268433
rect 171966 268359 172022 268368
rect 171876 240848 171928 240854
rect 171876 240790 171928 240796
rect 171980 224641 172008 268359
rect 172072 266354 172100 286282
rect 172440 269074 172468 338399
rect 172532 276010 172560 356759
rect 173162 339688 173218 339697
rect 173162 339623 173218 339632
rect 172520 276004 172572 276010
rect 172520 275946 172572 275952
rect 172428 269068 172480 269074
rect 172428 269010 172480 269016
rect 172060 266348 172112 266354
rect 172060 266290 172112 266296
rect 172428 262880 172480 262886
rect 172428 262822 172480 262828
rect 171966 224632 172022 224641
rect 171966 224567 172022 224576
rect 171782 224360 171838 224369
rect 171782 224295 171838 224304
rect 170954 219192 171010 219201
rect 170954 219127 171010 219136
rect 172440 204921 172468 262822
rect 173176 231713 173204 339623
rect 173268 325694 173296 369854
rect 173268 325666 173756 325694
rect 173728 321609 173756 325666
rect 173714 321600 173770 321609
rect 173714 321535 173770 321544
rect 173254 313304 173310 313313
rect 173254 313239 173310 313248
rect 173268 299470 173296 313239
rect 173256 299464 173308 299470
rect 173256 299406 173308 299412
rect 173256 284368 173308 284374
rect 173256 284310 173308 284316
rect 173268 231810 173296 284310
rect 173728 276185 173756 321535
rect 173820 313313 173848 382327
rect 174556 360505 174584 569910
rect 177948 568608 178000 568614
rect 177948 568550 178000 568556
rect 177856 547936 177908 547942
rect 177856 547878 177908 547884
rect 177302 537024 177358 537033
rect 177302 536959 177358 536968
rect 174636 445800 174688 445806
rect 174636 445742 174688 445748
rect 174542 360496 174598 360505
rect 174542 360431 174598 360440
rect 174648 344457 174676 445742
rect 177316 429146 177344 536959
rect 177304 429140 177356 429146
rect 177304 429082 177356 429088
rect 176200 418192 176252 418198
rect 176200 418134 176252 418140
rect 176106 376816 176162 376825
rect 176106 376751 176162 376760
rect 174726 360496 174782 360505
rect 174726 360431 174782 360440
rect 174634 344448 174690 344457
rect 174634 344383 174690 344392
rect 174544 336864 174596 336870
rect 174544 336806 174596 336812
rect 173806 313304 173862 313313
rect 173806 313239 173862 313248
rect 173714 276176 173770 276185
rect 173714 276111 173770 276120
rect 173348 273284 173400 273290
rect 173348 273226 173400 273232
rect 173360 250510 173388 273226
rect 173808 255332 173860 255338
rect 173808 255274 173860 255280
rect 173440 252000 173492 252006
rect 173440 251942 173492 251948
rect 173348 250504 173400 250510
rect 173348 250446 173400 250452
rect 173452 240553 173480 251942
rect 173820 251938 173848 255274
rect 173808 251932 173860 251938
rect 173808 251874 173860 251880
rect 173438 240544 173494 240553
rect 173438 240479 173494 240488
rect 173256 231804 173308 231810
rect 173256 231746 173308 231752
rect 173162 231704 173218 231713
rect 173162 231639 173218 231648
rect 172426 204912 172482 204921
rect 172426 204847 172482 204856
rect 171784 203584 171836 203590
rect 171784 203526 171836 203532
rect 170862 185600 170918 185609
rect 170862 185535 170918 185544
rect 170588 178152 170640 178158
rect 170588 178094 170640 178100
rect 170496 167000 170548 167006
rect 170496 166942 170548 166948
rect 170600 165578 170628 178094
rect 170588 165572 170640 165578
rect 170588 165514 170640 165520
rect 170404 155916 170456 155922
rect 170404 155858 170456 155864
rect 169024 146940 169076 146946
rect 169024 146882 169076 146888
rect 169116 146328 169168 146334
rect 169116 146270 169168 146276
rect 167736 129056 167788 129062
rect 167736 128998 167788 129004
rect 167644 123480 167696 123486
rect 167644 123422 167696 123428
rect 167656 111761 167684 123422
rect 167642 111752 167698 111761
rect 167642 111687 167698 111696
rect 167748 110129 167776 128998
rect 169024 126268 169076 126274
rect 169024 126210 169076 126216
rect 167734 110120 167790 110129
rect 167734 110055 167790 110064
rect 167644 109064 167696 109070
rect 167644 109006 167696 109012
rect 167552 108996 167604 109002
rect 167552 108938 167604 108944
rect 167564 108769 167592 108938
rect 167550 108760 167606 108769
rect 167550 108695 167606 108704
rect 167656 88097 167684 109006
rect 167736 104236 167788 104242
rect 167736 104178 167788 104184
rect 167748 89593 167776 104178
rect 167828 97300 167880 97306
rect 167828 97242 167880 97248
rect 167840 89622 167868 97242
rect 168378 90400 168434 90409
rect 168378 90335 168434 90344
rect 168392 89622 168420 90335
rect 167828 89616 167880 89622
rect 167734 89584 167790 89593
rect 167828 89558 167880 89564
rect 168380 89616 168432 89622
rect 168380 89558 168432 89564
rect 167734 89519 167790 89528
rect 167642 88088 167698 88097
rect 167642 88023 167698 88032
rect 169036 66162 169064 126210
rect 169128 92410 169156 146270
rect 170404 144220 170456 144226
rect 170404 144162 170456 144168
rect 169208 114572 169260 114578
rect 169208 114514 169260 114520
rect 169116 92404 169168 92410
rect 169116 92346 169168 92352
rect 169220 79966 169248 114514
rect 169300 100768 169352 100774
rect 169300 100710 169352 100716
rect 169312 82657 169340 100710
rect 170416 94489 170444 144162
rect 170680 137284 170732 137290
rect 170680 137226 170732 137232
rect 170588 116000 170640 116006
rect 170588 115942 170640 115948
rect 170496 110492 170548 110498
rect 170496 110434 170548 110440
rect 170402 94480 170458 94489
rect 170402 94415 170458 94424
rect 170402 91760 170458 91769
rect 170402 91695 170458 91704
rect 169298 82648 169354 82657
rect 169298 82583 169354 82592
rect 169208 79960 169260 79966
rect 169208 79902 169260 79908
rect 169024 66156 169076 66162
rect 169024 66098 169076 66104
rect 166998 6216 167054 6225
rect 166998 6151 167054 6160
rect 140044 3528 140096 3534
rect 140044 3470 140096 3476
rect 141424 3528 141476 3534
rect 141424 3470 141476 3476
rect 143540 3528 143592 3534
rect 143540 3470 143592 3476
rect 144828 3528 144880 3534
rect 170416 3505 170444 91695
rect 170508 74458 170536 110434
rect 170600 88262 170628 115942
rect 170692 109002 170720 137226
rect 171796 133210 171824 203526
rect 173162 194168 173218 194177
rect 173162 194103 173218 194112
rect 171876 182232 171928 182238
rect 171876 182174 171928 182180
rect 171888 158710 171916 182174
rect 171876 158704 171928 158710
rect 171876 158646 171928 158652
rect 171876 143608 171928 143614
rect 171876 143550 171928 143556
rect 171784 133204 171836 133210
rect 171784 133146 171836 133152
rect 171784 121508 171836 121514
rect 171784 121450 171836 121456
rect 170680 108996 170732 109002
rect 170680 108938 170732 108944
rect 170772 107704 170824 107710
rect 170772 107646 170824 107652
rect 170784 93809 170812 107646
rect 170770 93800 170826 93809
rect 170770 93735 170826 93744
rect 171796 89690 171824 121450
rect 171888 99890 171916 143550
rect 173176 141438 173204 194103
rect 173268 172417 173296 231746
rect 174556 223582 174584 336806
rect 174634 316840 174690 316849
rect 174634 316775 174690 316784
rect 174648 241505 174676 316775
rect 174740 306374 174768 360431
rect 174820 355360 174872 355366
rect 174820 355302 174872 355308
rect 174832 309777 174860 355302
rect 176014 348120 176070 348129
rect 176014 348055 176070 348064
rect 174910 345128 174966 345137
rect 174910 345063 174966 345072
rect 174924 320958 174952 345063
rect 174912 320952 174964 320958
rect 174912 320894 174964 320900
rect 174818 309768 174874 309777
rect 174818 309703 174874 309712
rect 174740 306346 175136 306374
rect 175108 294001 175136 306346
rect 175188 304360 175240 304366
rect 175188 304302 175240 304308
rect 175200 303686 175228 304302
rect 175188 303680 175240 303686
rect 175188 303622 175240 303628
rect 175094 293992 175150 294001
rect 175094 293927 175150 293936
rect 175108 273222 175136 293927
rect 175096 273216 175148 273222
rect 175096 273158 175148 273164
rect 174726 271144 174782 271153
rect 174726 271079 174782 271088
rect 174740 258738 174768 271079
rect 174728 258732 174780 258738
rect 174728 258674 174780 258680
rect 175096 258596 175148 258602
rect 175096 258538 175148 258544
rect 174634 241496 174690 241505
rect 174634 241431 174690 241440
rect 174648 235142 174676 241431
rect 174636 235136 174688 235142
rect 174636 235078 174688 235084
rect 174544 223576 174596 223582
rect 174544 223518 174596 223524
rect 173808 209704 173860 209710
rect 173808 209646 173860 209652
rect 173820 208457 173848 209646
rect 173806 208448 173862 208457
rect 173806 208383 173862 208392
rect 174544 189100 174596 189106
rect 174544 189042 174596 189048
rect 173346 180840 173402 180849
rect 173346 180775 173402 180784
rect 173254 172408 173310 172417
rect 173254 172343 173310 172352
rect 173360 161362 173388 180775
rect 174556 168366 174584 189042
rect 175108 182073 175136 258538
rect 175094 182064 175150 182073
rect 175094 181999 175150 182008
rect 175108 181393 175136 181999
rect 175094 181384 175150 181393
rect 175094 181319 175150 181328
rect 174544 168360 174596 168366
rect 174544 168302 174596 168308
rect 173348 161356 173400 161362
rect 173348 161298 173400 161304
rect 173256 142180 173308 142186
rect 173256 142122 173308 142128
rect 173164 141432 173216 141438
rect 173164 141374 173216 141380
rect 173164 117972 173216 117978
rect 173164 117914 173216 117920
rect 171968 104168 172020 104174
rect 171968 104110 172020 104116
rect 171876 99884 171928 99890
rect 171876 99826 171928 99832
rect 171876 91860 171928 91866
rect 171876 91802 171928 91808
rect 171784 89684 171836 89690
rect 171784 89626 171836 89632
rect 170588 88256 170640 88262
rect 170588 88198 170640 88204
rect 170496 74452 170548 74458
rect 170496 74394 170548 74400
rect 171888 70378 171916 91802
rect 171980 85474 172008 104110
rect 172060 99408 172112 99414
rect 172060 99350 172112 99356
rect 172072 86970 172100 99350
rect 172060 86964 172112 86970
rect 172060 86906 172112 86912
rect 171968 85468 172020 85474
rect 171968 85410 172020 85416
rect 173176 71670 173204 117914
rect 173268 92478 173296 142122
rect 174544 139460 174596 139466
rect 174544 139402 174596 139408
rect 173348 127628 173400 127634
rect 173348 127570 173400 127576
rect 173256 92472 173308 92478
rect 173256 92414 173308 92420
rect 173360 92313 173388 127570
rect 173440 105596 173492 105602
rect 173440 105538 173492 105544
rect 173346 92304 173402 92313
rect 173346 92239 173402 92248
rect 173452 78674 173480 105538
rect 174556 94081 174584 139402
rect 174636 118720 174688 118726
rect 174636 118662 174688 118668
rect 174542 94072 174598 94081
rect 174542 94007 174598 94016
rect 174648 91050 174676 118662
rect 174726 97064 174782 97073
rect 174726 96999 174782 97008
rect 174636 91044 174688 91050
rect 174636 90986 174688 90992
rect 173440 78668 173492 78674
rect 173440 78610 173492 78616
rect 174740 74526 174768 96999
rect 174728 74520 174780 74526
rect 174728 74462 174780 74468
rect 173164 71664 173216 71670
rect 173164 71606 173216 71612
rect 171876 70372 171928 70378
rect 171876 70314 171928 70320
rect 175200 10305 175228 303622
rect 175924 248532 175976 248538
rect 175924 248474 175976 248480
rect 175936 234433 175964 248474
rect 175922 234424 175978 234433
rect 175922 234359 175978 234368
rect 175936 173913 175964 234359
rect 176028 217977 176056 348055
rect 176120 337618 176148 376751
rect 176108 337612 176160 337618
rect 176108 337554 176160 337560
rect 176108 331288 176160 331294
rect 176108 331230 176160 331236
rect 176120 323785 176148 331230
rect 176106 323776 176162 323785
rect 176106 323711 176162 323720
rect 176108 288448 176160 288454
rect 176108 288390 176160 288396
rect 176120 274650 176148 288390
rect 176108 274644 176160 274650
rect 176108 274586 176160 274592
rect 176108 272332 176160 272338
rect 176108 272274 176160 272280
rect 176120 258602 176148 272274
rect 176108 258596 176160 258602
rect 176108 258538 176160 258544
rect 176108 252680 176160 252686
rect 176108 252622 176160 252628
rect 176120 233918 176148 252622
rect 176212 246430 176240 418134
rect 177396 393984 177448 393990
rect 177396 393926 177448 393932
rect 177304 382968 177356 382974
rect 177304 382910 177356 382916
rect 176658 349888 176714 349897
rect 176658 349823 176714 349832
rect 176672 309913 176700 349823
rect 176658 309904 176714 309913
rect 176658 309839 176714 309848
rect 177316 307737 177344 382910
rect 177408 380186 177436 393926
rect 177396 380180 177448 380186
rect 177396 380122 177448 380128
rect 177394 363624 177450 363633
rect 177394 363559 177450 363568
rect 177302 307728 177358 307737
rect 177302 307663 177358 307672
rect 177408 295322 177436 363559
rect 177868 353977 177896 547878
rect 177960 363798 177988 568550
rect 191104 563100 191156 563106
rect 191104 563042 191156 563048
rect 186964 561740 187016 561746
rect 186964 561682 187016 561688
rect 178684 560380 178736 560386
rect 178684 560322 178736 560328
rect 178696 529922 178724 560322
rect 180156 556300 180208 556306
rect 180156 556242 180208 556248
rect 178776 536852 178828 536858
rect 178776 536794 178828 536800
rect 178684 529916 178736 529922
rect 178684 529858 178736 529864
rect 178684 495508 178736 495514
rect 178684 495450 178736 495456
rect 178040 400988 178092 400994
rect 178040 400930 178092 400936
rect 178052 379409 178080 400930
rect 178038 379400 178094 379409
rect 178038 379335 178094 379344
rect 178406 379400 178462 379409
rect 178406 379335 178462 379344
rect 178420 378729 178448 379335
rect 178406 378720 178462 378729
rect 178406 378655 178462 378664
rect 177948 363792 178000 363798
rect 177948 363734 178000 363740
rect 177960 363662 177988 363734
rect 177948 363656 178000 363662
rect 177948 363598 178000 363604
rect 178696 359553 178724 495450
rect 178788 421598 178816 536794
rect 180064 530664 180116 530670
rect 180064 530606 180116 530612
rect 179420 460964 179472 460970
rect 179420 460906 179472 460912
rect 179328 433356 179380 433362
rect 179328 433298 179380 433304
rect 178776 421592 178828 421598
rect 178776 421534 178828 421540
rect 178866 375456 178922 375465
rect 178866 375391 178922 375400
rect 178774 366480 178830 366489
rect 178774 366415 178830 366424
rect 178682 359544 178738 359553
rect 178682 359479 178738 359488
rect 177854 353968 177910 353977
rect 177854 353903 177910 353912
rect 177868 353569 177896 353903
rect 177854 353560 177910 353569
rect 177854 353495 177910 353504
rect 178682 336968 178738 336977
rect 178682 336903 178738 336912
rect 177486 335608 177542 335617
rect 177486 335543 177542 335552
rect 177500 315314 177528 335543
rect 177488 315308 177540 315314
rect 177488 315250 177540 315256
rect 177488 309868 177540 309874
rect 177488 309810 177540 309816
rect 177396 295316 177448 295322
rect 177396 295258 177448 295264
rect 177304 294092 177356 294098
rect 177304 294034 177356 294040
rect 176660 282192 176712 282198
rect 176660 282134 176712 282140
rect 176672 281586 176700 282134
rect 176660 281580 176712 281586
rect 176660 281522 176712 281528
rect 177316 264246 177344 294034
rect 177396 275324 177448 275330
rect 177396 275266 177448 275272
rect 177304 264240 177356 264246
rect 177304 264182 177356 264188
rect 176200 246424 176252 246430
rect 176200 246366 176252 246372
rect 177304 244316 177356 244322
rect 177304 244258 177356 244264
rect 177316 236774 177344 244258
rect 177304 236768 177356 236774
rect 177304 236710 177356 236716
rect 177304 235136 177356 235142
rect 177304 235078 177356 235084
rect 176108 233912 176160 233918
rect 176108 233854 176160 233860
rect 176014 217968 176070 217977
rect 176014 217903 176070 217912
rect 176016 195356 176068 195362
rect 176016 195298 176068 195304
rect 175922 173904 175978 173913
rect 175922 173839 175978 173848
rect 175924 163532 175976 163538
rect 175924 163474 175976 163480
rect 175936 150414 175964 163474
rect 175924 150408 175976 150414
rect 175924 150350 175976 150356
rect 175924 138032 175976 138038
rect 175924 137974 175976 137980
rect 175936 89049 175964 137974
rect 176028 137465 176056 195298
rect 176106 178120 176162 178129
rect 176106 178055 176162 178064
rect 176120 164218 176148 178055
rect 176108 164212 176160 164218
rect 176108 164154 176160 164160
rect 176014 137456 176070 137465
rect 176014 137391 176070 137400
rect 176016 122868 176068 122874
rect 176016 122810 176068 122816
rect 176028 93974 176056 122810
rect 176108 100836 176160 100842
rect 176108 100778 176160 100784
rect 176016 93968 176068 93974
rect 176016 93910 176068 93916
rect 175922 89040 175978 89049
rect 175922 88975 175978 88984
rect 176120 80034 176148 100778
rect 176200 94512 176252 94518
rect 176200 94454 176252 94460
rect 176108 80028 176160 80034
rect 176108 79970 176160 79976
rect 176212 77246 176240 94454
rect 176200 77240 176252 77246
rect 176200 77182 176252 77188
rect 175186 10296 175242 10305
rect 175186 10231 175242 10240
rect 177316 4049 177344 235078
rect 177408 229770 177436 275266
rect 177500 247625 177528 309810
rect 177578 307728 177634 307737
rect 177578 307663 177634 307672
rect 177592 307057 177620 307663
rect 177578 307048 177634 307057
rect 177578 306983 177634 306992
rect 177592 284986 177620 306983
rect 177580 284980 177632 284986
rect 177580 284922 177632 284928
rect 177948 281580 178000 281586
rect 177948 281522 178000 281528
rect 177486 247616 177542 247625
rect 177486 247551 177542 247560
rect 177488 242276 177540 242282
rect 177488 242218 177540 242224
rect 177396 229764 177448 229770
rect 177396 229706 177448 229712
rect 177500 227050 177528 242218
rect 177488 227044 177540 227050
rect 177488 226986 177540 226992
rect 177762 202872 177818 202881
rect 177762 202807 177764 202816
rect 177816 202807 177818 202816
rect 177764 202778 177816 202784
rect 177856 199436 177908 199442
rect 177856 199378 177908 199384
rect 177394 198248 177450 198257
rect 177394 198183 177450 198192
rect 177408 118046 177436 198183
rect 177868 195362 177896 199378
rect 177856 195356 177908 195362
rect 177856 195298 177908 195304
rect 177580 188352 177632 188358
rect 177580 188294 177632 188300
rect 177488 178084 177540 178090
rect 177488 178026 177540 178032
rect 177500 164150 177528 178026
rect 177592 177313 177620 188294
rect 177960 178702 177988 281522
rect 178696 272338 178724 336903
rect 178684 272332 178736 272338
rect 178684 272274 178736 272280
rect 178684 269068 178736 269074
rect 178684 269010 178736 269016
rect 178040 256692 178092 256698
rect 178040 256634 178092 256640
rect 178052 256018 178080 256634
rect 178040 256012 178092 256018
rect 178040 255954 178092 255960
rect 178038 228440 178094 228449
rect 178038 228375 178040 228384
rect 178092 228375 178094 228384
rect 178040 228346 178092 228352
rect 177948 178696 178000 178702
rect 177948 178638 178000 178644
rect 177578 177304 177634 177313
rect 177578 177239 177634 177248
rect 177488 164144 177540 164150
rect 177488 164086 177540 164092
rect 177488 135312 177540 135318
rect 177488 135254 177540 135260
rect 177396 118040 177448 118046
rect 177396 117982 177448 117988
rect 177500 91633 177528 135254
rect 178696 134638 178724 269010
rect 178788 262206 178816 366415
rect 178880 336025 178908 375391
rect 178866 336016 178922 336025
rect 178866 335951 178922 335960
rect 178866 273320 178922 273329
rect 178866 273255 178922 273264
rect 178776 262200 178828 262206
rect 178776 262142 178828 262148
rect 178774 250472 178830 250481
rect 178774 250407 178830 250416
rect 178788 236065 178816 250407
rect 178774 236056 178830 236065
rect 178774 235991 178830 236000
rect 178776 200796 178828 200802
rect 178776 200738 178828 200744
rect 178788 138718 178816 200738
rect 178880 199442 178908 273255
rect 179340 256698 179368 433298
rect 179432 320113 179460 460906
rect 180076 350577 180104 530606
rect 180168 504422 180196 556242
rect 184846 554840 184902 554849
rect 184846 554775 184902 554784
rect 184296 552152 184348 552158
rect 184296 552094 184348 552100
rect 182916 550724 182968 550730
rect 182916 550666 182968 550672
rect 182822 533352 182878 533361
rect 182822 533287 182878 533296
rect 180156 504416 180208 504422
rect 180156 504358 180208 504364
rect 180156 483676 180208 483682
rect 180156 483618 180208 483624
rect 180168 392018 180196 483618
rect 182088 477556 182140 477562
rect 182088 477498 182140 477504
rect 181444 414044 181496 414050
rect 181444 413986 181496 413992
rect 180156 392012 180208 392018
rect 180156 391954 180208 391960
rect 180062 350568 180118 350577
rect 180062 350503 180118 350512
rect 180076 326466 180104 350503
rect 180064 326460 180116 326466
rect 180064 326402 180116 326408
rect 179418 320104 179474 320113
rect 179418 320039 179474 320048
rect 179420 279540 179472 279546
rect 179420 279482 179472 279488
rect 179432 278798 179460 279482
rect 179420 278792 179472 278798
rect 179420 278734 179472 278740
rect 179328 256692 179380 256698
rect 179328 256634 179380 256640
rect 180168 244934 180196 391954
rect 180430 331256 180486 331265
rect 180430 331191 180486 331200
rect 180246 320104 180302 320113
rect 180246 320039 180302 320048
rect 180260 318889 180288 320039
rect 180246 318880 180302 318889
rect 180246 318815 180302 318824
rect 180260 298858 180288 318815
rect 180248 298852 180300 298858
rect 180248 298794 180300 298800
rect 180248 297492 180300 297498
rect 180248 297434 180300 297440
rect 180260 272542 180288 297434
rect 180248 272536 180300 272542
rect 180248 272478 180300 272484
rect 180156 244928 180208 244934
rect 180156 244870 180208 244876
rect 179418 241360 179474 241369
rect 179418 241295 179474 241304
rect 179432 240786 179460 241295
rect 179420 240780 179472 240786
rect 179420 240722 179472 240728
rect 178958 236056 179014 236065
rect 178958 235991 179014 236000
rect 178868 199436 178920 199442
rect 178868 199378 178920 199384
rect 178972 198694 179000 235991
rect 180062 231840 180118 231849
rect 180062 231775 180118 231784
rect 180076 230518 180104 231775
rect 180064 230512 180116 230518
rect 180064 230454 180116 230460
rect 178960 198688 179012 198694
rect 178960 198630 179012 198636
rect 180154 185056 180210 185065
rect 180154 184991 180210 185000
rect 178866 182200 178922 182209
rect 178866 182135 178922 182144
rect 178880 155854 178908 182135
rect 180168 157282 180196 184991
rect 180246 176896 180302 176905
rect 180246 176831 180302 176840
rect 180260 158642 180288 176831
rect 180248 158636 180300 158642
rect 180248 158578 180300 158584
rect 180156 157276 180208 157282
rect 180156 157218 180208 157224
rect 178868 155848 178920 155854
rect 178868 155790 178920 155796
rect 180340 150476 180392 150482
rect 180340 150418 180392 150424
rect 178776 138712 178828 138718
rect 178776 138654 178828 138660
rect 178684 134632 178736 134638
rect 178684 134574 178736 134580
rect 178776 131776 178828 131782
rect 178776 131718 178828 131724
rect 177580 113892 177632 113898
rect 177580 113834 177632 113840
rect 177486 91624 177542 91633
rect 177486 91559 177542 91568
rect 177396 84856 177448 84862
rect 177396 84798 177448 84804
rect 177302 4040 177358 4049
rect 177302 3975 177358 3984
rect 144828 3470 144880 3476
rect 170402 3496 170458 3505
rect 140056 480 140084 3470
rect 143552 480 143580 3470
rect 170402 3431 170458 3440
rect 177408 2009 177436 84798
rect 177592 75818 177620 113834
rect 177672 109132 177724 109138
rect 177672 109074 177724 109080
rect 177684 84182 177712 109074
rect 178684 104916 178736 104922
rect 178684 104858 178736 104864
rect 178040 91792 178092 91798
rect 178040 91734 178092 91740
rect 178052 86737 178080 91734
rect 178696 88233 178724 104858
rect 178682 88224 178738 88233
rect 178682 88159 178738 88168
rect 178038 86728 178094 86737
rect 178038 86663 178094 86672
rect 178682 86184 178738 86193
rect 178682 86119 178738 86128
rect 177672 84176 177724 84182
rect 177672 84118 177724 84124
rect 177580 75812 177632 75818
rect 177580 75754 177632 75760
rect 178696 28354 178724 86119
rect 178788 82754 178816 131718
rect 180248 131164 180300 131170
rect 180248 131106 180300 131112
rect 180156 130416 180208 130422
rect 180156 130358 180208 130364
rect 178868 95940 178920 95946
rect 178868 95882 178920 95888
rect 178776 82748 178828 82754
rect 178776 82690 178828 82696
rect 178880 67522 178908 95882
rect 178960 87712 179012 87718
rect 178960 87654 179012 87660
rect 178868 67516 178920 67522
rect 178868 67458 178920 67464
rect 178972 64802 179000 87654
rect 178960 64796 179012 64802
rect 178960 64738 179012 64744
rect 180168 50998 180196 130358
rect 180260 68950 180288 131106
rect 180352 123486 180380 150418
rect 180340 123480 180392 123486
rect 180340 123422 180392 123428
rect 180340 121576 180392 121582
rect 180340 121518 180392 121524
rect 180352 93158 180380 121518
rect 180340 93152 180392 93158
rect 180340 93094 180392 93100
rect 180248 68944 180300 68950
rect 180248 68886 180300 68892
rect 180156 50992 180208 50998
rect 180156 50934 180208 50940
rect 178684 28348 178736 28354
rect 178684 28290 178736 28296
rect 180444 9654 180472 331191
rect 181456 289134 181484 413986
rect 182100 369238 182128 477498
rect 182088 369232 182140 369238
rect 182088 369174 182140 369180
rect 181628 368552 181680 368558
rect 181628 368494 181680 368500
rect 181536 355360 181588 355366
rect 181536 355302 181588 355308
rect 181548 346390 181576 355302
rect 181640 354657 181668 368494
rect 181626 354648 181682 354657
rect 181626 354583 181682 354592
rect 181536 346384 181588 346390
rect 181536 346326 181588 346332
rect 181444 289128 181496 289134
rect 181444 289070 181496 289076
rect 181442 285016 181498 285025
rect 181442 284951 181498 284960
rect 180708 278792 180760 278798
rect 180708 278734 180760 278740
rect 180616 265736 180668 265742
rect 180616 265678 180668 265684
rect 180524 245608 180576 245614
rect 180524 245550 180576 245556
rect 180536 241369 180564 245550
rect 180522 241360 180578 241369
rect 180522 241295 180578 241304
rect 180628 231849 180656 265678
rect 180614 231840 180670 231849
rect 180614 231775 180670 231784
rect 180720 182850 180748 278734
rect 181456 265742 181484 284951
rect 181548 269074 181576 346326
rect 182836 336977 182864 533287
rect 182928 365838 182956 550666
rect 184202 539880 184258 539889
rect 184202 539815 184258 539824
rect 183560 454708 183612 454714
rect 183560 454650 183612 454656
rect 183098 369880 183154 369889
rect 183098 369815 183154 369824
rect 182916 365832 182968 365838
rect 182916 365774 182968 365780
rect 182822 336968 182878 336977
rect 182822 336903 182878 336912
rect 182180 329112 182232 329118
rect 182180 329054 182232 329060
rect 182192 312497 182220 329054
rect 182824 315376 182876 315382
rect 182824 315318 182876 315324
rect 182178 312488 182234 312497
rect 182178 312423 182234 312432
rect 181720 273964 181772 273970
rect 181720 273906 181772 273912
rect 181626 273456 181682 273465
rect 181626 273391 181682 273400
rect 181536 269068 181588 269074
rect 181536 269010 181588 269016
rect 181444 265736 181496 265742
rect 181444 265678 181496 265684
rect 181444 262268 181496 262274
rect 181444 262210 181496 262216
rect 180708 182844 180760 182850
rect 180708 182786 180760 182792
rect 181456 177342 181484 262210
rect 181536 249416 181588 249422
rect 181536 249358 181588 249364
rect 181548 223514 181576 249358
rect 181640 245614 181668 273391
rect 181732 248538 181760 273906
rect 182088 263628 182140 263634
rect 182088 263570 182140 263576
rect 182100 262274 182128 263570
rect 182088 262268 182140 262274
rect 182088 262210 182140 262216
rect 182088 259412 182140 259418
rect 182088 259354 182140 259360
rect 182100 258194 182128 259354
rect 182088 258188 182140 258194
rect 182088 258130 182140 258136
rect 181720 248532 181772 248538
rect 181720 248474 181772 248480
rect 181628 245608 181680 245614
rect 181628 245550 181680 245556
rect 181720 243024 181772 243030
rect 181720 242966 181772 242972
rect 181628 230512 181680 230518
rect 181628 230454 181680 230460
rect 181536 223508 181588 223514
rect 181536 223450 181588 223456
rect 181548 185638 181576 223450
rect 181640 200705 181668 230454
rect 181732 226302 181760 242966
rect 182100 235278 182128 258130
rect 182088 235272 182140 235278
rect 182088 235214 182140 235220
rect 181720 226296 181772 226302
rect 181720 226238 181772 226244
rect 182180 210452 182232 210458
rect 182180 210394 182232 210400
rect 182192 206825 182220 210394
rect 182178 206816 182234 206825
rect 182178 206751 182234 206760
rect 181626 200696 181682 200705
rect 181626 200631 181682 200640
rect 181628 196648 181680 196654
rect 181628 196590 181680 196596
rect 181536 185632 181588 185638
rect 181536 185574 181588 185580
rect 181640 177410 181668 196590
rect 181628 177404 181680 177410
rect 181628 177346 181680 177352
rect 181444 177336 181496 177342
rect 181444 177278 181496 177284
rect 181628 110560 181680 110566
rect 181628 110502 181680 110508
rect 181534 103864 181590 103873
rect 181534 103799 181590 103808
rect 181442 93120 181498 93129
rect 181442 93055 181498 93064
rect 181456 64297 181484 93055
rect 181548 84153 181576 103799
rect 181640 91089 181668 110502
rect 181626 91080 181682 91089
rect 181626 91015 181682 91024
rect 181534 84144 181590 84153
rect 181534 84079 181590 84088
rect 181442 64288 181498 64297
rect 181442 64223 181498 64232
rect 180432 9648 180484 9654
rect 180432 9590 180484 9596
rect 182836 6905 182864 315318
rect 182928 305697 182956 365774
rect 183008 337612 183060 337618
rect 183008 337554 183060 337560
rect 182914 305688 182970 305697
rect 182914 305623 182970 305632
rect 183020 283121 183048 337554
rect 183112 337414 183140 369815
rect 183192 342372 183244 342378
rect 183192 342314 183244 342320
rect 183100 337408 183152 337414
rect 183100 337350 183152 337356
rect 183204 316713 183232 342314
rect 183190 316704 183246 316713
rect 183190 316639 183246 316648
rect 183376 297492 183428 297498
rect 183376 297434 183428 297440
rect 183006 283112 183062 283121
rect 183006 283047 183062 283056
rect 183282 282976 183338 282985
rect 183282 282911 183338 282920
rect 183296 282878 183324 282911
rect 183284 282872 183336 282878
rect 183284 282814 183336 282820
rect 183284 276684 183336 276690
rect 183284 276626 183336 276632
rect 183296 276146 183324 276626
rect 183284 276140 183336 276146
rect 183284 276082 183336 276088
rect 183296 258074 183324 276082
rect 183204 258046 183324 258074
rect 183204 171057 183232 258046
rect 183284 251864 183336 251870
rect 183284 251806 183336 251812
rect 183296 231849 183324 251806
rect 183388 238678 183416 297434
rect 183466 287192 183522 287201
rect 183466 287127 183522 287136
rect 183480 274582 183508 287127
rect 183468 274576 183520 274582
rect 183468 274518 183520 274524
rect 183572 251870 183600 454650
rect 184216 267073 184244 539815
rect 184308 454714 184336 552094
rect 184296 454708 184348 454714
rect 184296 454650 184348 454656
rect 184860 447137 184888 554775
rect 185674 549400 185730 549409
rect 185674 549335 185730 549344
rect 185584 546508 185636 546514
rect 185584 546450 185636 546456
rect 185400 487824 185452 487830
rect 185400 487766 185452 487772
rect 185412 487218 185440 487766
rect 184940 487212 184992 487218
rect 184940 487154 184992 487160
rect 185400 487212 185452 487218
rect 185400 487154 185452 487160
rect 184846 447128 184902 447137
rect 184846 447063 184902 447072
rect 184388 384396 184440 384402
rect 184388 384338 184440 384344
rect 184296 376032 184348 376038
rect 184296 375974 184348 375980
rect 184308 345953 184336 375974
rect 184400 370569 184428 384338
rect 184386 370560 184442 370569
rect 184386 370495 184442 370504
rect 184294 345944 184350 345953
rect 184294 345879 184350 345888
rect 184294 340096 184350 340105
rect 184294 340031 184350 340040
rect 184308 318753 184336 340031
rect 184294 318744 184350 318753
rect 184294 318679 184350 318688
rect 184846 318744 184902 318753
rect 184846 318679 184902 318688
rect 184860 317529 184888 318679
rect 184846 317520 184902 317529
rect 184846 317455 184902 317464
rect 184296 304292 184348 304298
rect 184296 304234 184348 304240
rect 184308 273465 184336 304234
rect 184860 283257 184888 317455
rect 184846 283248 184902 283257
rect 184846 283183 184902 283192
rect 184386 283112 184442 283121
rect 184386 283047 184442 283056
rect 184294 273456 184350 273465
rect 184294 273391 184350 273400
rect 184400 270502 184428 283047
rect 184756 271176 184808 271182
rect 184756 271118 184808 271124
rect 184388 270496 184440 270502
rect 184388 270438 184440 270444
rect 184296 269068 184348 269074
rect 184296 269010 184348 269016
rect 184202 267064 184258 267073
rect 184202 266999 184258 267008
rect 184204 257372 184256 257378
rect 184204 257314 184256 257320
rect 184216 256766 184244 257314
rect 184204 256760 184256 256766
rect 184204 256702 184256 256708
rect 183560 251864 183612 251870
rect 183560 251806 183612 251812
rect 184204 246424 184256 246430
rect 184204 246366 184256 246372
rect 183376 238672 183428 238678
rect 183376 238614 183428 238620
rect 183388 238513 183416 238614
rect 183374 238504 183430 238513
rect 183374 238439 183430 238448
rect 183282 231840 183338 231849
rect 183282 231775 183338 231784
rect 183190 171048 183246 171057
rect 183190 170983 183246 170992
rect 182916 135380 182968 135386
rect 182916 135322 182968 135328
rect 182928 87961 182956 135322
rect 182914 87952 182970 87961
rect 182914 87887 182970 87896
rect 184216 7585 184244 246366
rect 184308 245857 184336 269010
rect 184664 256760 184716 256766
rect 184664 256702 184716 256708
rect 184294 245848 184350 245857
rect 184294 245783 184350 245792
rect 184676 230450 184704 256702
rect 184768 239737 184796 271118
rect 184846 247616 184902 247625
rect 184846 247551 184902 247560
rect 184754 239728 184810 239737
rect 184754 239663 184810 239672
rect 184768 238377 184796 239663
rect 184754 238368 184810 238377
rect 184754 238303 184810 238312
rect 184756 234660 184808 234666
rect 184756 234602 184808 234608
rect 184664 230444 184716 230450
rect 184664 230386 184716 230392
rect 184294 229800 184350 229809
rect 184294 229735 184350 229744
rect 184308 219434 184336 229735
rect 184296 219428 184348 219434
rect 184296 219370 184348 219376
rect 184664 204944 184716 204950
rect 184664 204886 184716 204892
rect 184676 191185 184704 204886
rect 184768 203658 184796 234602
rect 184756 203652 184808 203658
rect 184756 203594 184808 203600
rect 184662 191176 184718 191185
rect 184662 191111 184718 191120
rect 184860 151065 184888 247551
rect 184952 235249 184980 487154
rect 185596 383654 185624 546450
rect 185688 522986 185716 549335
rect 185676 522980 185728 522986
rect 185676 522922 185728 522928
rect 185596 383626 185716 383654
rect 185584 382288 185636 382294
rect 185584 382230 185636 382236
rect 185596 376009 185624 382230
rect 185688 376786 185716 383626
rect 185676 376780 185728 376786
rect 185676 376722 185728 376728
rect 185582 376000 185638 376009
rect 185582 375935 185638 375944
rect 185584 370524 185636 370530
rect 185584 370466 185636 370472
rect 185596 282169 185624 370466
rect 185688 327865 185716 376722
rect 186412 374672 186464 374678
rect 186412 374614 186464 374620
rect 186424 368490 186452 374614
rect 186412 368484 186464 368490
rect 186412 368426 186464 368432
rect 186976 358834 187004 561682
rect 188344 557592 188396 557598
rect 188344 557534 188396 557540
rect 187054 556200 187110 556209
rect 187054 556135 187110 556144
rect 187068 520946 187096 556135
rect 187148 550656 187200 550662
rect 187148 550598 187200 550604
rect 187160 528562 187188 550598
rect 187148 528556 187200 528562
rect 187148 528498 187200 528504
rect 187056 520940 187108 520946
rect 187056 520882 187108 520888
rect 187148 502376 187200 502382
rect 187148 502318 187200 502324
rect 187056 489932 187108 489938
rect 187056 489874 187108 489880
rect 186964 358828 187016 358834
rect 186964 358770 187016 358776
rect 186228 343664 186280 343670
rect 186228 343606 186280 343612
rect 185674 327856 185730 327865
rect 185674 327791 185730 327800
rect 186240 295361 186268 343606
rect 186976 329118 187004 358770
rect 186964 329112 187016 329118
rect 186964 329054 187016 329060
rect 186964 327752 187016 327758
rect 186964 327694 187016 327700
rect 186320 325032 186372 325038
rect 186320 324974 186372 324980
rect 186332 317422 186360 324974
rect 186320 317416 186372 317422
rect 186320 317358 186372 317364
rect 186226 295352 186282 295361
rect 186226 295287 186282 295296
rect 185676 284436 185728 284442
rect 185676 284378 185728 284384
rect 185582 282160 185638 282169
rect 185582 282095 185638 282104
rect 185032 274576 185084 274582
rect 185032 274518 185084 274524
rect 184938 235240 184994 235249
rect 184938 235175 184994 235184
rect 185044 234666 185072 274518
rect 185688 259418 185716 284378
rect 186240 276078 186268 295287
rect 186976 289814 187004 327694
rect 187068 296070 187096 489874
rect 187160 377369 187188 502318
rect 187240 462392 187292 462398
rect 187240 462334 187292 462340
rect 187252 448526 187280 462334
rect 187240 448520 187292 448526
rect 187240 448462 187292 448468
rect 187146 377360 187202 377369
rect 187146 377295 187202 377304
rect 187146 363080 187202 363089
rect 187146 363015 187202 363024
rect 187056 296064 187108 296070
rect 187056 296006 187108 296012
rect 186964 289808 187016 289814
rect 186964 289750 187016 289756
rect 187054 289776 187110 289785
rect 187054 289711 187110 289720
rect 187068 289105 187096 289711
rect 187054 289096 187110 289105
rect 187054 289031 187110 289040
rect 187068 278089 187096 289031
rect 187054 278080 187110 278089
rect 187054 278015 187110 278024
rect 186228 276072 186280 276078
rect 186228 276014 186280 276020
rect 185768 270496 185820 270502
rect 185768 270438 185820 270444
rect 185676 259412 185728 259418
rect 185676 259354 185728 259360
rect 185584 258120 185636 258126
rect 185584 258062 185636 258068
rect 185032 234660 185084 234666
rect 185032 234602 185084 234608
rect 185596 204950 185624 258062
rect 185780 253230 185808 270438
rect 187160 268569 187188 363015
rect 188356 360369 188384 557534
rect 190368 554872 190420 554878
rect 190368 554814 190420 554820
rect 188436 545216 188488 545222
rect 188436 545158 188488 545164
rect 188448 518906 188476 545158
rect 189724 541068 189776 541074
rect 189724 541010 189776 541016
rect 188894 538248 188950 538257
rect 188894 538183 188950 538192
rect 188436 518900 188488 518906
rect 188436 518842 188488 518848
rect 188804 388544 188856 388550
rect 188804 388486 188856 388492
rect 188816 373318 188844 388486
rect 188804 373312 188856 373318
rect 188804 373254 188856 373260
rect 188434 367160 188490 367169
rect 188434 367095 188490 367104
rect 188342 360360 188398 360369
rect 188342 360295 188398 360304
rect 187238 345808 187294 345817
rect 187238 345743 187294 345752
rect 187252 331906 187280 345743
rect 187240 331900 187292 331906
rect 187240 331842 187292 331848
rect 188356 320929 188384 360295
rect 188448 341562 188476 367095
rect 188908 351257 188936 538183
rect 188986 534168 189042 534177
rect 188986 534103 189042 534112
rect 188894 351248 188950 351257
rect 188894 351183 188950 351192
rect 188528 349852 188580 349858
rect 188528 349794 188580 349800
rect 188436 341556 188488 341562
rect 188436 341498 188488 341504
rect 188436 334620 188488 334626
rect 188436 334562 188488 334568
rect 188342 320920 188398 320929
rect 188342 320855 188398 320864
rect 187608 311228 187660 311234
rect 187608 311170 187660 311176
rect 187516 291372 187568 291378
rect 187516 291314 187568 291320
rect 187240 276072 187292 276078
rect 187240 276014 187292 276020
rect 187146 268560 187202 268569
rect 187146 268495 187202 268504
rect 187252 264217 187280 276014
rect 187332 268388 187384 268394
rect 187332 268330 187384 268336
rect 187344 267782 187372 268330
rect 187332 267776 187384 267782
rect 187384 267724 187464 267734
rect 187332 267718 187464 267724
rect 187344 267706 187464 267718
rect 187238 264208 187294 264217
rect 187238 264143 187294 264152
rect 186962 263800 187018 263809
rect 186962 263735 187018 263744
rect 185768 253224 185820 253230
rect 185768 253166 185820 253172
rect 186226 245848 186282 245857
rect 186226 245783 186282 245792
rect 185676 230444 185728 230450
rect 185676 230386 185728 230392
rect 185584 204944 185636 204950
rect 185584 204886 185636 204892
rect 185688 192506 185716 230386
rect 185676 192500 185728 192506
rect 185676 192442 185728 192448
rect 186240 182889 186268 245783
rect 186318 241360 186374 241369
rect 186318 241295 186374 241304
rect 186332 240174 186360 241295
rect 186320 240168 186372 240174
rect 186320 240110 186372 240116
rect 186226 182880 186282 182889
rect 186226 182815 186282 182824
rect 184846 151056 184902 151065
rect 184846 150991 184902 151000
rect 185676 144968 185728 144974
rect 185676 144910 185728 144916
rect 184296 141432 184348 141438
rect 184296 141374 184348 141380
rect 184308 26897 184336 141374
rect 185584 134564 185636 134570
rect 185584 134506 185636 134512
rect 184386 118824 184442 118833
rect 184386 118759 184442 118768
rect 184400 81394 184428 118759
rect 185596 93401 185624 134506
rect 185688 104242 185716 144910
rect 185768 106412 185820 106418
rect 185768 106354 185820 106360
rect 185676 104236 185728 104242
rect 185676 104178 185728 104184
rect 185582 93392 185638 93401
rect 185582 93327 185638 93336
rect 185584 90432 185636 90438
rect 185584 90374 185636 90380
rect 184388 81388 184440 81394
rect 184388 81330 184440 81336
rect 185596 26926 185624 90374
rect 185780 86873 185808 106354
rect 185766 86864 185822 86873
rect 185766 86799 185822 86808
rect 186976 50386 187004 263735
rect 187148 248464 187200 248470
rect 187148 248406 187200 248412
rect 187056 240848 187108 240854
rect 187056 240790 187108 240796
rect 187068 210458 187096 240790
rect 187160 235657 187188 248406
rect 187146 235648 187202 235657
rect 187146 235583 187202 235592
rect 187436 211993 187464 267706
rect 187528 242214 187556 291314
rect 187620 267714 187648 311170
rect 188342 307184 188398 307193
rect 188342 307119 188398 307128
rect 188356 282849 188384 307119
rect 188448 304366 188476 334562
rect 188540 325650 188568 349794
rect 188528 325644 188580 325650
rect 188528 325586 188580 325592
rect 188436 304360 188488 304366
rect 188436 304302 188488 304308
rect 188436 289808 188488 289814
rect 188436 289750 188488 289756
rect 188342 282840 188398 282849
rect 188342 282775 188398 282784
rect 187608 267708 187660 267714
rect 187608 267650 187660 267656
rect 188342 265160 188398 265169
rect 188342 265095 188398 265104
rect 187516 242208 187568 242214
rect 187516 242150 187568 242156
rect 188356 234569 188384 265095
rect 188448 261526 188476 289750
rect 188526 285152 188582 285161
rect 188526 285087 188582 285096
rect 188540 264926 188568 285087
rect 188528 264920 188580 264926
rect 188528 264862 188580 264868
rect 188436 261520 188488 261526
rect 188436 261462 188488 261468
rect 188436 259480 188488 259486
rect 188436 259422 188488 259428
rect 188342 234560 188398 234569
rect 188342 234495 188398 234504
rect 187422 211984 187478 211993
rect 187422 211919 187478 211928
rect 187056 210452 187108 210458
rect 187056 210394 187108 210400
rect 188356 188465 188384 234495
rect 188448 233238 188476 259422
rect 188436 233232 188488 233238
rect 188436 233174 188488 233180
rect 187054 188456 187110 188465
rect 187054 188391 187110 188400
rect 188342 188456 188398 188465
rect 188448 188426 188476 233174
rect 189000 212401 189028 534103
rect 189736 508570 189764 541010
rect 189724 508564 189776 508570
rect 189724 508506 189776 508512
rect 190276 448588 190328 448594
rect 190276 448530 190328 448536
rect 189816 404388 189868 404394
rect 189816 404330 189868 404336
rect 189724 374060 189776 374066
rect 189724 374002 189776 374008
rect 189736 345710 189764 374002
rect 189724 345704 189776 345710
rect 189724 345646 189776 345652
rect 189722 333024 189778 333033
rect 189722 332959 189778 332968
rect 189736 258194 189764 332959
rect 189828 331945 189856 404330
rect 190288 377466 190316 448530
rect 190276 377460 190328 377466
rect 190276 377402 190328 377408
rect 189908 368484 189960 368490
rect 189908 368426 189960 368432
rect 189920 363730 189948 368426
rect 190380 367810 190408 554814
rect 191116 534070 191144 563042
rect 195888 558952 195940 558958
rect 195888 558894 195940 558900
rect 192484 552084 192536 552090
rect 192484 552026 192536 552032
rect 191194 550896 191250 550905
rect 191194 550831 191250 550840
rect 191104 534064 191156 534070
rect 191104 534006 191156 534012
rect 191208 528554 191236 550831
rect 191746 534984 191802 534993
rect 191746 534919 191802 534928
rect 191116 528526 191236 528554
rect 191116 525094 191144 528526
rect 191104 525088 191156 525094
rect 191104 525030 191156 525036
rect 190460 378208 190512 378214
rect 190460 378150 190512 378156
rect 190368 367804 190420 367810
rect 190368 367746 190420 367752
rect 189908 363724 189960 363730
rect 189908 363666 189960 363672
rect 190472 343670 190500 378150
rect 191116 367849 191144 525030
rect 191760 460902 191788 534919
rect 191748 460896 191800 460902
rect 191748 460838 191800 460844
rect 191760 460222 191788 460838
rect 191748 460216 191800 460222
rect 191748 460158 191800 460164
rect 191288 455456 191340 455462
rect 191288 455398 191340 455404
rect 191196 386436 191248 386442
rect 191196 386378 191248 386384
rect 191102 367840 191158 367849
rect 191102 367775 191158 367784
rect 190460 343664 190512 343670
rect 190460 343606 190512 343612
rect 189906 340912 189962 340921
rect 189906 340847 189962 340856
rect 189814 331936 189870 331945
rect 189814 331871 189870 331880
rect 189920 295390 189948 340847
rect 191104 331968 191156 331974
rect 191104 331910 191156 331916
rect 190276 307080 190328 307086
rect 190276 307022 190328 307028
rect 189908 295384 189960 295390
rect 189908 295326 189960 295332
rect 189816 265736 189868 265742
rect 189816 265678 189868 265684
rect 189724 258188 189776 258194
rect 189724 258130 189776 258136
rect 189724 256828 189776 256834
rect 189724 256770 189776 256776
rect 189736 254590 189764 256770
rect 189724 254584 189776 254590
rect 189724 254526 189776 254532
rect 189080 244928 189132 244934
rect 189736 244905 189764 254526
rect 189828 249422 189856 265678
rect 189816 249416 189868 249422
rect 189816 249358 189868 249364
rect 189080 244870 189132 244876
rect 189722 244896 189778 244905
rect 189092 242321 189120 244870
rect 189722 244831 189778 244840
rect 190184 243024 190236 243030
rect 190184 242966 190236 242972
rect 189078 242312 189134 242321
rect 189078 242247 189134 242256
rect 190196 220561 190224 242966
rect 190288 238377 190316 307022
rect 191116 297537 191144 331910
rect 191102 297528 191158 297537
rect 191102 297463 191158 297472
rect 190368 295384 190420 295390
rect 190368 295326 190420 295332
rect 190380 264926 190408 295326
rect 191104 285728 191156 285734
rect 191104 285670 191156 285676
rect 190368 264920 190420 264926
rect 190368 264862 190420 264868
rect 191116 258126 191144 285670
rect 191104 258120 191156 258126
rect 191104 258062 191156 258068
rect 191104 249824 191156 249830
rect 191104 249766 191156 249772
rect 190368 244928 190420 244934
rect 190368 244870 190420 244876
rect 190274 238368 190330 238377
rect 190274 238303 190330 238312
rect 190182 220552 190238 220561
rect 190182 220487 190238 220496
rect 190196 219473 190224 220487
rect 190182 219464 190238 219473
rect 190182 219399 190238 219408
rect 188986 212392 189042 212401
rect 188986 212327 189042 212336
rect 189724 196648 189776 196654
rect 189724 196590 189776 196596
rect 188342 188391 188398 188400
rect 188436 188420 188488 188426
rect 187068 98705 187096 188391
rect 188436 188362 188488 188368
rect 187148 186380 187200 186386
rect 187148 186322 187200 186328
rect 187160 162790 187188 186322
rect 187148 162784 187200 162790
rect 187148 162726 187200 162732
rect 187148 127016 187200 127022
rect 187148 126958 187200 126964
rect 187054 98696 187110 98705
rect 187054 98631 187110 98640
rect 187160 91866 187188 126958
rect 188344 118040 188396 118046
rect 188344 117982 188396 117988
rect 187148 91860 187200 91866
rect 187148 91802 187200 91808
rect 186964 50380 187016 50386
rect 186964 50322 187016 50328
rect 186964 35284 187016 35290
rect 186964 35226 187016 35232
rect 185584 26920 185636 26926
rect 184294 26888 184350 26897
rect 185584 26862 185636 26868
rect 184294 26823 184350 26832
rect 184202 7576 184258 7585
rect 184202 7511 184258 7520
rect 182822 6896 182878 6905
rect 182822 6831 182878 6840
rect 186976 4826 187004 35226
rect 188356 28286 188384 117982
rect 188436 116068 188488 116074
rect 188436 116010 188488 116016
rect 188448 85542 188476 116010
rect 188436 85536 188488 85542
rect 188436 85478 188488 85484
rect 188344 28280 188396 28286
rect 189736 28257 189764 196590
rect 190380 172446 190408 244870
rect 190458 231296 190514 231305
rect 190458 231231 190514 231240
rect 190472 227730 190500 231231
rect 190460 227724 190512 227730
rect 190460 227666 190512 227672
rect 191116 213926 191144 249766
rect 191208 242962 191236 386378
rect 191300 378214 191328 455398
rect 191380 385688 191432 385694
rect 191380 385630 191432 385636
rect 191288 378208 191340 378214
rect 191288 378150 191340 378156
rect 191392 375358 191420 385630
rect 191380 375352 191432 375358
rect 191380 375294 191432 375300
rect 191288 369232 191340 369238
rect 191288 369174 191340 369180
rect 191300 266966 191328 369174
rect 192496 355026 192524 552026
rect 193954 550760 194010 550769
rect 193954 550695 194010 550704
rect 193864 548004 193916 548010
rect 193864 547946 193916 547952
rect 192574 537160 192630 537169
rect 192574 537095 192630 537104
rect 192588 443698 192616 537095
rect 192666 451888 192722 451897
rect 192666 451823 192722 451832
rect 192576 443692 192628 443698
rect 192576 443634 192628 443640
rect 192680 441454 192708 451823
rect 192668 441448 192720 441454
rect 192668 441390 192720 441396
rect 192576 427848 192628 427854
rect 192576 427790 192628 427796
rect 192484 355020 192536 355026
rect 192484 354962 192536 354968
rect 192496 354754 192524 354962
rect 192484 354748 192536 354754
rect 192484 354690 192536 354696
rect 192484 313336 192536 313342
rect 192484 313278 192536 313284
rect 191840 279472 191892 279478
rect 191840 279414 191892 279420
rect 191852 273494 191880 279414
rect 191840 273488 191892 273494
rect 191840 273430 191892 273436
rect 191380 272536 191432 272542
rect 191380 272478 191432 272484
rect 191288 266960 191340 266966
rect 191288 266902 191340 266908
rect 191288 260160 191340 260166
rect 191288 260102 191340 260108
rect 191196 242956 191248 242962
rect 191196 242898 191248 242904
rect 191208 235249 191236 242898
rect 191194 235240 191250 235249
rect 191194 235175 191250 235184
rect 191196 233912 191248 233918
rect 191196 233854 191248 233860
rect 191208 223514 191236 233854
rect 191300 233238 191328 260102
rect 191392 251258 191420 272478
rect 191840 258528 191892 258534
rect 191840 258470 191892 258476
rect 191852 258194 191880 258470
rect 191840 258188 191892 258194
rect 191840 258130 191892 258136
rect 191380 251252 191432 251258
rect 191380 251194 191432 251200
rect 191748 250504 191800 250510
rect 191748 250446 191800 250452
rect 191760 249558 191788 250446
rect 191748 249552 191800 249558
rect 191748 249494 191800 249500
rect 191654 246528 191710 246537
rect 191654 246463 191710 246472
rect 191668 245721 191696 246463
rect 191654 245712 191710 245721
rect 191852 245698 191880 258130
rect 191654 245647 191710 245656
rect 191760 245670 191880 245698
rect 192206 245712 192262 245721
rect 191288 233232 191340 233238
rect 191288 233174 191340 233180
rect 191656 232552 191708 232558
rect 191656 232494 191708 232500
rect 191668 231810 191696 232494
rect 191656 231804 191708 231810
rect 191656 231746 191708 231752
rect 191196 223508 191248 223514
rect 191196 223450 191248 223456
rect 191104 213920 191156 213926
rect 191104 213862 191156 213868
rect 191116 185706 191144 213862
rect 191760 186998 191788 245670
rect 192206 245647 192262 245656
rect 192220 240281 192248 245647
rect 192206 240272 192262 240281
rect 192206 240207 192262 240216
rect 191840 239420 191892 239426
rect 191840 239362 191892 239368
rect 191852 237726 191880 239362
rect 191840 237720 191892 237726
rect 191840 237662 191892 237668
rect 192496 233170 192524 313278
rect 192588 291378 192616 427790
rect 192668 399492 192720 399498
rect 192668 399434 192720 399440
rect 192680 376825 192708 399434
rect 193128 383716 193180 383722
rect 193128 383658 193180 383664
rect 193140 382401 193168 383658
rect 193126 382392 193182 382401
rect 193126 382327 193182 382336
rect 192666 376816 192722 376825
rect 192666 376751 192722 376760
rect 192760 355020 192812 355026
rect 192760 354962 192812 354968
rect 192668 334008 192720 334014
rect 192668 333950 192720 333956
rect 192576 291372 192628 291378
rect 192576 291314 192628 291320
rect 192680 278730 192708 333950
rect 192772 304366 192800 354962
rect 193876 349178 193904 547946
rect 193968 507142 193996 550695
rect 194508 543856 194560 543862
rect 194508 543798 194560 543804
rect 193956 507136 194008 507142
rect 193956 507078 194008 507084
rect 193956 453552 194008 453558
rect 193956 453494 194008 453500
rect 193968 400926 193996 453494
rect 193956 400920 194008 400926
rect 193956 400862 194008 400868
rect 193864 349172 193916 349178
rect 193864 349114 193916 349120
rect 192760 304360 192812 304366
rect 192760 304302 192812 304308
rect 193404 302932 193456 302938
rect 193404 302874 193456 302880
rect 193416 297430 193444 302874
rect 193876 301510 193904 349114
rect 193968 338745 193996 400862
rect 194048 398880 194100 398886
rect 194048 398822 194100 398828
rect 194060 388550 194088 398822
rect 194048 388544 194100 388550
rect 194048 388486 194100 388492
rect 194416 380180 194468 380186
rect 194416 380122 194468 380128
rect 193954 338736 194010 338745
rect 193954 338671 194010 338680
rect 194046 336832 194102 336841
rect 194046 336767 194102 336776
rect 194060 318170 194088 336767
rect 193956 318164 194008 318170
rect 193956 318106 194008 318112
rect 194048 318164 194100 318170
rect 194048 318106 194100 318112
rect 193864 301504 193916 301510
rect 193864 301446 193916 301452
rect 193968 297566 193996 318106
rect 194324 298172 194376 298178
rect 194324 298114 194376 298120
rect 193956 297560 194008 297566
rect 193956 297502 194008 297508
rect 193404 297424 193456 297430
rect 193404 297366 193456 297372
rect 193126 293176 193182 293185
rect 193126 293111 193182 293120
rect 192668 278724 192720 278730
rect 192668 278666 192720 278672
rect 193036 273488 193088 273494
rect 193036 273430 193088 273436
rect 192944 236768 192996 236774
rect 192944 236710 192996 236716
rect 192956 233889 192984 236710
rect 192666 233880 192722 233889
rect 192666 233815 192722 233824
rect 192942 233880 192998 233889
rect 192942 233815 192998 233824
rect 192484 233164 192536 233170
rect 192484 233106 192536 233112
rect 192482 219464 192538 219473
rect 192482 219399 192538 219408
rect 192496 211138 192524 219399
rect 192574 218648 192630 218657
rect 192574 218583 192630 218592
rect 192484 211132 192536 211138
rect 192484 211074 192536 211080
rect 191838 202192 191894 202201
rect 191838 202127 191894 202136
rect 191852 197305 191880 202127
rect 191838 197296 191894 197305
rect 191838 197231 191894 197240
rect 191748 186992 191800 186998
rect 191748 186934 191800 186940
rect 191104 185700 191156 185706
rect 191104 185642 191156 185648
rect 191104 184952 191156 184958
rect 191104 184894 191156 184900
rect 190368 172440 190420 172446
rect 190368 172382 190420 172388
rect 191116 150346 191144 184894
rect 191104 150340 191156 150346
rect 191104 150282 191156 150288
rect 191104 142248 191156 142254
rect 191104 142190 191156 142196
rect 191116 117978 191144 142190
rect 191288 140820 191340 140826
rect 191288 140762 191340 140768
rect 191196 120216 191248 120222
rect 191196 120158 191248 120164
rect 191104 117972 191156 117978
rect 191104 117914 191156 117920
rect 189816 98048 189868 98054
rect 189816 97990 189868 97996
rect 189828 82822 189856 97990
rect 191102 94480 191158 94489
rect 191102 94415 191158 94424
rect 189816 82816 189868 82822
rect 189816 82758 189868 82764
rect 188344 28222 188396 28228
rect 189722 28248 189778 28257
rect 189722 28183 189778 28192
rect 189724 20052 189776 20058
rect 189724 19994 189776 20000
rect 186964 4820 187016 4826
rect 186964 4762 187016 4768
rect 189736 3369 189764 19994
rect 191116 6254 191144 94415
rect 191208 52426 191236 120158
rect 191300 90953 191328 140762
rect 192484 140072 192536 140078
rect 192484 140014 192536 140020
rect 191286 90944 191342 90953
rect 191286 90879 191342 90888
rect 191196 52420 191248 52426
rect 191196 52362 191248 52368
rect 192496 48278 192524 140014
rect 192588 130490 192616 218583
rect 192680 218074 192708 233815
rect 192942 220280 192998 220289
rect 192942 220215 192998 220224
rect 192956 220114 192984 220215
rect 192944 220108 192996 220114
rect 192944 220050 192996 220056
rect 192668 218068 192720 218074
rect 192668 218010 192720 218016
rect 193048 217734 193076 273430
rect 193140 262274 193168 293111
rect 193864 292664 193916 292670
rect 193864 292606 193916 292612
rect 193220 266960 193272 266966
rect 193220 266902 193272 266908
rect 193128 262268 193180 262274
rect 193128 262210 193180 262216
rect 193232 255377 193260 266902
rect 193218 255368 193274 255377
rect 193218 255303 193274 255312
rect 193128 251252 193180 251258
rect 193128 251194 193180 251200
rect 193140 248742 193168 251194
rect 193128 248736 193180 248742
rect 193128 248678 193180 248684
rect 193036 217728 193088 217734
rect 193036 217670 193088 217676
rect 193140 178673 193168 248678
rect 193876 241505 193904 292606
rect 194336 267170 194364 298114
rect 194428 269074 194456 380122
rect 194520 377505 194548 543798
rect 195242 542736 195298 542745
rect 195242 542671 195298 542680
rect 195152 539708 195204 539714
rect 195152 539650 195204 539656
rect 195164 538966 195192 539650
rect 195152 538960 195204 538966
rect 195152 538902 195204 538908
rect 195256 538898 195284 542671
rect 195336 542496 195388 542502
rect 195336 542438 195388 542444
rect 195244 538892 195296 538898
rect 195244 538834 195296 538840
rect 195244 538348 195296 538354
rect 195244 538290 195296 538296
rect 195256 380225 195284 538290
rect 195348 523734 195376 542438
rect 195336 523728 195388 523734
rect 195336 523670 195388 523676
rect 195520 380928 195572 380934
rect 195520 380870 195572 380876
rect 195242 380216 195298 380225
rect 195242 380151 195298 380160
rect 195336 379636 195388 379642
rect 195336 379578 195388 379584
rect 195242 378720 195298 378729
rect 195242 378655 195298 378664
rect 194506 377496 194562 377505
rect 194506 377431 194562 377440
rect 195256 369238 195284 378655
rect 195244 369232 195296 369238
rect 195244 369174 195296 369180
rect 194600 367124 194652 367130
rect 194600 367066 194652 367072
rect 194612 311234 194640 367066
rect 195242 362264 195298 362273
rect 195242 362199 195298 362208
rect 195256 329089 195284 362199
rect 195348 359582 195376 379578
rect 195428 363724 195480 363730
rect 195428 363666 195480 363672
rect 195336 359576 195388 359582
rect 195336 359518 195388 359524
rect 195334 338192 195390 338201
rect 195334 338127 195390 338136
rect 195242 329080 195298 329089
rect 195242 329015 195298 329024
rect 195244 326392 195296 326398
rect 195244 326334 195296 326340
rect 194600 311228 194652 311234
rect 194600 311170 194652 311176
rect 194600 310548 194652 310554
rect 194600 310490 194652 310496
rect 194506 287464 194562 287473
rect 194506 287399 194562 287408
rect 194416 269068 194468 269074
rect 194416 269010 194468 269016
rect 194324 267164 194376 267170
rect 194324 267106 194376 267112
rect 194336 265674 194364 267106
rect 194324 265668 194376 265674
rect 194324 265610 194376 265616
rect 194414 255368 194470 255377
rect 194414 255303 194470 255312
rect 194428 255270 194456 255303
rect 194416 255264 194468 255270
rect 194416 255206 194468 255212
rect 194324 251932 194376 251938
rect 194324 251874 194376 251880
rect 194336 251666 194364 251874
rect 194324 251660 194376 251666
rect 194324 251602 194376 251608
rect 194232 245676 194284 245682
rect 194232 245618 194284 245624
rect 193862 241496 193918 241505
rect 193862 241431 193918 241440
rect 194244 230450 194272 245618
rect 194232 230444 194284 230450
rect 194232 230386 194284 230392
rect 194232 229764 194284 229770
rect 194232 229706 194284 229712
rect 194244 229022 194272 229706
rect 194232 229016 194284 229022
rect 194232 228958 194284 228964
rect 194336 221474 194364 251602
rect 194416 237720 194468 237726
rect 194416 237662 194468 237668
rect 194324 221468 194376 221474
rect 194324 221410 194376 221416
rect 193862 215928 193918 215937
rect 193862 215863 193918 215872
rect 193876 208350 193904 215863
rect 193864 208344 193916 208350
rect 193864 208286 193916 208292
rect 194428 199510 194456 237662
rect 194520 200122 194548 287399
rect 194612 245682 194640 310490
rect 195152 291304 195204 291310
rect 195152 291246 195204 291252
rect 195164 290494 195192 291246
rect 195152 290488 195204 290494
rect 195152 290430 195204 290436
rect 195150 288552 195206 288561
rect 195150 288487 195206 288496
rect 195164 287706 195192 288487
rect 195152 287700 195204 287706
rect 195152 287642 195204 287648
rect 195150 285696 195206 285705
rect 195150 285631 195206 285640
rect 195164 282878 195192 285631
rect 195152 282872 195204 282878
rect 195152 282814 195204 282820
rect 194692 269068 194744 269074
rect 194692 269010 194744 269016
rect 194704 268054 194732 269010
rect 194692 268048 194744 268054
rect 194692 267990 194744 267996
rect 194704 262886 194732 267990
rect 195150 265568 195206 265577
rect 195150 265503 195206 265512
rect 195164 265033 195192 265503
rect 195150 265024 195206 265033
rect 195150 264959 195206 264968
rect 194692 262880 194744 262886
rect 194692 262822 194744 262828
rect 194784 262268 194836 262274
rect 194784 262210 194836 262216
rect 194796 251841 194824 262210
rect 194782 251832 194838 251841
rect 194782 251767 194838 251776
rect 194600 245676 194652 245682
rect 194600 245618 194652 245624
rect 195256 240106 195284 326334
rect 195348 301753 195376 338127
rect 195440 331294 195468 363666
rect 195532 362302 195560 380870
rect 195900 376145 195928 558894
rect 197176 553512 197228 553518
rect 197176 553454 197228 553460
rect 196714 541104 196770 541113
rect 196714 541039 196770 541048
rect 196624 534812 196676 534818
rect 196624 534754 196676 534760
rect 195886 376136 195942 376145
rect 195886 376071 195942 376080
rect 195888 375420 195940 375426
rect 195888 375362 195940 375368
rect 195900 368393 195928 375362
rect 195886 368384 195942 368393
rect 195886 368319 195942 368328
rect 195520 362296 195572 362302
rect 195520 362238 195572 362244
rect 195518 358864 195574 358873
rect 195518 358799 195574 358808
rect 195532 342922 195560 358799
rect 196636 351966 196664 534754
rect 196728 519586 196756 541039
rect 196716 519580 196768 519586
rect 196716 519522 196768 519528
rect 197082 470928 197138 470937
rect 197082 470863 197138 470872
rect 196714 384976 196770 384985
rect 196714 384911 196770 384920
rect 196728 383722 196756 384911
rect 196716 383716 196768 383722
rect 196716 383658 196768 383664
rect 196728 364313 196756 383658
rect 197096 375698 197124 470863
rect 197084 375692 197136 375698
rect 197084 375634 197136 375640
rect 197188 373386 197216 553454
rect 197280 444258 197308 702646
rect 213920 565888 213972 565894
rect 213920 565830 213972 565836
rect 197360 562352 197412 562358
rect 197360 562294 197412 562300
rect 197372 561814 197400 562294
rect 197360 561808 197412 561814
rect 197360 561750 197412 561756
rect 197372 453558 197400 561750
rect 205638 559056 205694 559065
rect 205638 558991 205694 559000
rect 209780 559020 209832 559026
rect 198648 558204 198700 558210
rect 198648 558146 198700 558152
rect 198554 554024 198610 554033
rect 198554 553959 198610 553968
rect 197544 536920 197596 536926
rect 197544 536862 197596 536868
rect 197452 532704 197504 532710
rect 197452 532646 197504 532652
rect 197464 532273 197492 532646
rect 197450 532264 197506 532273
rect 197450 532199 197506 532208
rect 197556 530670 197584 536862
rect 197544 530664 197596 530670
rect 197544 530606 197596 530612
rect 197452 529848 197504 529854
rect 197450 529816 197452 529825
rect 198568 529825 198596 553959
rect 197504 529816 197506 529825
rect 197450 529751 197506 529760
rect 198554 529816 198610 529825
rect 198554 529751 198610 529760
rect 197452 528556 197504 528562
rect 197452 528498 197504 528504
rect 197464 527377 197492 528498
rect 197450 527368 197506 527377
rect 197450 527303 197506 527312
rect 197542 524784 197598 524793
rect 197542 524719 197598 524728
rect 197450 522336 197506 522345
rect 197450 522271 197506 522280
rect 197464 521694 197492 522271
rect 197452 521688 197504 521694
rect 197452 521630 197504 521636
rect 197556 521014 197584 524719
rect 197544 521008 197596 521014
rect 197544 520950 197596 520956
rect 197450 517440 197506 517449
rect 197450 517375 197506 517384
rect 197464 516186 197492 517375
rect 197452 516180 197504 516186
rect 197452 516122 197504 516128
rect 197452 510604 197504 510610
rect 197452 510546 197504 510552
rect 197464 510241 197492 510546
rect 197450 510232 197506 510241
rect 197450 510167 197506 510176
rect 197450 507648 197506 507657
rect 197450 507583 197506 507592
rect 197464 502994 197492 507583
rect 197452 502988 197504 502994
rect 197452 502930 197504 502936
rect 197450 502752 197506 502761
rect 197450 502687 197506 502696
rect 197464 502382 197492 502687
rect 197452 502376 197504 502382
rect 197452 502318 197504 502324
rect 197452 500948 197504 500954
rect 197452 500890 197504 500896
rect 197464 500449 197492 500890
rect 198660 500449 198688 558146
rect 198832 551336 198884 551342
rect 198832 551278 198884 551284
rect 198738 538384 198794 538393
rect 198738 538319 198794 538328
rect 198752 534750 198780 538319
rect 198740 534744 198792 534750
rect 198740 534686 198792 534692
rect 197450 500440 197506 500449
rect 197450 500375 197506 500384
rect 198646 500440 198702 500449
rect 198646 500375 198702 500384
rect 197450 495544 197506 495553
rect 197450 495479 197452 495488
rect 197504 495479 197506 495488
rect 197452 495450 197504 495456
rect 197450 492960 197506 492969
rect 197450 492895 197506 492904
rect 197464 492726 197492 492895
rect 197452 492720 197504 492726
rect 197452 492662 197504 492668
rect 197450 490512 197506 490521
rect 197450 490447 197506 490456
rect 197464 489938 197492 490447
rect 197452 489932 197504 489938
rect 197452 489874 197504 489880
rect 197450 488064 197506 488073
rect 197450 487999 197506 488008
rect 197464 487218 197492 487999
rect 197452 487212 197504 487218
rect 197452 487154 197504 487160
rect 197450 485616 197506 485625
rect 197450 485551 197506 485560
rect 197464 483682 197492 485551
rect 197452 483676 197504 483682
rect 197452 483618 197504 483624
rect 198002 483168 198058 483177
rect 198002 483103 198058 483112
rect 197450 480720 197506 480729
rect 197450 480655 197506 480664
rect 197464 480282 197492 480655
rect 197452 480276 197504 480282
rect 197452 480218 197504 480224
rect 197450 478272 197506 478281
rect 197450 478207 197506 478216
rect 197464 477562 197492 478207
rect 197452 477556 197504 477562
rect 197452 477498 197504 477504
rect 197450 475824 197506 475833
rect 197450 475759 197506 475768
rect 197464 474774 197492 475759
rect 197452 474768 197504 474774
rect 197452 474710 197504 474716
rect 197452 473408 197504 473414
rect 197450 473376 197452 473385
rect 197504 473376 197506 473385
rect 197450 473311 197506 473320
rect 197450 468480 197506 468489
rect 197450 468415 197506 468424
rect 197464 467906 197492 468415
rect 197452 467900 197504 467906
rect 197452 467842 197504 467848
rect 197450 466032 197506 466041
rect 197450 465967 197506 465976
rect 197464 465730 197492 465967
rect 197452 465724 197504 465730
rect 197452 465666 197504 465672
rect 197450 463312 197506 463321
rect 197450 463247 197506 463256
rect 197464 462398 197492 463247
rect 197452 462392 197504 462398
rect 197452 462334 197504 462340
rect 197452 460896 197504 460902
rect 197450 460864 197452 460873
rect 197504 460864 197506 460873
rect 197450 460799 197506 460808
rect 197450 455968 197506 455977
rect 197450 455903 197506 455912
rect 197464 455462 197492 455903
rect 197452 455456 197504 455462
rect 197452 455398 197504 455404
rect 197360 453552 197412 453558
rect 197360 453494 197412 453500
rect 197358 448624 197414 448633
rect 197358 448559 197360 448568
rect 197412 448559 197414 448568
rect 197360 448530 197412 448536
rect 197358 446176 197414 446185
rect 197358 446111 197414 446120
rect 197372 445806 197400 446111
rect 197360 445800 197412 445806
rect 197360 445742 197412 445748
rect 197280 444230 197400 444258
rect 197372 443766 197400 444230
rect 197360 443760 197412 443766
rect 197358 443728 197360 443737
rect 197412 443728 197414 443737
rect 197358 443663 197414 443672
rect 197728 441448 197780 441454
rect 197726 441416 197728 441425
rect 197780 441416 197782 441425
rect 197726 441351 197782 441360
rect 197358 436384 197414 436393
rect 197358 436319 197414 436328
rect 197372 436150 197400 436319
rect 197360 436144 197412 436150
rect 197360 436086 197412 436092
rect 197358 433936 197414 433945
rect 197358 433871 197414 433880
rect 197372 433362 197400 433871
rect 197360 433356 197412 433362
rect 197360 433298 197412 433304
rect 197358 429040 197414 429049
rect 197358 428975 197414 428984
rect 197372 427854 197400 428975
rect 197360 427848 197412 427854
rect 197360 427790 197412 427796
rect 197358 426592 197414 426601
rect 197358 426527 197414 426536
rect 197372 426494 197400 426527
rect 197360 426488 197412 426494
rect 197360 426430 197412 426436
rect 197358 424144 197414 424153
rect 197358 424079 197414 424088
rect 197372 423706 197400 424079
rect 197360 423700 197412 423706
rect 197360 423642 197412 423648
rect 197358 419248 197414 419257
rect 197358 419183 197414 419192
rect 197372 418198 197400 419183
rect 197360 418192 197412 418198
rect 197360 418134 197412 418140
rect 197358 414352 197414 414361
rect 197358 414287 197414 414296
rect 197372 414050 197400 414287
rect 197360 414044 197412 414050
rect 197360 413986 197412 413992
rect 197358 411904 197414 411913
rect 197358 411839 197414 411848
rect 197372 411330 197400 411839
rect 197360 411324 197412 411330
rect 197360 411266 197412 411272
rect 197360 409828 197412 409834
rect 197360 409770 197412 409776
rect 197372 409601 197400 409770
rect 197358 409592 197414 409601
rect 197358 409527 197414 409536
rect 197358 407008 197414 407017
rect 197358 406943 197414 406952
rect 197372 405754 197400 406943
rect 197360 405748 197412 405754
rect 197360 405690 197412 405696
rect 197358 404560 197414 404569
rect 197358 404495 197414 404504
rect 197372 404394 197400 404495
rect 197360 404388 197412 404394
rect 197360 404330 197412 404336
rect 197358 399664 197414 399673
rect 197358 399599 197414 399608
rect 197372 398886 197400 399599
rect 197360 398880 197412 398886
rect 197360 398822 197412 398828
rect 197358 394768 197414 394777
rect 197358 394703 197360 394712
rect 197412 394703 197414 394712
rect 197360 394674 197412 394680
rect 197360 390516 197412 390522
rect 197360 390458 197412 390464
rect 197372 390017 197400 390458
rect 197358 390008 197414 390017
rect 197358 389943 197414 389952
rect 197358 387424 197414 387433
rect 197358 387359 197414 387368
rect 197372 386442 197400 387359
rect 197360 386436 197412 386442
rect 197360 386378 197412 386384
rect 197358 385112 197414 385121
rect 197358 385047 197360 385056
rect 197412 385047 197414 385056
rect 197360 385018 197412 385024
rect 197358 380216 197414 380225
rect 197358 380151 197360 380160
rect 197412 380151 197414 380160
rect 197360 380122 197412 380128
rect 197176 373380 197228 373386
rect 197176 373322 197228 373328
rect 196808 372632 196860 372638
rect 196808 372574 196860 372580
rect 196714 364304 196770 364313
rect 196714 364239 196770 364248
rect 196820 355434 196848 372574
rect 196808 355428 196860 355434
rect 196808 355370 196860 355376
rect 196624 351960 196676 351966
rect 196624 351902 196676 351908
rect 195520 342916 195572 342922
rect 195520 342858 195572 342864
rect 195428 331288 195480 331294
rect 195428 331230 195480 331236
rect 196636 319433 196664 351902
rect 197268 349852 197320 349858
rect 197268 349794 197320 349800
rect 196714 347032 196770 347041
rect 196714 346967 196770 346976
rect 196622 319424 196678 319433
rect 196622 319359 196678 319368
rect 195980 314696 196032 314702
rect 195980 314638 196032 314644
rect 195992 306374 196020 314638
rect 196728 314129 196756 346967
rect 196714 314120 196770 314129
rect 196714 314055 196770 314064
rect 197176 311160 197228 311166
rect 197176 311102 197228 311108
rect 197084 307148 197136 307154
rect 197084 307090 197136 307096
rect 195900 306346 196020 306374
rect 195334 301744 195390 301753
rect 195334 301679 195390 301688
rect 195336 294024 195388 294030
rect 195336 293966 195388 293972
rect 195348 286346 195376 293966
rect 195900 292618 195928 306346
rect 195900 292590 196020 292618
rect 195992 287054 196020 292590
rect 196622 287328 196678 287337
rect 196622 287263 196678 287272
rect 195900 287026 196020 287054
rect 195336 286340 195388 286346
rect 195336 286282 195388 286288
rect 195900 278662 195928 287026
rect 195888 278656 195940 278662
rect 195888 278598 195940 278604
rect 196636 265742 196664 287263
rect 196624 265736 196676 265742
rect 196624 265678 196676 265684
rect 196808 261520 196860 261526
rect 196808 261462 196860 261468
rect 195888 252612 195940 252618
rect 195888 252554 195940 252560
rect 195336 247104 195388 247110
rect 195336 247046 195388 247052
rect 195244 240100 195296 240106
rect 195244 240042 195296 240048
rect 195242 231976 195298 231985
rect 195242 231911 195298 231920
rect 195256 231577 195284 231911
rect 195242 231568 195298 231577
rect 195242 231503 195298 231512
rect 195244 224256 195296 224262
rect 195244 224198 195296 224204
rect 195256 222154 195284 224198
rect 195244 222148 195296 222154
rect 195244 222090 195296 222096
rect 195244 221536 195296 221542
rect 195244 221478 195296 221484
rect 195256 219201 195284 221478
rect 195242 219192 195298 219201
rect 195242 219127 195298 219136
rect 195244 218068 195296 218074
rect 195244 218010 195296 218016
rect 195256 202201 195284 218010
rect 195348 216578 195376 247046
rect 195794 241496 195850 241505
rect 195794 241431 195850 241440
rect 195808 240854 195836 241431
rect 195796 240848 195848 240854
rect 195796 240790 195848 240796
rect 195808 224913 195836 240790
rect 195794 224904 195850 224913
rect 195794 224839 195850 224848
rect 195704 223508 195756 223514
rect 195704 223450 195756 223456
rect 195428 222216 195480 222222
rect 195428 222158 195480 222164
rect 195440 221921 195468 222158
rect 195426 221912 195482 221921
rect 195426 221847 195482 221856
rect 195716 220726 195744 223450
rect 195704 220720 195756 220726
rect 195704 220662 195756 220668
rect 195426 220144 195482 220153
rect 195426 220079 195482 220088
rect 195336 216572 195388 216578
rect 195336 216514 195388 216520
rect 195242 202192 195298 202201
rect 195242 202127 195298 202136
rect 195348 200870 195376 216514
rect 195336 200864 195388 200870
rect 195336 200806 195388 200812
rect 194508 200116 194560 200122
rect 194508 200058 194560 200064
rect 194416 199504 194468 199510
rect 194416 199446 194468 199452
rect 194520 199442 194548 200058
rect 195150 199472 195206 199481
rect 194508 199436 194560 199442
rect 195150 199407 195206 199416
rect 194508 199378 194560 199384
rect 193862 196752 193918 196761
rect 193862 196687 193918 196696
rect 193126 178664 193182 178673
rect 193126 178599 193182 178608
rect 192576 130484 192628 130490
rect 192576 130426 192628 130432
rect 192576 118788 192628 118794
rect 192576 118730 192628 118736
rect 192588 86902 192616 118730
rect 193876 90370 193904 196687
rect 195164 190454 195192 199407
rect 195242 198792 195298 198801
rect 195242 198727 195298 198736
rect 195256 198694 195284 198727
rect 195244 198688 195296 198694
rect 195244 198630 195296 198636
rect 195440 198082 195468 220079
rect 195900 219434 195928 252554
rect 196716 247172 196768 247178
rect 196716 247114 196768 247120
rect 195978 235784 196034 235793
rect 195978 235719 196034 235728
rect 195992 234938 196020 235719
rect 196624 235272 196676 235278
rect 196624 235214 196676 235220
rect 195980 234932 196032 234938
rect 195980 234874 196032 234880
rect 196070 233336 196126 233345
rect 196070 233271 196126 233280
rect 196084 232529 196112 233271
rect 196070 232520 196126 232529
rect 196070 232455 196126 232464
rect 195888 219428 195940 219434
rect 195888 219370 195940 219376
rect 195428 198076 195480 198082
rect 195428 198018 195480 198024
rect 195164 190426 195284 190454
rect 194048 117360 194100 117366
rect 194048 117302 194100 117308
rect 193954 110528 194010 110537
rect 193954 110463 194010 110472
rect 193864 90364 193916 90370
rect 193864 90306 193916 90312
rect 192668 89004 192720 89010
rect 192668 88946 192720 88952
rect 192576 86896 192628 86902
rect 192576 86838 192628 86844
rect 192680 66230 192708 88946
rect 192668 66224 192720 66230
rect 192668 66166 192720 66172
rect 193968 63442 193996 110463
rect 194060 89729 194088 117302
rect 194046 89720 194102 89729
rect 194046 89655 194102 89664
rect 195256 86290 195284 190426
rect 196636 184210 196664 235214
rect 196728 214713 196756 247114
rect 196820 235929 196848 261462
rect 196898 254416 196954 254425
rect 196898 254351 196954 254360
rect 196806 235920 196862 235929
rect 196806 235855 196862 235864
rect 196912 232529 196940 254351
rect 197096 251705 197124 307090
rect 197188 280838 197216 311102
rect 197176 280832 197228 280838
rect 197176 280774 197228 280780
rect 197176 278724 197228 278730
rect 197176 278666 197228 278672
rect 197082 251696 197138 251705
rect 197082 251631 197084 251640
rect 197136 251631 197138 251640
rect 197084 251602 197136 251608
rect 197096 251571 197124 251602
rect 196898 232520 196954 232529
rect 196898 232455 196954 232464
rect 196714 214704 196770 214713
rect 196714 214639 196770 214648
rect 196716 213240 196768 213246
rect 196716 213182 196768 213188
rect 196728 193118 196756 213182
rect 196716 193112 196768 193118
rect 196716 193054 196768 193060
rect 196624 184204 196676 184210
rect 196624 184146 196676 184152
rect 197188 180169 197216 278666
rect 197280 276010 197308 349794
rect 198016 345030 198044 483103
rect 198844 463321 198872 551278
rect 205652 550905 205680 558991
rect 209780 558962 209832 558968
rect 209792 557534 209820 558962
rect 209792 557506 210464 557534
rect 207020 556232 207072 556238
rect 207020 556174 207072 556180
rect 205638 550896 205694 550905
rect 205638 550831 205694 550840
rect 199844 549364 199896 549370
rect 199844 549306 199896 549312
rect 199660 535424 199712 535430
rect 199660 535366 199712 535372
rect 199750 535392 199806 535401
rect 199672 530602 199700 535366
rect 199750 535327 199806 535336
rect 199764 533361 199792 535327
rect 199750 533352 199806 533361
rect 199750 533287 199806 533296
rect 199660 530596 199712 530602
rect 199660 530538 199712 530544
rect 199014 505200 199070 505209
rect 199014 505135 199070 505144
rect 198830 463312 198886 463321
rect 198830 463247 198886 463256
rect 198094 453520 198150 453529
rect 198094 453455 198150 453464
rect 198004 345024 198056 345030
rect 198004 344966 198056 344972
rect 198016 318889 198044 344966
rect 198108 329798 198136 453455
rect 198646 421696 198702 421705
rect 198646 421631 198702 421640
rect 198554 392320 198610 392329
rect 198554 392255 198610 392264
rect 198096 329792 198148 329798
rect 198096 329734 198148 329740
rect 198002 318880 198058 318889
rect 198002 318815 198058 318824
rect 198108 317665 198136 329734
rect 198094 317656 198150 317665
rect 198094 317591 198150 317600
rect 198108 316034 198136 317591
rect 198108 316006 198504 316034
rect 198370 307728 198426 307737
rect 198370 307663 198426 307672
rect 198384 306513 198412 307663
rect 198370 306504 198426 306513
rect 198370 306439 198426 306448
rect 197358 282432 197414 282441
rect 197358 282367 197414 282376
rect 197372 281586 197400 282367
rect 197360 281580 197412 281586
rect 197360 281522 197412 281528
rect 197360 281444 197412 281450
rect 197360 281386 197412 281392
rect 197372 280809 197400 281386
rect 197452 280832 197504 280838
rect 197358 280800 197414 280809
rect 197452 280774 197504 280780
rect 197358 280735 197414 280744
rect 197464 280265 197492 280774
rect 197450 280256 197506 280265
rect 197450 280191 197506 280200
rect 197358 279440 197414 279449
rect 197358 279375 197414 279384
rect 197372 278798 197400 279375
rect 197360 278792 197412 278798
rect 197360 278734 197412 278740
rect 197452 278724 197504 278730
rect 197452 278666 197504 278672
rect 197360 278656 197412 278662
rect 197464 278633 197492 278666
rect 197360 278598 197412 278604
rect 197450 278624 197506 278633
rect 197268 276004 197320 276010
rect 197268 275946 197320 275952
rect 197266 250064 197322 250073
rect 197266 249999 197322 250008
rect 197280 247178 197308 249999
rect 197268 247172 197320 247178
rect 197268 247114 197320 247120
rect 197372 245177 197400 278598
rect 197450 278559 197506 278568
rect 198384 278089 198412 306439
rect 198370 278080 198426 278089
rect 198370 278015 198426 278024
rect 197450 276720 197506 276729
rect 197450 276655 197506 276664
rect 197464 276078 197492 276655
rect 197452 276072 197504 276078
rect 197452 276014 197504 276020
rect 197544 276004 197596 276010
rect 197544 275946 197596 275952
rect 197556 275913 197584 275946
rect 197542 275904 197598 275913
rect 197542 275839 197598 275848
rect 197450 274544 197506 274553
rect 197450 274479 197506 274488
rect 197464 273494 197492 274479
rect 197452 273488 197504 273494
rect 197452 273430 197504 273436
rect 197452 273216 197504 273222
rect 197452 273158 197504 273164
rect 197464 272921 197492 273158
rect 197450 272912 197506 272921
rect 197450 272847 197506 272856
rect 197450 271552 197506 271561
rect 197450 271487 197506 271496
rect 197464 270570 197492 271487
rect 197452 270564 197504 270570
rect 197452 270506 197504 270512
rect 197450 270192 197506 270201
rect 197450 270127 197506 270136
rect 197464 269142 197492 270127
rect 197452 269136 197504 269142
rect 197452 269078 197504 269084
rect 197542 268832 197598 268841
rect 197542 268767 197598 268776
rect 197556 267782 197584 268767
rect 198280 268048 198332 268054
rect 198278 268016 198280 268025
rect 198332 268016 198334 268025
rect 198278 267951 198334 267960
rect 197544 267776 197596 267782
rect 197544 267718 197596 267724
rect 197452 267708 197504 267714
rect 197452 267650 197504 267656
rect 197464 266665 197492 267650
rect 197542 267200 197598 267209
rect 197542 267135 197544 267144
rect 197596 267135 197598 267144
rect 197544 267106 197596 267112
rect 197450 266656 197506 266665
rect 197450 266591 197506 266600
rect 197452 264920 197504 264926
rect 197452 264862 197504 264868
rect 197464 264489 197492 264862
rect 197450 264480 197506 264489
rect 197450 264415 197506 264424
rect 197450 263664 197506 263673
rect 197450 263599 197452 263608
rect 197504 263599 197506 263608
rect 197452 263570 197504 263576
rect 198476 262313 198504 316006
rect 198462 262304 198518 262313
rect 198462 262239 198518 262248
rect 198096 262200 198148 262206
rect 198096 262142 198148 262148
rect 197450 261488 197506 261497
rect 197450 261423 197506 261432
rect 197464 260914 197492 261423
rect 198108 260953 198136 262142
rect 198094 260944 198150 260953
rect 197452 260908 197504 260914
rect 198094 260879 198150 260888
rect 197452 260850 197504 260856
rect 197450 260128 197506 260137
rect 197450 260063 197506 260072
rect 197464 259486 197492 260063
rect 197452 259480 197504 259486
rect 197452 259422 197504 259428
rect 197450 259312 197506 259321
rect 197450 259247 197506 259256
rect 197464 258534 197492 259247
rect 197452 258528 197504 258534
rect 197452 258470 197504 258476
rect 197450 257952 197506 257961
rect 197450 257887 197506 257896
rect 197464 256834 197492 257887
rect 197542 257408 197598 257417
rect 197542 257343 197598 257352
rect 197452 256828 197504 256834
rect 197452 256770 197504 256776
rect 197556 256766 197584 257343
rect 197544 256760 197596 256766
rect 197544 256702 197596 256708
rect 197452 256692 197504 256698
rect 197452 256634 197504 256640
rect 197464 256601 197492 256634
rect 197450 256592 197506 256601
rect 197450 256527 197506 256536
rect 197452 255264 197504 255270
rect 197450 255232 197452 255241
rect 197504 255232 197506 255241
rect 197450 255167 197506 255176
rect 197910 253600 197966 253609
rect 197910 253535 197966 253544
rect 197924 253230 197952 253535
rect 197912 253224 197964 253230
rect 197912 253166 197964 253172
rect 198372 253224 198424 253230
rect 198372 253166 198424 253172
rect 197450 253056 197506 253065
rect 197450 252991 197506 253000
rect 197464 252618 197492 252991
rect 197452 252612 197504 252618
rect 197452 252554 197504 252560
rect 197450 250880 197506 250889
rect 197450 250815 197506 250824
rect 197464 249830 197492 250815
rect 197452 249824 197504 249830
rect 197452 249766 197504 249772
rect 197452 249552 197504 249558
rect 197450 249520 197452 249529
rect 197504 249520 197506 249529
rect 197450 249455 197506 249464
rect 197452 248736 197504 248742
rect 197450 248704 197452 248713
rect 197504 248704 197506 248713
rect 197450 248639 197506 248648
rect 197726 247888 197782 247897
rect 197726 247823 197782 247832
rect 197740 247110 197768 247823
rect 197728 247104 197780 247110
rect 197728 247046 197780 247052
rect 197358 245168 197414 245177
rect 197358 245103 197414 245112
rect 197372 244934 197400 245103
rect 197360 244928 197412 244934
rect 197360 244870 197412 244876
rect 197358 243808 197414 243817
rect 197358 243743 197414 243752
rect 197372 243030 197400 243743
rect 197360 243024 197412 243030
rect 197360 242966 197412 242972
rect 197912 240848 197964 240854
rect 197910 240816 197912 240825
rect 197964 240816 197966 240825
rect 197910 240751 197966 240760
rect 197268 231124 197320 231130
rect 197268 231066 197320 231072
rect 197280 230382 197308 231066
rect 197268 230376 197320 230382
rect 197268 230318 197320 230324
rect 197174 180160 197230 180169
rect 197174 180095 197230 180104
rect 196622 178800 196678 178809
rect 196622 178735 196678 178744
rect 195428 153264 195480 153270
rect 195428 153206 195480 153212
rect 195336 114640 195388 114646
rect 195336 114582 195388 114588
rect 195244 86284 195296 86290
rect 195244 86226 195296 86232
rect 195244 80708 195296 80714
rect 195244 80650 195296 80656
rect 193956 63436 194008 63442
rect 193956 63378 194008 63384
rect 192484 48272 192536 48278
rect 192484 48214 192536 48220
rect 195256 10402 195284 80650
rect 195348 51066 195376 114582
rect 195440 104174 195468 153206
rect 195428 104168 195480 104174
rect 195428 104110 195480 104116
rect 195336 51060 195388 51066
rect 195336 51002 195388 51008
rect 196636 13802 196664 178735
rect 196808 132524 196860 132530
rect 196808 132466 196860 132472
rect 196716 122936 196768 122942
rect 196716 122878 196768 122884
rect 196728 88330 196756 122878
rect 196820 100026 196848 132466
rect 197280 115161 197308 230318
rect 198096 217728 198148 217734
rect 198096 217670 198148 217676
rect 198004 216708 198056 216714
rect 198004 216650 198056 216656
rect 198016 186289 198044 216650
rect 198108 193866 198136 217670
rect 198384 195401 198412 253166
rect 198568 244361 198596 392255
rect 198660 252249 198688 421631
rect 198922 416800 198978 416809
rect 198922 416735 198978 416744
rect 198830 382528 198886 382537
rect 198830 382463 198886 382472
rect 198844 332586 198872 382463
rect 198936 376038 198964 416735
rect 198924 376032 198976 376038
rect 198924 375974 198976 375980
rect 199028 348430 199056 505135
rect 199384 375284 199436 375290
rect 199384 375226 199436 375232
rect 199016 348424 199068 348430
rect 199016 348366 199068 348372
rect 198832 332580 198884 332586
rect 198832 332522 198884 332528
rect 198740 331288 198792 331294
rect 198740 331230 198792 331236
rect 198752 314702 198780 331230
rect 198740 314696 198792 314702
rect 198740 314638 198792 314644
rect 198740 287088 198792 287094
rect 198792 287036 198872 287054
rect 198740 287030 198872 287036
rect 198752 287026 198872 287030
rect 198740 284368 198792 284374
rect 198740 284310 198792 284316
rect 198752 278225 198780 284310
rect 198844 283626 198872 287026
rect 198832 283620 198884 283626
rect 198832 283562 198884 283568
rect 198738 278216 198794 278225
rect 198738 278151 198794 278160
rect 198646 252240 198702 252249
rect 198646 252175 198702 252184
rect 198646 246528 198702 246537
rect 198646 246463 198702 246472
rect 198554 244352 198610 244361
rect 198554 244287 198610 244296
rect 198462 242176 198518 242185
rect 198462 242111 198518 242120
rect 198476 229809 198504 242111
rect 198660 238754 198688 246463
rect 198568 238726 198688 238754
rect 198568 231130 198596 238726
rect 199396 238066 199424 375226
rect 199856 374678 199884 549306
rect 201038 546680 201094 546689
rect 201038 546615 201094 546624
rect 201052 535401 201080 546615
rect 203614 541104 203670 541113
rect 203614 541039 203670 541048
rect 203628 535922 203656 541039
rect 205652 538214 205680 550831
rect 205652 538186 205772 538214
rect 203628 535894 204102 535922
rect 205744 535908 205772 538186
rect 207032 535922 207060 556174
rect 210436 535922 210464 557506
rect 212540 553444 212592 553450
rect 212540 553386 212592 553392
rect 207032 535894 207414 535922
rect 210436 535894 210910 535922
rect 212552 535908 212580 553386
rect 213932 535922 213960 565830
rect 231858 557560 231914 557569
rect 231914 557506 231992 557534
rect 231858 557495 231914 557504
rect 226984 552152 227036 552158
rect 226984 552094 227036 552100
rect 225326 545320 225382 545329
rect 225326 545255 225382 545264
rect 223672 543856 223724 543862
rect 223672 543798 223724 543804
rect 218704 542496 218756 542502
rect 218704 542438 218756 542444
rect 215852 539708 215904 539714
rect 215852 539650 215904 539656
rect 213932 535894 214222 535922
rect 215864 535908 215892 539650
rect 217506 538248 217562 538257
rect 217506 538183 217562 538192
rect 217520 535908 217548 538183
rect 218716 535922 218744 542438
rect 222474 538520 222530 538529
rect 222474 538455 222530 538464
rect 223210 538520 223266 538529
rect 223210 538455 223266 538464
rect 221094 538248 221150 538257
rect 221094 538183 221150 538192
rect 220820 536920 220872 536926
rect 220820 536862 220872 536868
rect 218716 535894 219190 535922
rect 220832 535908 220860 536862
rect 208674 535528 208730 535537
rect 202064 535486 202446 535514
rect 202064 535430 202092 535486
rect 208730 535486 209070 535514
rect 208674 535463 208730 535472
rect 202052 535424 202104 535430
rect 200394 535392 200450 535401
rect 201038 535392 201094 535401
rect 200450 535350 200790 535378
rect 200394 535327 200450 535336
rect 221108 535401 221136 538183
rect 222488 535908 222516 538455
rect 223224 538354 223252 538455
rect 223212 538348 223264 538354
rect 223212 538290 223264 538296
rect 223684 535922 223712 543798
rect 225340 535922 225368 545255
rect 226248 538280 226300 538286
rect 226248 538222 226300 538228
rect 223684 535894 224158 535922
rect 225340 535894 225814 535922
rect 202052 535366 202104 535372
rect 221094 535392 221150 535401
rect 201038 535327 201094 535336
rect 221094 535327 221150 535336
rect 226260 535294 226288 538222
rect 226996 535922 227024 552094
rect 229100 546508 229152 546514
rect 229100 546450 229152 546456
rect 226996 535894 227470 535922
rect 229112 535908 229140 546450
rect 230480 541068 230532 541074
rect 230480 541010 230532 541016
rect 230492 535922 230520 541010
rect 231964 535922 231992 557506
rect 233896 536858 233924 702714
rect 235184 702574 235212 703520
rect 267660 703050 267688 703520
rect 267648 703044 267700 703050
rect 267648 702986 267700 702992
rect 283852 702982 283880 703520
rect 281540 702976 281592 702982
rect 281540 702918 281592 702924
rect 283840 702976 283892 702982
rect 283840 702918 283892 702924
rect 273260 702908 273312 702914
rect 273260 702850 273312 702856
rect 276020 702908 276072 702914
rect 276020 702850 276072 702856
rect 235172 702568 235224 702574
rect 235172 702510 235224 702516
rect 264244 702568 264296 702574
rect 264244 702510 264296 702516
rect 259460 599004 259512 599010
rect 259460 598946 259512 598952
rect 255962 589384 256018 589393
rect 255962 589319 256018 589328
rect 241520 561808 241572 561814
rect 241520 561750 241572 561756
rect 241532 557534 241560 561750
rect 241532 557506 241928 557534
rect 235264 554872 235316 554878
rect 235264 554814 235316 554820
rect 240230 554840 240286 554849
rect 233884 536852 233936 536858
rect 233884 536794 233936 536800
rect 234068 536852 234120 536858
rect 234068 536794 234120 536800
rect 230492 535894 230782 535922
rect 231964 535894 232438 535922
rect 234080 535908 234108 536794
rect 235276 535922 235304 554814
rect 240230 554775 240286 554784
rect 238760 550724 238812 550730
rect 238760 550666 238812 550672
rect 237380 548004 237432 548010
rect 237380 547946 237432 547952
rect 235276 535894 235750 535922
rect 237392 535908 237420 547946
rect 238772 535922 238800 550666
rect 240244 535922 240272 554775
rect 241900 535922 241928 557506
rect 248512 556300 248564 556306
rect 248512 556242 248564 556248
rect 243542 556200 243598 556209
rect 243542 556135 243598 556144
rect 243556 535922 243584 556135
rect 247040 554804 247092 554810
rect 247040 554746 247092 554752
rect 245660 547188 245712 547194
rect 245660 547130 245712 547136
rect 238772 535894 239062 535922
rect 240244 535894 240718 535922
rect 241900 535894 242374 535922
rect 243556 535894 244030 535922
rect 245672 535908 245700 547130
rect 247052 535922 247080 554746
rect 248524 535922 248552 556242
rect 253938 550760 253994 550769
rect 253938 550695 253994 550704
rect 251824 549364 251876 549370
rect 251824 549306 251876 549312
rect 250628 539640 250680 539646
rect 250628 539582 250680 539588
rect 247052 535894 247342 535922
rect 248524 535894 248998 535922
rect 250640 535908 250668 539582
rect 251836 535922 251864 549306
rect 251836 535894 252310 535922
rect 253952 535908 253980 550695
rect 255318 545184 255374 545193
rect 255318 545119 255374 545128
rect 255332 535922 255360 545119
rect 255976 542502 256004 589319
rect 259472 557534 259500 598946
rect 264256 561678 264284 702510
rect 267740 561740 267792 561746
rect 267740 561682 267792 561688
rect 263600 561672 263652 561678
rect 263600 561614 263652 561620
rect 264244 561672 264296 561678
rect 264244 561614 264296 561620
rect 263612 560386 263640 561614
rect 263600 560380 263652 560386
rect 263600 560322 263652 560328
rect 259472 557506 260144 557534
rect 255964 542496 256016 542502
rect 255964 542438 256016 542444
rect 257344 542496 257396 542502
rect 257344 542438 257396 542444
rect 257356 535922 257384 542438
rect 258448 541000 258500 541006
rect 258448 540942 258500 540948
rect 255332 535894 255622 535922
rect 257278 535894 257384 535922
rect 258460 535922 258488 540942
rect 260116 535922 260144 557506
rect 261758 542736 261814 542745
rect 261758 542671 261814 542680
rect 261772 541686 261800 542671
rect 261760 541680 261812 541686
rect 261760 541622 261812 541628
rect 262218 541240 262274 541249
rect 262218 541175 262274 541184
rect 258460 535894 258934 535922
rect 260116 535894 260590 535922
rect 262232 535908 262260 541175
rect 263612 535922 263640 560322
rect 267752 557534 267780 561682
rect 268384 557592 268436 557598
rect 268384 557534 268436 557540
rect 267752 557506 268332 557534
rect 266728 542428 266780 542434
rect 266728 542370 266780 542376
rect 265530 538520 265586 538529
rect 265530 538455 265586 538464
rect 263612 535894 263902 535922
rect 265544 535908 265572 538455
rect 266740 535922 266768 542370
rect 268304 538214 268332 557506
rect 268396 539578 268424 557534
rect 270500 552084 270552 552090
rect 270500 552026 270552 552032
rect 268384 539572 268436 539578
rect 268384 539514 268436 539520
rect 268304 538186 268608 538214
rect 268580 535922 268608 538186
rect 270512 535922 270540 552026
rect 273272 546689 273300 702850
rect 273258 546680 273314 546689
rect 273258 546615 273314 546624
rect 270684 543788 270736 543794
rect 270684 543730 270736 543736
rect 270696 539617 270724 543730
rect 270682 539608 270738 539617
rect 273272 539578 273300 546615
rect 273994 539608 274050 539617
rect 270682 539543 270738 539552
rect 272340 539572 272392 539578
rect 272340 539514 272392 539520
rect 273260 539572 273312 539578
rect 273994 539543 274050 539552
rect 275652 539572 275704 539578
rect 273260 539514 273312 539520
rect 266740 535894 267214 535922
rect 268580 535894 269054 535922
rect 270512 535894 270710 535922
rect 272352 535908 272380 539514
rect 274008 535908 274036 539543
rect 275652 539514 275704 539520
rect 275664 535908 275692 539514
rect 276032 535673 276060 702850
rect 281552 557534 281580 702918
rect 300136 702642 300164 703520
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 300124 702636 300176 702642
rect 300124 702578 300176 702584
rect 327724 700324 327776 700330
rect 327724 700266 327776 700272
rect 320180 568608 320232 568614
rect 320180 568550 320232 568556
rect 311900 567248 311952 567254
rect 311900 567190 311952 567196
rect 291200 564460 291252 564466
rect 291200 564402 291252 564408
rect 288440 558952 288492 558958
rect 288440 558894 288492 558900
rect 281552 557506 281856 557534
rect 278044 549296 278096 549302
rect 278044 549238 278096 549244
rect 278056 539578 278084 549238
rect 280618 539880 280674 539889
rect 280618 539815 280674 539824
rect 278044 539572 278096 539578
rect 278044 539514 278096 539520
rect 278964 539572 279016 539578
rect 278964 539514 279016 539520
rect 278976 535908 279004 539514
rect 280632 535908 280660 539815
rect 281828 535922 281856 557506
rect 287060 553512 287112 553518
rect 287060 553454 287112 553460
rect 284300 547936 284352 547942
rect 284300 547878 284352 547884
rect 283470 542600 283526 542609
rect 283470 542535 283526 542544
rect 283484 535922 283512 542535
rect 284312 538214 284340 547878
rect 284312 538186 285168 538214
rect 285140 535922 285168 538186
rect 287072 535922 287100 553454
rect 288452 535922 288480 558894
rect 291212 557534 291240 564402
rect 291212 557506 291792 557534
rect 290094 552120 290150 552129
rect 290094 552055 290150 552064
rect 290108 535922 290136 552055
rect 291764 535922 291792 557506
rect 304998 549400 305054 549409
rect 304998 549335 305054 549344
rect 295338 546680 295394 546689
rect 295338 546615 295394 546624
rect 295352 535922 295380 546615
rect 300032 545148 300084 545154
rect 300032 545090 300084 545096
rect 298374 544096 298430 544105
rect 298374 544031 298430 544040
rect 297180 538280 297232 538286
rect 297180 538222 297232 538228
rect 281828 535894 282302 535922
rect 283484 535894 283958 535922
rect 285140 535894 285614 535922
rect 287072 535894 287270 535922
rect 288452 535894 288926 535922
rect 290108 535894 290582 535922
rect 291764 535894 292238 535922
rect 295352 535894 295550 535922
rect 297192 535908 297220 538222
rect 298388 535922 298416 544031
rect 300044 535922 300072 545090
rect 305012 535922 305040 549335
rect 309968 545148 310020 545154
rect 309968 545090 310020 545096
rect 306654 543960 306710 543969
rect 306654 543895 306710 543904
rect 306668 535922 306696 543895
rect 309980 535922 310008 545090
rect 311912 535922 311940 567190
rect 316592 543788 316644 543794
rect 316592 543730 316644 543736
rect 315396 539708 315448 539714
rect 315396 539650 315448 539656
rect 298388 535894 298862 535922
rect 300044 535894 300518 535922
rect 305012 535894 305486 535922
rect 306668 535894 307142 535922
rect 309980 535894 310454 535922
rect 311912 535894 312110 535922
rect 315408 535908 315436 539650
rect 316604 535922 316632 543730
rect 318246 541240 318302 541249
rect 318246 541175 318302 541184
rect 318260 535922 318288 541175
rect 320192 535922 320220 568550
rect 327736 545630 327764 700266
rect 331232 551342 331260 702986
rect 348804 700330 348832 703520
rect 351920 702976 351972 702982
rect 351920 702918 351972 702924
rect 349804 702840 349856 702846
rect 349804 702782 349856 702788
rect 348792 700324 348844 700330
rect 348792 700266 348844 700272
rect 349816 596222 349844 702782
rect 349804 596216 349856 596222
rect 349804 596158 349856 596164
rect 341524 569968 341576 569974
rect 341524 569910 341576 569916
rect 331220 551336 331272 551342
rect 331220 551278 331272 551284
rect 328458 547904 328514 547913
rect 328458 547839 328514 547848
rect 324320 545624 324372 545630
rect 324320 545566 324372 545572
rect 324872 545624 324924 545630
rect 324872 545566 324924 545572
rect 327724 545624 327776 545630
rect 327724 545566 327776 545572
rect 324332 545222 324360 545566
rect 324320 545216 324372 545222
rect 324320 545158 324372 545164
rect 323582 541512 323638 541521
rect 323582 541447 323638 541456
rect 322018 539744 322074 539753
rect 322018 539679 322074 539688
rect 316604 535894 317078 535922
rect 318260 535894 318734 535922
rect 320192 535894 320390 535922
rect 322032 535908 322060 539679
rect 323596 539646 323624 541447
rect 323584 539640 323636 539646
rect 323584 539582 323636 539588
rect 323596 538214 323624 539582
rect 323596 538186 323716 538214
rect 323688 535908 323716 538186
rect 324884 535922 324912 545566
rect 327080 545216 327132 545222
rect 327080 545158 327132 545164
rect 327092 538214 327120 545158
rect 327092 538186 327212 538214
rect 324884 535894 325358 535922
rect 327184 535908 327212 538186
rect 328472 535922 328500 547839
rect 339958 546544 340014 546553
rect 339958 546479 340014 546488
rect 338304 541000 338356 541006
rect 338304 540942 338356 540948
rect 337106 538520 337162 538529
rect 337106 538455 337162 538464
rect 335450 537160 335506 537169
rect 335450 537095 335506 537104
rect 333794 537024 333850 537033
rect 333794 536959 333850 536968
rect 330484 536920 330536 536926
rect 330484 536862 330536 536868
rect 328472 535894 328854 535922
rect 330496 535908 330524 536862
rect 333808 535908 333836 536959
rect 335464 535908 335492 537095
rect 337120 535908 337148 538455
rect 338316 535922 338344 540942
rect 339972 535922 340000 546479
rect 341536 539578 341564 569910
rect 349816 557534 349844 596158
rect 351932 587926 351960 702918
rect 364996 702710 365024 703520
rect 397472 702794 397500 703520
rect 397380 702778 397500 702794
rect 397368 702772 397500 702778
rect 397420 702766 397500 702772
rect 397368 702714 397420 702720
rect 364984 702704 365036 702710
rect 364984 702646 365036 702652
rect 381544 702704 381596 702710
rect 381544 702646 381596 702652
rect 356152 702636 356204 702642
rect 356152 702578 356204 702584
rect 360844 702636 360896 702642
rect 360844 702578 360896 702584
rect 351920 587920 351972 587926
rect 351920 587862 351972 587868
rect 349816 557506 350028 557534
rect 348238 542464 348294 542473
rect 348238 542399 348294 542408
rect 341524 539572 341576 539578
rect 341524 539514 341576 539520
rect 343732 539572 343784 539578
rect 343732 539514 343784 539520
rect 345388 539572 345440 539578
rect 345388 539514 345440 539520
rect 342076 536852 342128 536858
rect 342076 536794 342128 536800
rect 338316 535894 338790 535922
rect 339972 535894 340446 535922
rect 342088 535908 342116 536794
rect 343744 535908 343772 539514
rect 345400 535908 345428 539514
rect 347044 538348 347096 538354
rect 347044 538290 347096 538296
rect 347056 535908 347084 538290
rect 348252 535922 348280 542399
rect 350000 541113 350028 557506
rect 349986 541104 350042 541113
rect 349986 541039 350042 541048
rect 350000 539578 350028 541039
rect 349988 539572 350040 539578
rect 349988 539514 350040 539520
rect 350356 538280 350408 538286
rect 350356 538222 350408 538228
rect 348252 535894 348726 535922
rect 350368 535908 350396 538222
rect 351932 538214 351960 587862
rect 356060 542496 356112 542502
rect 356058 542464 356060 542473
rect 356112 542464 356114 542473
rect 356058 542399 356114 542408
rect 351932 538186 352052 538214
rect 352024 535908 352052 538186
rect 353666 536888 353722 536897
rect 353666 536823 353722 536832
rect 353680 535908 353708 536823
rect 308402 535800 308458 535809
rect 308458 535758 308798 535786
rect 308402 535735 308458 535744
rect 276018 535664 276074 535673
rect 276018 535599 276074 535608
rect 276938 535664 276994 535673
rect 276994 535622 277334 535650
rect 276938 535599 276994 535608
rect 313372 535560 313424 535566
rect 304078 535528 304134 535537
rect 293512 535498 293894 535514
rect 293500 535492 293894 535498
rect 293552 535486 293894 535492
rect 302174 535498 302372 535514
rect 302174 535492 302384 535498
rect 302174 535486 302332 535492
rect 293500 535434 293552 535440
rect 303830 535486 304078 535514
rect 332416 535560 332468 535566
rect 313424 535508 313766 535514
rect 313372 535502 313766 535508
rect 313384 535486 313766 535502
rect 332166 535508 332416 535514
rect 332166 535502 332468 535508
rect 332166 535486 332456 535502
rect 304078 535463 304134 535472
rect 302332 535434 302384 535440
rect 355350 535350 355640 535378
rect 355612 535294 355640 535350
rect 226248 535288 226300 535294
rect 226248 535230 226300 535236
rect 355600 535288 355652 535294
rect 355600 535230 355652 535236
rect 356164 519738 356192 702578
rect 357440 563100 357492 563106
rect 357440 563042 357492 563048
rect 357348 543720 357400 543726
rect 357348 543662 357400 543668
rect 357360 542502 357388 543662
rect 357348 542496 357400 542502
rect 357348 542438 357400 542444
rect 356242 538384 356298 538393
rect 356242 538319 356298 538328
rect 356256 520010 356284 538319
rect 357452 522345 357480 563042
rect 359004 560312 359056 560318
rect 359004 560254 359056 560260
rect 357622 543824 357678 543833
rect 357622 543759 357678 543768
rect 357530 540152 357586 540161
rect 357530 540087 357586 540096
rect 357438 522336 357494 522345
rect 357438 522271 357494 522280
rect 356256 519982 356468 520010
rect 356334 519888 356390 519897
rect 356334 519823 356390 519832
rect 356348 519738 356376 519823
rect 356164 519710 356376 519738
rect 356440 509234 356468 519982
rect 357544 512689 357572 540087
rect 357636 534721 357664 543759
rect 358820 538348 358872 538354
rect 358820 538290 358872 538296
rect 357622 534712 357678 534721
rect 357622 534647 357678 534656
rect 358726 532128 358782 532137
rect 358726 532063 358782 532072
rect 358740 532030 358768 532063
rect 358728 532024 358780 532030
rect 358728 531966 358780 531972
rect 358726 529680 358782 529689
rect 358726 529615 358782 529624
rect 358740 528630 358768 529615
rect 358728 528624 358780 528630
rect 358728 528566 358780 528572
rect 358726 527232 358782 527241
rect 358726 527167 358728 527176
rect 358780 527167 358782 527176
rect 358728 527138 358780 527144
rect 358726 524784 358782 524793
rect 358726 524719 358782 524728
rect 358740 524482 358768 524719
rect 358728 524476 358780 524482
rect 358728 524418 358780 524424
rect 358726 522336 358782 522345
rect 358726 522271 358782 522280
rect 358740 520946 358768 522271
rect 358728 520940 358780 520946
rect 358728 520882 358780 520888
rect 358634 519888 358690 519897
rect 358634 519823 358690 519832
rect 358648 518974 358676 519823
rect 358636 518968 358688 518974
rect 358636 518910 358688 518916
rect 358726 517440 358782 517449
rect 358726 517375 358782 517384
rect 358740 516186 358768 517375
rect 358728 516180 358780 516186
rect 358728 516122 358780 516128
rect 357530 512680 357586 512689
rect 357530 512615 357586 512624
rect 358082 510096 358138 510105
rect 358082 510031 358138 510040
rect 356256 509206 356468 509234
rect 356256 490929 356284 509206
rect 356242 490920 356298 490929
rect 356242 490855 356298 490864
rect 357898 482896 357954 482905
rect 357898 482831 357954 482840
rect 357912 481710 357940 482831
rect 357900 481704 357952 481710
rect 357900 481646 357952 481652
rect 357898 478000 357954 478009
rect 357898 477935 357954 477944
rect 357912 477562 357940 477935
rect 357900 477556 357952 477562
rect 357900 477498 357952 477504
rect 358096 473346 358124 510031
rect 358726 507648 358782 507657
rect 358726 507583 358782 507592
rect 358740 506530 358768 507583
rect 358728 506524 358780 506530
rect 358728 506466 358780 506472
rect 358726 505200 358782 505209
rect 358726 505135 358728 505144
rect 358780 505135 358782 505144
rect 358728 505106 358780 505112
rect 358726 502752 358782 502761
rect 358726 502687 358782 502696
rect 358740 502450 358768 502687
rect 358728 502444 358780 502450
rect 358728 502386 358780 502392
rect 358726 497856 358782 497865
rect 358726 497791 358782 497800
rect 358636 496800 358688 496806
rect 358636 496742 358688 496748
rect 358648 495553 358676 496742
rect 358634 495544 358690 495553
rect 358634 495479 358690 495488
rect 358740 494766 358768 497791
rect 358728 494760 358780 494766
rect 358728 494702 358780 494708
rect 358726 492960 358782 492969
rect 358726 492895 358782 492904
rect 358740 492726 358768 492895
rect 358728 492720 358780 492726
rect 358728 492662 358780 492668
rect 358726 487792 358782 487801
rect 358726 487727 358782 487736
rect 358740 487218 358768 487727
rect 358728 487212 358780 487218
rect 358728 487154 358780 487160
rect 358174 485344 358230 485353
rect 358174 485279 358230 485288
rect 358188 484430 358216 485279
rect 358176 484424 358228 484430
rect 358176 484366 358228 484372
rect 358726 475552 358782 475561
rect 358726 475487 358782 475496
rect 358740 474774 358768 475487
rect 358728 474768 358780 474774
rect 358728 474710 358780 474716
rect 358084 473340 358136 473346
rect 358084 473282 358136 473288
rect 358726 473104 358782 473113
rect 358726 473039 358782 473048
rect 358740 472054 358768 473039
rect 358728 472048 358780 472054
rect 358728 471990 358780 471996
rect 358726 470656 358782 470665
rect 358726 470591 358728 470600
rect 358780 470591 358782 470600
rect 358728 470562 358780 470568
rect 356242 467936 356298 467945
rect 356242 467871 356298 467880
rect 356256 451274 356284 467871
rect 358726 465760 358782 465769
rect 358726 465695 358782 465704
rect 358740 465118 358768 465695
rect 358728 465112 358780 465118
rect 358728 465054 358780 465060
rect 358634 463312 358690 463321
rect 358634 463247 358690 463256
rect 358648 462398 358676 463247
rect 358636 462392 358688 462398
rect 358636 462334 358688 462340
rect 358726 460864 358782 460873
rect 358726 460799 358782 460808
rect 358740 459610 358768 460799
rect 358728 459604 358780 459610
rect 358728 459546 358780 459552
rect 357438 458416 357494 458425
rect 357438 458351 357494 458360
rect 356164 451246 356284 451274
rect 201314 377632 201370 377641
rect 199948 377590 200054 377618
rect 199948 375290 199976 377590
rect 201314 377567 201370 377576
rect 201512 377590 201710 377618
rect 202892 377590 203366 377618
rect 204272 377590 205022 377618
rect 200026 376544 200082 376553
rect 200026 376479 200082 376488
rect 200040 375306 200068 376479
rect 200304 375692 200356 375698
rect 200304 375634 200356 375640
rect 199936 375284 199988 375290
rect 200040 375278 200160 375306
rect 199936 375226 199988 375232
rect 199844 374672 199896 374678
rect 199844 374614 199896 374620
rect 199476 336048 199528 336054
rect 199476 335990 199528 335996
rect 199488 305114 199516 335990
rect 199568 318096 199620 318102
rect 199568 318038 199620 318044
rect 199580 307834 199608 318038
rect 200132 310457 200160 375278
rect 200210 367840 200266 367849
rect 200210 367775 200266 367784
rect 200118 310448 200174 310457
rect 200118 310383 200174 310392
rect 199568 307828 199620 307834
rect 199568 307770 199620 307776
rect 200028 307828 200080 307834
rect 200028 307770 200080 307776
rect 199476 305108 199528 305114
rect 199476 305050 199528 305056
rect 199568 290828 199620 290834
rect 199568 290770 199620 290776
rect 199476 283960 199528 283966
rect 199476 283902 199528 283908
rect 199488 273970 199516 283902
rect 199476 273964 199528 273970
rect 199476 273906 199528 273912
rect 199474 272368 199530 272377
rect 199474 272303 199530 272312
rect 199488 250481 199516 272303
rect 199580 271182 199608 290770
rect 200040 288522 200068 307770
rect 200120 305108 200172 305114
rect 200120 305050 200172 305056
rect 200028 288516 200080 288522
rect 200028 288458 200080 288464
rect 200132 285326 200160 305050
rect 200120 285320 200172 285326
rect 200120 285262 200172 285268
rect 200224 283914 200252 367775
rect 200316 298178 200344 375634
rect 201328 373994 201356 377567
rect 201328 373966 201448 373994
rect 201420 362273 201448 373966
rect 201406 362264 201462 362273
rect 201406 362199 201462 362208
rect 200488 319524 200540 319530
rect 200488 319466 200540 319472
rect 200304 298172 200356 298178
rect 200304 298114 200356 298120
rect 200394 291952 200450 291961
rect 200394 291887 200450 291896
rect 200408 284172 200436 291887
rect 200500 291009 200528 319466
rect 201408 305108 201460 305114
rect 201408 305050 201460 305056
rect 201420 305017 201448 305050
rect 201406 305008 201462 305017
rect 201406 304943 201462 304952
rect 201316 298784 201368 298790
rect 201316 298726 201368 298732
rect 201328 298178 201356 298726
rect 201316 298172 201368 298178
rect 201316 298114 201368 298120
rect 200486 291000 200542 291009
rect 200486 290935 200542 290944
rect 201512 290834 201540 377590
rect 201590 377496 201646 377505
rect 201590 377431 201646 377440
rect 201604 364750 201632 377431
rect 202234 376000 202290 376009
rect 202234 375935 202290 375944
rect 201592 364744 201644 364750
rect 201592 364686 201644 364692
rect 202144 364744 202196 364750
rect 202144 364686 202196 364692
rect 201604 364478 201632 364686
rect 201592 364472 201644 364478
rect 201592 364414 201644 364420
rect 202156 311914 202184 364686
rect 202248 363662 202276 375935
rect 202892 363769 202920 377590
rect 203616 377460 203668 377466
rect 203616 377402 203668 377408
rect 203524 365832 203576 365838
rect 203524 365774 203576 365780
rect 202878 363760 202934 363769
rect 202878 363695 202934 363704
rect 202236 363656 202288 363662
rect 202236 363598 202288 363604
rect 202236 362296 202288 362302
rect 202236 362238 202288 362244
rect 202248 332382 202276 362238
rect 202880 337408 202932 337414
rect 202880 337350 202932 337356
rect 202328 332580 202380 332586
rect 202328 332522 202380 332528
rect 202788 332580 202840 332586
rect 202788 332522 202840 332528
rect 202236 332376 202288 332382
rect 202236 332318 202288 332324
rect 202144 311908 202196 311914
rect 202144 311850 202196 311856
rect 202340 306374 202368 332522
rect 202800 332382 202828 332522
rect 202788 332376 202840 332382
rect 202788 332318 202840 332324
rect 202800 318850 202828 332318
rect 202788 318844 202840 318850
rect 202788 318786 202840 318792
rect 202248 306346 202368 306374
rect 202248 302326 202276 306346
rect 202236 302320 202288 302326
rect 202236 302262 202288 302268
rect 202248 294098 202276 302262
rect 202236 294092 202288 294098
rect 202236 294034 202288 294040
rect 202142 291408 202198 291417
rect 202142 291343 202198 291352
rect 201500 290828 201552 290834
rect 201500 290770 201552 290776
rect 201684 288516 201736 288522
rect 201684 288458 201736 288464
rect 201408 285864 201460 285870
rect 201408 285806 201460 285812
rect 200948 285320 201000 285326
rect 200948 285262 201000 285268
rect 200960 284186 200988 285262
rect 200960 284158 201342 284186
rect 200486 284064 200542 284073
rect 200542 284022 200790 284050
rect 200486 283999 200542 284008
rect 201420 283966 201448 285806
rect 201696 284172 201724 288458
rect 202156 284889 202184 291343
rect 202142 284880 202198 284889
rect 202142 284815 202198 284824
rect 202248 284172 202276 294034
rect 202800 284172 202828 318786
rect 202892 291961 202920 337350
rect 203536 297498 203564 365774
rect 203628 322998 203656 377402
rect 203616 322992 203668 322998
rect 203616 322934 203668 322940
rect 203524 297492 203576 297498
rect 203524 297434 203576 297440
rect 203628 293185 203656 322934
rect 204272 307086 204300 377590
rect 205730 376136 205786 376145
rect 205730 376071 205786 376080
rect 204352 376032 204404 376038
rect 204352 375974 204404 375980
rect 204364 307154 204392 375974
rect 205640 373380 205692 373386
rect 205640 373322 205692 373328
rect 204904 363792 204956 363798
rect 204904 363734 204956 363740
rect 204916 315382 204944 363734
rect 205652 347750 205680 373322
rect 205744 353326 205772 376071
rect 206664 375358 206692 377604
rect 208320 375358 208348 377604
rect 209792 377590 209990 377618
rect 211172 377590 211646 377618
rect 205824 375352 205876 375358
rect 205824 375294 205876 375300
rect 206652 375352 206704 375358
rect 206652 375294 206704 375300
rect 207020 375352 207072 375358
rect 207020 375294 207072 375300
rect 208308 375352 208360 375358
rect 208308 375294 208360 375300
rect 205836 366489 205864 375294
rect 207032 370598 207060 375294
rect 207112 374672 207164 374678
rect 207112 374614 207164 374620
rect 209044 374672 209096 374678
rect 209044 374614 209096 374620
rect 207020 370592 207072 370598
rect 207020 370534 207072 370540
rect 207032 370326 207060 370534
rect 207020 370320 207072 370326
rect 207020 370262 207072 370268
rect 205822 366480 205878 366489
rect 205822 366415 205878 366424
rect 207124 358562 207152 374614
rect 208308 370320 208360 370326
rect 208360 370268 208440 370274
rect 208308 370262 208440 370268
rect 208320 370246 208440 370262
rect 208412 366353 208440 370246
rect 208398 366344 208454 366353
rect 208398 366279 208454 366288
rect 207112 358556 207164 358562
rect 207112 358498 207164 358504
rect 207664 358556 207716 358562
rect 207664 358498 207716 358504
rect 207676 357542 207704 358498
rect 207664 357536 207716 357542
rect 207664 357478 207716 357484
rect 205732 353320 205784 353326
rect 205732 353262 205784 353268
rect 206284 353320 206336 353326
rect 206284 353262 206336 353268
rect 205640 347744 205692 347750
rect 205640 347686 205692 347692
rect 204996 325712 205048 325718
rect 204996 325654 205048 325660
rect 205008 317422 205036 325654
rect 204996 317416 205048 317422
rect 204996 317358 205048 317364
rect 204904 315376 204956 315382
rect 204904 315318 204956 315324
rect 204352 307148 204404 307154
rect 204352 307090 204404 307096
rect 204260 307080 204312 307086
rect 204260 307022 204312 307028
rect 204260 297560 204312 297566
rect 204260 297502 204312 297508
rect 203614 293176 203670 293185
rect 203614 293111 203670 293120
rect 202878 291952 202934 291961
rect 202878 291887 202934 291896
rect 204272 289785 204300 297502
rect 204902 295488 204958 295497
rect 204902 295423 204958 295432
rect 203154 289776 203210 289785
rect 203154 289711 203210 289720
rect 204258 289776 204314 289785
rect 204258 289711 204314 289720
rect 203168 284172 203196 289711
rect 204272 289241 204300 289711
rect 204258 289232 204314 289241
rect 204258 289167 204314 289176
rect 204258 285016 204314 285025
rect 204258 284951 204314 284960
rect 203340 284300 203392 284306
rect 203340 284242 203392 284248
rect 203352 284186 203380 284242
rect 203352 284158 203734 284186
rect 204272 284172 204300 284951
rect 204916 284889 204944 295423
rect 205008 285802 205036 317358
rect 206296 296721 206324 353262
rect 206376 347744 206428 347750
rect 206376 347686 206428 347692
rect 206388 346458 206416 347686
rect 206376 346452 206428 346458
rect 206376 346394 206428 346400
rect 206388 315353 206416 346394
rect 206468 326460 206520 326466
rect 206468 326402 206520 326408
rect 206374 315344 206430 315353
rect 206374 315279 206430 315288
rect 206480 298081 206508 326402
rect 207676 305833 207704 357478
rect 207754 338736 207810 338745
rect 207754 338671 207810 338680
rect 207768 306474 207796 338671
rect 208124 316124 208176 316130
rect 208124 316066 208176 316072
rect 207756 306468 207808 306474
rect 207756 306410 207808 306416
rect 207662 305824 207718 305833
rect 207662 305759 207718 305768
rect 206466 298072 206522 298081
rect 206466 298007 206522 298016
rect 207570 298072 207626 298081
rect 207570 298007 207626 298016
rect 206650 297528 206706 297537
rect 206650 297463 206706 297472
rect 206282 296712 206338 296721
rect 206282 296647 206338 296656
rect 205548 285864 205600 285870
rect 205548 285806 205600 285812
rect 204996 285796 205048 285802
rect 204996 285738 205048 285744
rect 205178 285696 205234 285705
rect 205178 285631 205234 285640
rect 204902 284880 204958 284889
rect 204902 284815 204958 284824
rect 204628 284368 204680 284374
rect 204628 284310 204680 284316
rect 204640 284172 204668 284310
rect 200132 283886 200252 283914
rect 201408 283960 201460 283966
rect 201408 283902 201460 283908
rect 205192 283914 205220 285631
rect 205560 284172 205588 285806
rect 206664 284374 206692 297463
rect 207584 296857 207612 298007
rect 207570 296848 207626 296857
rect 207570 296783 207626 296792
rect 207020 285796 207072 285802
rect 207020 285738 207072 285744
rect 206652 284368 206704 284374
rect 206098 284336 206154 284345
rect 206652 284310 206704 284316
rect 206098 284271 206154 284280
rect 206112 284172 206140 284271
rect 206664 284172 206692 284310
rect 207032 284172 207060 285738
rect 207584 284172 207612 296783
rect 207768 291145 207796 306410
rect 207754 291136 207810 291145
rect 207754 291071 207810 291080
rect 208136 284172 208164 316066
rect 208492 309188 208544 309194
rect 208492 309130 208544 309136
rect 208504 284172 208532 309130
rect 209056 306374 209084 374614
rect 209134 369200 209190 369209
rect 209134 369135 209190 369144
rect 209148 337482 209176 369135
rect 209792 365838 209820 377590
rect 209780 365832 209832 365838
rect 209780 365774 209832 365780
rect 211172 355366 211200 377590
rect 213288 374678 213316 377604
rect 214576 377590 214958 377618
rect 215312 377590 216614 377618
rect 213276 374672 213328 374678
rect 213276 374614 213328 374620
rect 214576 374105 214604 377590
rect 215206 375184 215262 375193
rect 215206 375119 215262 375128
rect 214562 374096 214618 374105
rect 213276 374060 213328 374066
rect 214562 374031 214618 374040
rect 213276 374002 213328 374008
rect 213184 367804 213236 367810
rect 213184 367746 213236 367752
rect 211160 355360 211212 355366
rect 211160 355302 211212 355308
rect 211894 351248 211950 351257
rect 211894 351183 211950 351192
rect 209780 345704 209832 345710
rect 209780 345646 209832 345652
rect 209136 337476 209188 337482
rect 209136 337418 209188 337424
rect 209134 327856 209190 327865
rect 209134 327791 209190 327800
rect 208964 306346 209084 306374
rect 209148 306374 209176 327791
rect 209792 316130 209820 345646
rect 211804 341556 211856 341562
rect 211804 341498 211856 341504
rect 210424 319456 210476 319462
rect 210424 319398 210476 319404
rect 209780 316124 209832 316130
rect 209780 316066 209832 316072
rect 209228 311908 209280 311914
rect 209228 311850 209280 311856
rect 209240 309194 209268 311850
rect 209228 309188 209280 309194
rect 209228 309130 209280 309136
rect 209412 306400 209464 306406
rect 209148 306348 209412 306374
rect 209148 306346 209464 306348
rect 208964 304298 208992 306346
rect 209412 306342 209464 306346
rect 208952 304292 209004 304298
rect 208952 304234 209004 304240
rect 209044 304292 209096 304298
rect 209044 304234 209096 304240
rect 209056 296002 209084 304234
rect 209044 295996 209096 296002
rect 209044 295938 209096 295944
rect 209056 284172 209084 295938
rect 209424 284172 209452 306342
rect 210436 289950 210464 319398
rect 210974 317384 211030 317393
rect 210974 317319 211030 317328
rect 210988 316130 211016 317319
rect 210976 316124 211028 316130
rect 210976 316066 211028 316072
rect 210606 310584 210662 310593
rect 210606 310519 210662 310528
rect 210424 289944 210476 289950
rect 210424 289886 210476 289892
rect 209962 289096 210018 289105
rect 209962 289031 210018 289040
rect 209976 284172 210004 289031
rect 210436 284186 210464 289886
rect 210620 289105 210648 310519
rect 211434 305688 211490 305697
rect 211434 305623 211490 305632
rect 211448 303793 211476 305623
rect 211434 303784 211490 303793
rect 211434 303719 211490 303728
rect 210606 289096 210662 289105
rect 210606 289031 210662 289040
rect 210884 285728 210936 285734
rect 210884 285670 210936 285676
rect 210436 284158 210542 284186
rect 210896 284172 210924 285670
rect 211448 284172 211476 303719
rect 211816 285734 211844 341498
rect 211908 338745 211936 351183
rect 211894 338736 211950 338745
rect 211894 338671 211950 338680
rect 213196 314945 213224 367746
rect 213288 359553 213316 374002
rect 213274 359544 213330 359553
rect 213274 359479 213330 359488
rect 213276 339584 213328 339590
rect 213276 339526 213328 339532
rect 213288 318102 213316 339526
rect 214576 326398 214604 374031
rect 215116 327820 215168 327826
rect 215116 327762 215168 327768
rect 214564 326392 214616 326398
rect 214564 326334 214616 326340
rect 214564 325644 214616 325650
rect 214564 325586 214616 325592
rect 214576 325174 214604 325586
rect 215128 325174 215156 327762
rect 214564 325168 214616 325174
rect 214564 325110 214616 325116
rect 215116 325168 215168 325174
rect 215116 325110 215168 325116
rect 213368 319456 213420 319462
rect 213368 319398 213420 319404
rect 213276 318096 213328 318102
rect 213276 318038 213328 318044
rect 213182 314936 213238 314945
rect 213182 314871 213238 314880
rect 212724 305108 212776 305114
rect 212724 305050 212776 305056
rect 212736 302938 212764 305050
rect 212724 302932 212776 302938
rect 212724 302874 212776 302880
rect 212354 292768 212410 292777
rect 212354 292703 212410 292712
rect 211986 289776 212042 289785
rect 211986 289711 212042 289720
rect 212000 288561 212028 289711
rect 211986 288552 212042 288561
rect 211986 288487 212042 288496
rect 211804 285728 211856 285734
rect 211804 285670 211856 285676
rect 212000 284172 212028 288487
rect 212368 284172 212396 292703
rect 213196 289785 213224 314871
rect 213380 307057 213408 319398
rect 213366 307048 213422 307057
rect 213366 306983 213422 306992
rect 213380 306374 213408 306983
rect 214576 306374 214604 325110
rect 214656 323060 214708 323066
rect 214656 323002 214708 323008
rect 214668 308689 214696 323002
rect 214654 308680 214710 308689
rect 214654 308615 214710 308624
rect 213380 306346 213500 306374
rect 214576 306346 214788 306374
rect 213182 289776 213238 289785
rect 213182 289711 213238 289720
rect 212908 285796 212960 285802
rect 212908 285738 212960 285744
rect 212920 284172 212948 285738
rect 213472 284172 213500 306346
rect 214760 299577 214788 306346
rect 215220 304298 215248 375119
rect 215312 350441 215340 377590
rect 218256 376825 218284 377604
rect 218242 376816 218298 376825
rect 218242 376751 218298 376760
rect 218256 375193 218284 376751
rect 218242 375184 218298 375193
rect 218242 375119 218298 375128
rect 217324 374672 217376 374678
rect 217324 374614 217376 374620
rect 215944 373312 215996 373318
rect 215944 373254 215996 373260
rect 215392 355428 215444 355434
rect 215392 355370 215444 355376
rect 215298 350432 215354 350441
rect 215298 350367 215354 350376
rect 215312 350033 215340 350367
rect 215298 350024 215354 350033
rect 215298 349959 215354 349968
rect 215298 305824 215354 305833
rect 215298 305759 215354 305768
rect 215208 304292 215260 304298
rect 215208 304234 215260 304240
rect 215312 302258 215340 305759
rect 215300 302252 215352 302258
rect 215300 302194 215352 302200
rect 214746 299568 214802 299577
rect 214746 299503 214802 299512
rect 214562 296712 214618 296721
rect 214562 296647 214618 296656
rect 214576 295458 214604 296647
rect 214564 295452 214616 295458
rect 214564 295394 214616 295400
rect 213828 285728 213880 285734
rect 213828 285670 213880 285676
rect 213840 284172 213868 285670
rect 214760 284172 214788 299503
rect 215404 293865 215432 355370
rect 215852 302252 215904 302258
rect 215852 302194 215904 302200
rect 215390 293856 215446 293865
rect 215390 293791 215446 293800
rect 215404 292777 215432 293791
rect 215390 292768 215446 292777
rect 215390 292703 215446 292712
rect 215298 288416 215354 288425
rect 215298 288351 215354 288360
rect 215312 287609 215340 288351
rect 215298 287600 215354 287609
rect 215298 287535 215354 287544
rect 215206 287464 215262 287473
rect 215206 287399 215262 287408
rect 215220 285734 215248 287399
rect 215208 285728 215260 285734
rect 215208 285670 215260 285676
rect 215312 284172 215340 287535
rect 215864 284172 215892 302194
rect 215956 285705 215984 373254
rect 216034 350024 216090 350033
rect 216034 349959 216090 349968
rect 216048 330585 216076 349959
rect 216034 330576 216090 330585
rect 216034 330511 216090 330520
rect 216036 318164 216088 318170
rect 216036 318106 216088 318112
rect 216048 288425 216076 318106
rect 217336 296714 217364 374614
rect 219912 374066 219940 377604
rect 220832 377590 221582 377618
rect 222212 377590 223238 377618
rect 223592 377590 224894 377618
rect 226352 377590 226550 377618
rect 227732 377590 228206 377618
rect 229112 377590 229862 377618
rect 230492 377590 231518 377618
rect 231872 377590 233174 377618
rect 234632 377590 234830 377618
rect 236012 377590 236486 377618
rect 237392 377590 238142 377618
rect 219900 374060 219952 374066
rect 219900 374002 219952 374008
rect 220832 371385 220860 377590
rect 220818 371376 220874 371385
rect 220818 371311 220874 371320
rect 221462 371376 221518 371385
rect 221462 371311 221518 371320
rect 218702 370832 218758 370841
rect 218702 370767 218758 370776
rect 217244 296686 217364 296714
rect 216680 289876 216732 289882
rect 216680 289818 216732 289824
rect 216692 289134 216720 289818
rect 216680 289128 216732 289134
rect 216680 289070 216732 289076
rect 216680 288448 216732 288454
rect 216034 288416 216090 288425
rect 216680 288390 216732 288396
rect 216034 288351 216090 288360
rect 216692 287745 216720 288390
rect 216678 287736 216734 287745
rect 216678 287671 216734 287680
rect 217244 285841 217272 296686
rect 218058 289096 218114 289105
rect 218058 289031 218114 289040
rect 217322 287328 217378 287337
rect 217322 287263 217378 287272
rect 217230 285832 217286 285841
rect 217230 285767 217286 285776
rect 215942 285696 215998 285705
rect 215942 285631 215998 285640
rect 216772 284436 216824 284442
rect 216772 284378 216824 284384
rect 216784 284172 216812 284378
rect 217336 284172 217364 287263
rect 217690 287192 217746 287201
rect 217690 287127 217746 287136
rect 217704 284172 217732 287127
rect 218072 285802 218100 289031
rect 218716 287054 218744 370767
rect 221476 353977 221504 371311
rect 222212 354006 222240 377590
rect 222200 354000 222252 354006
rect 221462 353968 221518 353977
rect 222200 353942 222252 353948
rect 221462 353903 221518 353912
rect 223592 349042 223620 377590
rect 223580 349036 223632 349042
rect 223580 348978 223632 348984
rect 224224 349036 224276 349042
rect 224224 348978 224276 348984
rect 224236 347818 224264 348978
rect 224224 347812 224276 347818
rect 224224 347754 224276 347760
rect 222842 343768 222898 343777
rect 222842 343703 222898 343712
rect 220084 342304 220136 342310
rect 220084 342246 220136 342252
rect 219716 324352 219768 324358
rect 219716 324294 219768 324300
rect 218532 287026 218744 287054
rect 218060 285796 218112 285802
rect 218060 285738 218112 285744
rect 218532 284481 218560 287026
rect 218612 286680 218664 286686
rect 218612 286622 218664 286628
rect 218518 284472 218574 284481
rect 218518 284407 218574 284416
rect 218532 284186 218560 284407
rect 218270 284158 218560 284186
rect 218624 284172 218652 286622
rect 219164 285728 219216 285734
rect 219164 285670 219216 285676
rect 219176 284172 219204 285670
rect 219728 284172 219756 324294
rect 220096 291009 220124 342246
rect 220176 329112 220228 329118
rect 220176 329054 220228 329060
rect 220188 324358 220216 329054
rect 220176 324352 220228 324358
rect 220176 324294 220228 324300
rect 220176 322312 220228 322318
rect 220176 322254 220228 322260
rect 220188 307057 220216 322254
rect 221462 320920 221518 320929
rect 221462 320855 221518 320864
rect 220174 307048 220230 307057
rect 220174 306983 220230 306992
rect 220176 304360 220228 304366
rect 220176 304302 220228 304308
rect 220188 295497 220216 304302
rect 221476 296714 221504 320855
rect 222476 314696 222528 314702
rect 222476 314638 222528 314644
rect 221556 301504 221608 301510
rect 221556 301446 221608 301452
rect 221200 296686 221504 296714
rect 220174 295488 220230 295497
rect 220174 295423 220230 295432
rect 220818 295488 220874 295497
rect 220818 295423 220874 295432
rect 220176 292596 220228 292602
rect 220176 292538 220228 292544
rect 220082 291000 220138 291009
rect 220082 290935 220138 290944
rect 220096 286686 220124 290935
rect 220188 288561 220216 292538
rect 220174 288552 220230 288561
rect 220174 288487 220230 288496
rect 220084 286680 220136 286686
rect 220084 286622 220136 286628
rect 220188 284186 220216 288487
rect 220832 285326 220860 295423
rect 221200 292777 221228 296686
rect 221186 292768 221242 292777
rect 221186 292703 221242 292712
rect 220820 285320 220872 285326
rect 220820 285262 220872 285268
rect 220188 284158 220662 284186
rect 221200 284172 221228 292703
rect 221568 292602 221596 301446
rect 221556 292596 221608 292602
rect 221556 292538 221608 292544
rect 222108 292596 222160 292602
rect 222108 292538 222160 292544
rect 221280 285320 221332 285326
rect 221280 285262 221332 285268
rect 221292 284186 221320 285262
rect 221292 284158 221582 284186
rect 222120 284172 222148 292538
rect 222488 284172 222516 314638
rect 222856 285841 222884 343703
rect 224236 340202 224264 347754
rect 224224 340196 224276 340202
rect 224224 340138 224276 340144
rect 224224 336796 224276 336802
rect 224224 336738 224276 336744
rect 223028 315308 223080 315314
rect 223028 315250 223080 315256
rect 223040 314702 223068 315250
rect 223028 314696 223080 314702
rect 223028 314638 223080 314644
rect 223488 313948 223540 313954
rect 223488 313890 223540 313896
rect 223500 309806 223528 313890
rect 223488 309800 223540 309806
rect 223488 309742 223540 309748
rect 223026 298752 223082 298761
rect 223026 298687 223082 298696
rect 223040 289921 223068 298687
rect 223026 289912 223082 289921
rect 223026 289847 223082 289856
rect 222842 285832 222898 285841
rect 222842 285767 222898 285776
rect 223040 284172 223068 289847
rect 223580 287088 223632 287094
rect 223580 287030 223632 287036
rect 205362 283928 205418 283937
rect 205192 283900 205362 283914
rect 205206 283886 205362 283900
rect 200132 283529 200160 283886
rect 214470 283928 214526 283937
rect 214406 283886 214470 283914
rect 205362 283863 205418 283872
rect 214470 283863 214526 283872
rect 216126 283928 216182 283937
rect 220266 283928 220322 283937
rect 216182 283886 216246 283914
rect 220110 283886 220266 283914
rect 216126 283863 216182 283872
rect 223592 283914 223620 287030
rect 224236 286414 224264 336738
rect 225604 330540 225656 330546
rect 225604 330482 225656 330488
rect 224316 295452 224368 295458
rect 224316 295394 224368 295400
rect 224224 286408 224276 286414
rect 224224 286350 224276 286356
rect 224328 285734 224356 295394
rect 224868 289128 224920 289134
rect 224868 289070 224920 289076
rect 224880 288454 224908 289070
rect 224868 288448 224920 288454
rect 225616 288425 225644 330482
rect 225694 315344 225750 315353
rect 225694 315279 225750 315288
rect 225708 294137 225736 315279
rect 226352 297537 226380 377590
rect 226984 356108 227036 356114
rect 226984 356050 227036 356056
rect 226996 329118 227024 356050
rect 227732 351393 227760 377590
rect 229112 362545 229140 377590
rect 230492 365809 230520 377590
rect 230478 365800 230534 365809
rect 230478 365735 230534 365744
rect 231122 365800 231178 365809
rect 231122 365735 231178 365744
rect 229098 362536 229154 362545
rect 229098 362471 229154 362480
rect 227718 351384 227774 351393
rect 227718 351319 227774 351328
rect 229744 339516 229796 339522
rect 229744 339458 229796 339464
rect 228364 333260 228416 333266
rect 228364 333202 228416 333208
rect 226984 329112 227036 329118
rect 226984 329054 227036 329060
rect 226982 319424 227038 319433
rect 226982 319359 227038 319368
rect 226338 297528 226394 297537
rect 226338 297463 226394 297472
rect 226706 296984 226762 296993
rect 226706 296919 226762 296928
rect 225694 294128 225750 294137
rect 225694 294063 225750 294072
rect 226720 291145 226748 296919
rect 226890 294128 226946 294137
rect 226890 294063 226946 294072
rect 226706 291136 226762 291145
rect 226706 291071 226762 291080
rect 224868 288390 224920 288396
rect 225602 288416 225658 288425
rect 224316 285728 224368 285734
rect 223946 285696 224002 285705
rect 224316 285670 224368 285676
rect 223946 285631 224002 285640
rect 223960 284172 223988 285631
rect 224880 284186 224908 288390
rect 225602 288351 225658 288360
rect 225052 286408 225104 286414
rect 225052 286350 225104 286356
rect 225064 285705 225092 286350
rect 225050 285696 225106 285705
rect 225050 285631 225106 285640
rect 224526 284158 224908 284186
rect 225064 284172 225092 285631
rect 225616 284186 225644 288351
rect 225970 285832 226026 285841
rect 225970 285767 226026 285776
rect 225446 284158 225644 284186
rect 225984 284172 226012 285767
rect 226524 285728 226576 285734
rect 226524 285670 226576 285676
rect 226536 284172 226564 285670
rect 226904 284172 226932 294063
rect 226996 291281 227024 319359
rect 227442 316704 227498 316713
rect 227442 316639 227498 316648
rect 227456 316169 227484 316639
rect 227442 316160 227498 316169
rect 227442 316095 227498 316104
rect 226982 291272 227038 291281
rect 226982 291207 227038 291216
rect 227456 284172 227484 316095
rect 227812 311908 227864 311914
rect 227812 311850 227864 311856
rect 227626 291272 227682 291281
rect 227626 291207 227682 291216
rect 227640 285802 227668 291207
rect 227628 285796 227680 285802
rect 227628 285738 227680 285744
rect 227824 284172 227852 311850
rect 227902 292496 227958 292505
rect 227902 292431 227958 292440
rect 227916 292097 227944 292431
rect 227902 292088 227958 292097
rect 227902 292023 227958 292032
rect 227916 284186 227944 292023
rect 228376 285734 228404 333202
rect 228548 320884 228600 320890
rect 228548 320826 228600 320832
rect 228456 317484 228508 317490
rect 228456 317426 228508 317432
rect 228468 292097 228496 317426
rect 228560 311914 228588 320826
rect 228548 311908 228600 311914
rect 228548 311850 228600 311856
rect 228454 292088 228510 292097
rect 228454 292023 228510 292032
rect 229756 289882 229784 339458
rect 231136 306513 231164 365735
rect 231872 361622 231900 377590
rect 233884 374740 233936 374746
rect 233884 374682 233936 374688
rect 233146 362400 233202 362409
rect 233146 362335 233202 362344
rect 233160 361729 233188 362335
rect 232502 361720 232558 361729
rect 232502 361655 232558 361664
rect 233146 361720 233202 361729
rect 233146 361655 233202 361664
rect 231860 361616 231912 361622
rect 231860 361558 231912 361564
rect 232226 320648 232282 320657
rect 232226 320583 232282 320592
rect 231122 306504 231178 306513
rect 231122 306439 231178 306448
rect 230294 301744 230350 301753
rect 230294 301679 230350 301688
rect 230308 296714 230336 301679
rect 230388 298852 230440 298858
rect 230388 298794 230440 298800
rect 230400 297401 230428 298794
rect 231136 297537 231164 306439
rect 231676 303680 231728 303686
rect 231676 303622 231728 303628
rect 231122 297528 231178 297537
rect 231122 297463 231178 297472
rect 230386 297392 230442 297401
rect 230386 297327 230442 297336
rect 231124 296744 231176 296750
rect 230308 296686 230428 296714
rect 231124 296686 231176 296692
rect 229744 289876 229796 289882
rect 229744 289818 229796 289824
rect 228916 285796 228968 285802
rect 228916 285738 228968 285744
rect 228364 285728 228416 285734
rect 228364 285670 228416 285676
rect 227916 284158 228390 284186
rect 228928 284172 228956 285738
rect 229284 285728 229336 285734
rect 229284 285670 229336 285676
rect 223762 283928 223818 283937
rect 223592 283900 223762 283914
rect 223606 283886 223762 283900
rect 220266 283863 220322 283872
rect 229296 283914 229324 285670
rect 229756 284186 229784 289818
rect 229756 284158 229862 284186
rect 230400 284172 230428 296686
rect 231136 288386 231164 296686
rect 231124 288380 231176 288386
rect 231124 288322 231176 288328
rect 231136 284186 231164 288322
rect 231136 284158 231334 284186
rect 231688 284172 231716 303622
rect 232240 284172 232268 320583
rect 232516 289105 232544 361655
rect 232596 361616 232648 361622
rect 232596 361558 232648 361564
rect 232608 315314 232636 361558
rect 233896 353258 233924 374682
rect 234632 366858 234660 377590
rect 234620 366852 234672 366858
rect 234620 366794 234672 366800
rect 235356 366852 235408 366858
rect 235356 366794 235408 366800
rect 235368 365770 235396 366794
rect 235356 365764 235408 365770
rect 235356 365706 235408 365712
rect 235264 363656 235316 363662
rect 235264 363598 235316 363604
rect 234528 359576 234580 359582
rect 234528 359518 234580 359524
rect 234540 357406 234568 359518
rect 234528 357400 234580 357406
rect 234528 357342 234580 357348
rect 233884 353252 233936 353258
rect 233884 353194 233936 353200
rect 232686 328672 232742 328681
rect 232686 328607 232742 328616
rect 232700 320657 232728 328607
rect 233896 323785 233924 353194
rect 234436 324964 234488 324970
rect 234436 324906 234488 324912
rect 233882 323776 233938 323785
rect 233882 323711 233938 323720
rect 232686 320648 232742 320657
rect 232686 320583 232742 320592
rect 232700 320249 232728 320583
rect 232686 320240 232742 320249
rect 232686 320175 232742 320184
rect 232688 315376 232740 315382
rect 232688 315318 232740 315324
rect 232596 315308 232648 315314
rect 232596 315250 232648 315256
rect 232502 289096 232558 289105
rect 232502 289031 232558 289040
rect 232700 287026 232728 315318
rect 232778 292632 232834 292641
rect 234448 292602 234476 324906
rect 234540 304366 234568 357342
rect 234618 314800 234674 314809
rect 234618 314735 234674 314744
rect 234528 304360 234580 304366
rect 234528 304302 234580 304308
rect 234540 303686 234568 304302
rect 234528 303680 234580 303686
rect 234528 303622 234580 303628
rect 234526 298208 234582 298217
rect 234526 298143 234582 298152
rect 232778 292567 232834 292576
rect 234436 292596 234488 292602
rect 232792 288561 232820 292567
rect 234436 292538 234488 292544
rect 233698 290456 233754 290465
rect 233698 290391 233754 290400
rect 232778 288552 232834 288561
rect 232778 288487 232834 288496
rect 232688 287020 232740 287026
rect 232688 286962 232740 286968
rect 232792 284172 232820 288487
rect 233148 287156 233200 287162
rect 233148 287098 233200 287104
rect 233160 284172 233188 287098
rect 233712 284172 233740 290391
rect 234250 287192 234306 287201
rect 234250 287127 234306 287136
rect 234264 287026 234292 287127
rect 234252 287020 234304 287026
rect 234252 286962 234304 286968
rect 234264 284172 234292 286962
rect 234448 285734 234476 292538
rect 234540 291009 234568 298143
rect 234526 291000 234582 291009
rect 234526 290935 234582 290944
rect 234436 285728 234488 285734
rect 234436 285670 234488 285676
rect 234632 284172 234660 314735
rect 235276 295322 235304 363598
rect 235368 348498 235396 365706
rect 235356 348492 235408 348498
rect 235356 348434 235408 348440
rect 235354 345944 235410 345953
rect 235354 345879 235410 345888
rect 235368 314809 235396 345879
rect 236012 322153 236040 377590
rect 237392 344457 237420 377590
rect 239784 374678 239812 377604
rect 240152 377590 241454 377618
rect 239772 374672 239824 374678
rect 239772 374614 239824 374620
rect 238022 364440 238078 364449
rect 238022 364375 238078 364384
rect 237378 344448 237434 344457
rect 237378 344383 237434 344392
rect 237932 339448 237984 339454
rect 237932 339390 237984 339396
rect 237944 338230 237972 339390
rect 237932 338224 237984 338230
rect 237932 338166 237984 338172
rect 236736 327140 236788 327146
rect 236736 327082 236788 327088
rect 235998 322144 236054 322153
rect 235998 322079 236054 322088
rect 235354 314800 235410 314809
rect 235354 314735 235410 314744
rect 235356 312588 235408 312594
rect 235356 312530 235408 312536
rect 235264 295316 235316 295322
rect 235264 295258 235316 295264
rect 235172 285728 235224 285734
rect 235172 285670 235224 285676
rect 235184 284172 235212 285670
rect 235276 284186 235304 295258
rect 235368 287706 235396 312530
rect 236642 308544 236698 308553
rect 236642 308479 236698 308488
rect 236000 305040 236052 305046
rect 236000 304982 236052 304988
rect 236092 305040 236144 305046
rect 236092 304982 236144 304988
rect 235356 287700 235408 287706
rect 235356 287642 235408 287648
rect 236012 285705 236040 304982
rect 235998 285696 236054 285705
rect 235998 285631 236054 285640
rect 235276 284158 235566 284186
rect 236104 284172 236132 304982
rect 236656 285841 236684 308479
rect 236748 305046 236776 327082
rect 238036 322318 238064 364375
rect 240152 339454 240180 377590
rect 241426 375320 241482 375329
rect 241426 375255 241482 375264
rect 241440 374105 241468 375255
rect 243096 374746 243124 377604
rect 244752 374814 244780 377604
rect 245672 377590 246422 377618
rect 244740 374808 244792 374814
rect 244740 374750 244792 374756
rect 242164 374740 242216 374746
rect 242164 374682 242216 374688
rect 243084 374740 243136 374746
rect 243084 374682 243136 374688
rect 241426 374096 241482 374105
rect 241426 374031 241482 374040
rect 241440 369170 241468 374031
rect 241428 369164 241480 369170
rect 241428 369106 241480 369112
rect 242176 356697 242204 374682
rect 245672 370705 245700 377590
rect 248064 376038 248092 377604
rect 248432 377590 249734 377618
rect 248052 376032 248104 376038
rect 248052 375974 248104 375980
rect 248064 374105 248092 375974
rect 248050 374096 248106 374105
rect 248050 374031 248106 374040
rect 245658 370696 245714 370705
rect 245658 370631 245714 370640
rect 246302 360224 246358 360233
rect 246302 360159 246358 360168
rect 244922 357640 244978 357649
rect 244922 357575 244978 357584
rect 242162 356688 242218 356697
rect 242162 356623 242218 356632
rect 242164 348424 242216 348430
rect 242164 348366 242216 348372
rect 240140 339448 240192 339454
rect 240140 339390 240192 339396
rect 238668 338224 238720 338230
rect 238668 338166 238720 338172
rect 238114 325000 238170 325009
rect 238114 324935 238170 324944
rect 238024 322312 238076 322318
rect 238024 322254 238076 322260
rect 238128 311846 238156 324935
rect 238576 313404 238628 313410
rect 238576 313346 238628 313352
rect 238116 311840 238168 311846
rect 238116 311782 238168 311788
rect 238024 311228 238076 311234
rect 238024 311170 238076 311176
rect 236736 305040 236788 305046
rect 236736 304982 236788 304988
rect 238036 301510 238064 311170
rect 238024 301504 238076 301510
rect 238024 301446 238076 301452
rect 238114 286104 238170 286113
rect 238114 286039 238170 286048
rect 237286 285968 237342 285977
rect 237654 285968 237710 285977
rect 237342 285926 237512 285954
rect 237286 285903 237342 285912
rect 236642 285832 236698 285841
rect 236642 285767 236698 285776
rect 237380 285796 237432 285802
rect 236656 284172 236684 285767
rect 237380 285738 237432 285744
rect 237392 285025 237420 285738
rect 237378 285016 237434 285025
rect 237484 284986 237512 285926
rect 237654 285903 237710 285912
rect 237564 285728 237616 285734
rect 237564 285670 237616 285676
rect 237378 284951 237434 284960
rect 237472 284980 237524 284986
rect 237472 284922 237524 284928
rect 237576 284172 237604 285670
rect 237668 285569 237696 285903
rect 237654 285560 237710 285569
rect 237654 285495 237710 285504
rect 238128 284172 238156 286039
rect 238484 285796 238536 285802
rect 238484 285738 238536 285744
rect 238496 284172 238524 285738
rect 238588 285734 238616 313346
rect 238680 310486 238708 338166
rect 240048 327140 240100 327146
rect 240048 327082 240100 327088
rect 239404 311840 239456 311846
rect 239404 311782 239456 311788
rect 239416 311234 239444 311782
rect 239404 311228 239456 311234
rect 239404 311170 239456 311176
rect 239588 311228 239640 311234
rect 239588 311170 239640 311176
rect 238668 310480 238720 310486
rect 238668 310422 238720 310428
rect 239034 309768 239090 309777
rect 239034 309703 239090 309712
rect 239048 307834 239076 309703
rect 239036 307828 239088 307834
rect 239036 307770 239088 307776
rect 238576 285728 238628 285734
rect 238576 285670 238628 285676
rect 239048 284172 239076 307770
rect 239600 284172 239628 311170
rect 240060 284186 240088 327082
rect 240876 320952 240928 320958
rect 240876 320894 240928 320900
rect 240888 320210 240916 320894
rect 240876 320204 240928 320210
rect 240876 320146 240928 320152
rect 240140 316124 240192 316130
rect 240140 316066 240192 316072
rect 240152 313954 240180 316066
rect 240140 313948 240192 313954
rect 240140 313890 240192 313896
rect 240232 310480 240284 310486
rect 240232 310422 240284 310428
rect 240244 290465 240272 310422
rect 240230 290456 240286 290465
rect 240230 290391 240286 290400
rect 240508 289128 240560 289134
rect 240508 289070 240560 289076
rect 239982 284158 240088 284186
rect 240520 284172 240548 289070
rect 240888 284172 240916 320146
rect 241980 313336 242032 313342
rect 241980 313278 242032 313284
rect 241426 288688 241482 288697
rect 241426 288623 241482 288632
rect 241440 284172 241468 288623
rect 241992 284172 242020 313278
rect 242176 306374 242204 348366
rect 243544 340196 243596 340202
rect 243544 340138 243596 340144
rect 242254 330440 242310 330449
rect 242254 330375 242310 330384
rect 242268 313342 242296 330375
rect 242256 313336 242308 313342
rect 242256 313278 242308 313284
rect 242176 306346 242388 306374
rect 242360 285734 242388 306346
rect 243452 298852 243504 298858
rect 243452 298794 243504 298800
rect 243082 287192 243138 287201
rect 243082 287127 243138 287136
rect 243096 287054 243124 287127
rect 243004 287026 243124 287054
rect 242348 285728 242400 285734
rect 242348 285670 242400 285676
rect 242898 285696 242954 285705
rect 242360 284172 242388 285670
rect 242898 285631 242954 285640
rect 242912 284172 242940 285631
rect 243004 284073 243032 287026
rect 243082 286104 243138 286113
rect 243082 286039 243138 286048
rect 243096 284209 243124 286039
rect 243082 284200 243138 284209
rect 243464 284172 243492 298794
rect 243556 285705 243584 340138
rect 244278 328400 244334 328409
rect 244278 328335 244334 328344
rect 244292 327729 244320 328335
rect 244278 327720 244334 327729
rect 244278 327655 244334 327664
rect 244292 315081 244320 327655
rect 244372 315308 244424 315314
rect 244372 315250 244424 315256
rect 244278 315072 244334 315081
rect 244278 315007 244334 315016
rect 244278 313984 244334 313993
rect 244278 313919 244334 313928
rect 244004 306468 244056 306474
rect 244004 306410 244056 306416
rect 243542 285696 243598 285705
rect 243542 285631 243598 285640
rect 243912 284980 243964 284986
rect 243912 284922 243964 284928
rect 243818 284880 243874 284889
rect 243818 284815 243874 284824
rect 243832 284345 243860 284815
rect 243818 284336 243874 284345
rect 243818 284271 243874 284280
rect 243832 284172 243860 284271
rect 243082 284135 243138 284144
rect 242990 284064 243046 284073
rect 242990 283999 243046 284008
rect 229466 283928 229522 283937
rect 229296 283900 229466 283914
rect 229310 283886 229466 283900
rect 223762 283863 223818 283872
rect 230938 283928 230994 283937
rect 230782 283886 230938 283914
rect 229466 283863 229522 283872
rect 230938 283863 230994 283872
rect 236734 283928 236790 283937
rect 236790 283886 237038 283914
rect 236734 283863 236790 283872
rect 200118 283520 200174 283529
rect 200118 283455 200174 283464
rect 199568 271176 199620 271182
rect 199568 271118 199620 271124
rect 243924 267734 243952 284922
rect 244016 279993 244044 306410
rect 244002 279984 244058 279993
rect 244002 279919 244058 279928
rect 244292 269657 244320 313919
rect 244384 278089 244412 315250
rect 244936 311137 244964 357575
rect 245014 356688 245070 356697
rect 245014 356623 245070 356632
rect 245028 344457 245056 356623
rect 245014 344448 245070 344457
rect 245014 344383 245070 344392
rect 245016 337408 245068 337414
rect 245016 337350 245068 337356
rect 245028 328409 245056 337350
rect 245658 334792 245714 334801
rect 245658 334727 245714 334736
rect 245014 328400 245070 328409
rect 245014 328335 245070 328344
rect 244922 311128 244978 311137
rect 244922 311063 244978 311072
rect 244464 300144 244516 300150
rect 244464 300086 244516 300092
rect 244370 278080 244426 278089
rect 244370 278015 244426 278024
rect 244384 277438 244412 278015
rect 244372 277432 244424 277438
rect 244372 277374 244424 277380
rect 244278 269648 244334 269657
rect 244278 269583 244334 269592
rect 244476 268841 244504 300086
rect 245672 298858 245700 334727
rect 246316 325009 246344 360159
rect 247038 334656 247094 334665
rect 247038 334591 247094 334600
rect 246302 325000 246358 325009
rect 246302 324935 246358 324944
rect 246304 322244 246356 322250
rect 246304 322186 246356 322192
rect 245752 300212 245804 300218
rect 245752 300154 245804 300160
rect 245660 298852 245712 298858
rect 245660 298794 245712 298800
rect 245658 294536 245714 294545
rect 245658 294471 245714 294480
rect 245016 285796 245068 285802
rect 245016 285738 245068 285744
rect 244922 273456 244978 273465
rect 244922 273391 244978 273400
rect 244462 268832 244518 268841
rect 244462 268767 244518 268776
rect 244476 267782 244504 268767
rect 244464 267776 244516 267782
rect 243924 267706 244044 267734
rect 244464 267718 244516 267724
rect 244016 259321 244044 267706
rect 244462 264480 244518 264489
rect 244462 264415 244518 264424
rect 244370 261760 244426 261769
rect 244370 261695 244426 261704
rect 244002 259312 244058 259321
rect 244002 259247 244058 259256
rect 199474 250472 199530 250481
rect 199474 250407 199530 250416
rect 200026 249520 200082 249529
rect 200026 249455 200082 249464
rect 199476 246356 199528 246362
rect 199476 246298 199528 246304
rect 199384 238060 199436 238066
rect 199384 238002 199436 238008
rect 199396 237726 199424 238002
rect 199384 237720 199436 237726
rect 199384 237662 199436 237668
rect 198738 237416 198794 237425
rect 198738 237351 198794 237360
rect 198556 231124 198608 231130
rect 198556 231066 198608 231072
rect 198462 229800 198518 229809
rect 198462 229735 198518 229744
rect 198752 216714 198780 237351
rect 199488 235890 199516 246298
rect 199934 242312 199990 242321
rect 199934 242247 199990 242256
rect 199568 242208 199620 242214
rect 199568 242150 199620 242156
rect 199580 237386 199608 242150
rect 199842 240272 199898 240281
rect 199842 240207 199898 240216
rect 199856 240038 199884 240207
rect 199948 240145 199976 242247
rect 199934 240136 199990 240145
rect 199934 240071 199990 240080
rect 199844 240032 199896 240038
rect 199844 239974 199896 239980
rect 199568 237380 199620 237386
rect 199568 237322 199620 237328
rect 199476 235884 199528 235890
rect 199476 235826 199528 235832
rect 199384 234932 199436 234938
rect 199384 234874 199436 234880
rect 199396 228857 199424 234874
rect 199382 228848 199438 228857
rect 199382 228783 199438 228792
rect 198740 216708 198792 216714
rect 198740 216650 198792 216656
rect 198370 195392 198426 195401
rect 198370 195327 198426 195336
rect 198096 193860 198148 193866
rect 198096 193802 198148 193808
rect 200040 192438 200068 249455
rect 244002 244216 244058 244225
rect 244002 244151 244058 244160
rect 200118 240544 200174 240553
rect 200118 240479 200174 240488
rect 200132 240242 200160 240479
rect 200120 240236 200172 240242
rect 200120 240178 200172 240184
rect 200118 240136 200174 240145
rect 200118 240071 200174 240080
rect 200132 237289 200160 240071
rect 200224 238066 200252 240244
rect 200592 239737 200620 240244
rect 201144 240106 201172 240244
rect 201132 240100 201184 240106
rect 201132 240042 201184 240048
rect 201040 240032 201092 240038
rect 201040 239974 201092 239980
rect 200578 239728 200634 239737
rect 200578 239663 200634 239672
rect 200592 238754 200620 239663
rect 200592 238726 200804 238754
rect 200212 238060 200264 238066
rect 200212 238002 200264 238008
rect 200118 237280 200174 237289
rect 200118 237215 200174 237224
rect 200776 224262 200804 238726
rect 201052 229094 201080 239974
rect 201144 235618 201172 240042
rect 201512 238754 201540 240244
rect 201512 238726 201632 238754
rect 201604 238377 201632 238726
rect 201590 238368 201646 238377
rect 201590 238303 201646 238312
rect 201314 237144 201370 237153
rect 201314 237079 201370 237088
rect 201328 235793 201356 237079
rect 201314 235784 201370 235793
rect 201314 235719 201370 235728
rect 201132 235612 201184 235618
rect 201132 235554 201184 235560
rect 201314 235240 201370 235249
rect 201314 235175 201370 235184
rect 201328 234530 201356 235175
rect 201316 234524 201368 234530
rect 201316 234466 201368 234472
rect 201052 229066 201172 229094
rect 200764 224256 200816 224262
rect 200764 224198 200816 224204
rect 200028 192432 200080 192438
rect 200028 192374 200080 192380
rect 198002 186280 198058 186289
rect 198002 186215 198058 186224
rect 197266 115152 197322 115161
rect 197266 115087 197322 115096
rect 198016 100065 198044 186215
rect 200764 183592 200816 183598
rect 200764 183534 200816 183540
rect 198096 179512 198148 179518
rect 198096 179454 198148 179460
rect 198108 166938 198136 179454
rect 200776 168298 200804 183534
rect 200764 168292 200816 168298
rect 200764 168234 200816 168240
rect 198096 166932 198148 166938
rect 198096 166874 198148 166880
rect 198096 150544 198148 150550
rect 198096 150486 198148 150492
rect 198108 129062 198136 150486
rect 198188 140888 198240 140894
rect 198188 140830 198240 140836
rect 198096 129056 198148 129062
rect 198096 128998 198148 129004
rect 198096 117428 198148 117434
rect 198096 117370 198148 117376
rect 198002 100056 198058 100065
rect 196808 100020 196860 100026
rect 198002 99991 198058 100000
rect 196808 99962 196860 99968
rect 196808 96688 196860 96694
rect 196808 96630 196860 96636
rect 196716 88324 196768 88330
rect 196716 88266 196768 88272
rect 196820 69018 196848 96630
rect 198002 82240 198058 82249
rect 198002 82175 198058 82184
rect 196808 69012 196860 69018
rect 196808 68954 196860 68960
rect 198016 15910 198044 82175
rect 198108 55214 198136 117370
rect 198200 110537 198228 140830
rect 200764 138712 200816 138718
rect 200764 138654 200816 138660
rect 199476 134632 199528 134638
rect 199476 134574 199528 134580
rect 199382 113384 199438 113393
rect 199382 113319 199438 113328
rect 198186 110528 198242 110537
rect 198186 110463 198242 110472
rect 198188 102196 198240 102202
rect 198188 102138 198240 102144
rect 198200 74497 198228 102138
rect 198186 74488 198242 74497
rect 198186 74423 198242 74432
rect 199396 67590 199424 113319
rect 199488 87553 199516 134574
rect 199474 87544 199530 87553
rect 199474 87479 199530 87488
rect 199384 67584 199436 67590
rect 199384 67526 199436 67532
rect 198096 55208 198148 55214
rect 198096 55150 198148 55156
rect 200776 25634 200804 138654
rect 201144 93809 201172 229066
rect 201604 219434 201632 238303
rect 202064 234433 202092 240244
rect 202616 238754 202644 240244
rect 202880 240168 202932 240174
rect 202880 240110 202932 240116
rect 202156 238726 202644 238754
rect 202156 238513 202184 238726
rect 202142 238504 202198 238513
rect 202142 238439 202198 238448
rect 202050 234424 202106 234433
rect 202050 234359 202106 234368
rect 201512 219406 201632 219434
rect 201512 218006 201540 219406
rect 201500 218000 201552 218006
rect 201500 217942 201552 217948
rect 202052 218000 202104 218006
rect 202052 217942 202104 217948
rect 202064 217394 202092 217942
rect 202052 217388 202104 217394
rect 202052 217330 202104 217336
rect 202156 192574 202184 238439
rect 202510 234424 202566 234433
rect 202510 234359 202566 234368
rect 202524 227089 202552 234359
rect 202326 227080 202382 227089
rect 202326 227015 202382 227024
rect 202510 227080 202566 227089
rect 202510 227015 202566 227024
rect 202236 224256 202288 224262
rect 202236 224198 202288 224204
rect 202144 192568 202196 192574
rect 202144 192510 202196 192516
rect 201500 192432 201552 192438
rect 201500 192374 201552 192380
rect 201512 188358 201540 192374
rect 201500 188352 201552 188358
rect 201500 188294 201552 188300
rect 202144 187740 202196 187746
rect 202144 187682 202196 187688
rect 202156 169658 202184 187682
rect 202248 185609 202276 224198
rect 202340 218006 202368 227015
rect 202328 218000 202380 218006
rect 202328 217942 202380 217948
rect 202234 185600 202290 185609
rect 202234 185535 202290 185544
rect 202144 169652 202196 169658
rect 202144 169594 202196 169600
rect 202236 151836 202288 151842
rect 202236 151778 202288 151784
rect 202144 133952 202196 133958
rect 202144 133894 202196 133900
rect 202156 113898 202184 133894
rect 202144 113892 202196 113898
rect 202144 113834 202196 113840
rect 202142 112432 202198 112441
rect 202142 112367 202198 112376
rect 201130 93800 201186 93809
rect 201130 93735 201186 93744
rect 202156 30297 202184 112367
rect 202248 97306 202276 151778
rect 202420 125656 202472 125662
rect 202420 125598 202472 125604
rect 202328 104984 202380 104990
rect 202328 104926 202380 104932
rect 202236 97300 202288 97306
rect 202236 97242 202288 97248
rect 202234 89040 202290 89049
rect 202234 88975 202290 88984
rect 202142 30288 202198 30297
rect 202142 30223 202198 30232
rect 200764 25628 200816 25634
rect 200764 25570 200816 25576
rect 198004 15904 198056 15910
rect 198004 15846 198056 15852
rect 196624 13796 196676 13802
rect 196624 13738 196676 13744
rect 195244 10396 195296 10402
rect 195244 10338 195296 10344
rect 202248 9042 202276 88975
rect 202340 71738 202368 104926
rect 202432 94518 202460 125598
rect 202604 111920 202656 111926
rect 202604 111862 202656 111868
rect 202616 105602 202644 111862
rect 202604 105596 202656 105602
rect 202604 105538 202656 105544
rect 202892 100026 202920 240110
rect 202984 237386 203012 240244
rect 203432 240168 203484 240174
rect 203536 240122 203564 240244
rect 203484 240116 203564 240122
rect 203432 240110 203564 240116
rect 203444 240094 203564 240110
rect 202972 237380 203024 237386
rect 202972 237322 203024 237328
rect 202984 236026 203012 237322
rect 204088 236026 204116 240244
rect 202972 236020 203024 236026
rect 202972 235962 203024 235968
rect 203524 236020 203576 236026
rect 203524 235962 203576 235968
rect 204076 236020 204128 236026
rect 204076 235962 204128 235968
rect 203536 208078 203564 235962
rect 204088 235929 204116 235962
rect 204074 235920 204130 235929
rect 204074 235855 204130 235864
rect 204456 228857 204484 240244
rect 205008 230382 205036 240244
rect 205376 237289 205404 240244
rect 205928 238754 205956 240244
rect 206008 239488 206060 239494
rect 206008 239430 206060 239436
rect 205836 238726 205956 238754
rect 205836 238649 205864 238726
rect 206020 238678 206048 239430
rect 206008 238672 206060 238678
rect 205822 238640 205878 238649
rect 206008 238614 206060 238620
rect 205822 238575 205878 238584
rect 205362 237280 205418 237289
rect 205362 237215 205418 237224
rect 204996 230376 205048 230382
rect 204996 230318 205048 230324
rect 205376 229094 205404 237215
rect 204916 229066 205404 229094
rect 204442 228848 204498 228857
rect 204442 228783 204498 228792
rect 204456 227769 204484 228783
rect 204442 227760 204498 227769
rect 204442 227695 204498 227704
rect 203524 208072 203576 208078
rect 203524 208014 203576 208020
rect 204536 188420 204588 188426
rect 204536 188362 204588 188368
rect 204548 186318 204576 188362
rect 204536 186312 204588 186318
rect 204536 186254 204588 186260
rect 203614 127256 203670 127265
rect 203614 127191 203670 127200
rect 203522 123584 203578 123593
rect 203522 123519 203578 123528
rect 202880 100020 202932 100026
rect 202880 99962 202932 99968
rect 202420 94512 202472 94518
rect 202420 94454 202472 94460
rect 202328 71732 202380 71738
rect 202328 71674 202380 71680
rect 203536 62082 203564 123519
rect 203628 95849 203656 127191
rect 203708 107772 203760 107778
rect 203708 107714 203760 107720
rect 203614 95840 203670 95849
rect 203614 95775 203670 95784
rect 203720 81433 203748 107714
rect 204916 95849 204944 229066
rect 204994 227760 205050 227769
rect 204994 227695 205050 227704
rect 205008 211857 205036 227695
rect 204994 211848 205050 211857
rect 204994 211783 205050 211792
rect 205836 205630 205864 238575
rect 206376 235612 206428 235618
rect 206376 235554 206428 235560
rect 205824 205624 205876 205630
rect 205824 205566 205876 205572
rect 205836 205154 205864 205566
rect 205824 205148 205876 205154
rect 205824 205090 205876 205096
rect 206284 198076 206336 198082
rect 206284 198018 206336 198024
rect 204996 185700 205048 185706
rect 204996 185642 205048 185648
rect 205008 180810 205036 185642
rect 204996 180804 205048 180810
rect 204996 180746 205048 180752
rect 204996 146940 205048 146946
rect 204996 146882 205048 146888
rect 204902 95840 204958 95849
rect 204902 95775 204958 95784
rect 204904 87644 204956 87650
rect 204904 87586 204956 87592
rect 203706 81424 203762 81433
rect 203706 81359 203762 81368
rect 203524 62076 203576 62082
rect 203524 62018 203576 62024
rect 204916 29714 204944 87586
rect 205008 84833 205036 146882
rect 205088 124908 205140 124914
rect 205088 124850 205140 124856
rect 204994 84824 205050 84833
rect 204994 84759 205050 84768
rect 205100 64870 205128 124850
rect 205180 98116 205232 98122
rect 205180 98058 205232 98064
rect 205088 64864 205140 64870
rect 205088 64806 205140 64812
rect 205192 49706 205220 98058
rect 206296 86329 206324 198018
rect 206388 188426 206416 235554
rect 206480 212498 206508 240244
rect 206848 233170 206876 240244
rect 207112 237448 207164 237454
rect 207112 237390 207164 237396
rect 206836 233164 206888 233170
rect 206836 233106 206888 233112
rect 206848 229158 206876 233106
rect 206836 229152 206888 229158
rect 206836 229094 206888 229100
rect 207124 216481 207152 237390
rect 207110 216472 207166 216481
rect 207110 216407 207166 216416
rect 207124 215393 207152 216407
rect 207110 215384 207166 215393
rect 207110 215319 207166 215328
rect 206468 212492 206520 212498
rect 206468 212434 206520 212440
rect 206480 195294 206508 212434
rect 207294 206272 207350 206281
rect 207294 206207 207350 206216
rect 206560 205148 206612 205154
rect 206560 205090 206612 205096
rect 206572 198082 206600 205090
rect 207308 204950 207336 206207
rect 207296 204944 207348 204950
rect 207296 204886 207348 204892
rect 207400 204338 207428 240244
rect 207952 240145 207980 240244
rect 208320 240145 208348 240244
rect 207938 240136 207994 240145
rect 207938 240071 207994 240080
rect 208306 240136 208362 240145
rect 208306 240071 208362 240080
rect 207952 237454 207980 240071
rect 208320 238241 208348 240071
rect 208306 238232 208362 238241
rect 208306 238167 208362 238176
rect 207940 237448 207992 237454
rect 207940 237390 207992 237396
rect 208872 235793 208900 240244
rect 209240 238754 209268 240244
rect 208964 238726 209268 238754
rect 208858 235784 208914 235793
rect 208858 235719 208914 235728
rect 208872 234977 208900 235719
rect 208858 234968 208914 234977
rect 208858 234903 208914 234912
rect 208964 227633 208992 238726
rect 209042 237280 209098 237289
rect 209042 237215 209098 237224
rect 208950 227624 209006 227633
rect 208950 227559 209006 227568
rect 207940 222216 207992 222222
rect 207940 222158 207992 222164
rect 207952 216073 207980 222158
rect 208964 221921 208992 227559
rect 208950 221912 209006 221921
rect 208950 221847 209006 221856
rect 207938 216064 207994 216073
rect 207938 215999 207994 216008
rect 207754 215384 207810 215393
rect 207754 215319 207810 215328
rect 207020 204332 207072 204338
rect 207020 204274 207072 204280
rect 207388 204332 207440 204338
rect 207388 204274 207440 204280
rect 207032 202842 207060 204274
rect 207020 202836 207072 202842
rect 207020 202778 207072 202784
rect 206560 198076 206612 198082
rect 206560 198018 206612 198024
rect 206560 195356 206612 195362
rect 206560 195298 206612 195304
rect 206468 195288 206520 195294
rect 206468 195230 206520 195236
rect 206376 188420 206428 188426
rect 206376 188362 206428 188368
rect 206572 181665 206600 195298
rect 207018 187232 207074 187241
rect 207018 187167 207074 187176
rect 207032 184890 207060 187167
rect 207020 184884 207072 184890
rect 207020 184826 207072 184832
rect 206558 181656 206614 181665
rect 206558 181591 206614 181600
rect 207768 177449 207796 215319
rect 209056 206281 209084 237215
rect 209226 234968 209282 234977
rect 209226 234903 209282 234912
rect 209240 206281 209268 234903
rect 209792 215257 209820 240244
rect 209870 239456 209926 239465
rect 209870 239391 209926 239400
rect 209884 238377 209912 239391
rect 210344 238754 210372 240244
rect 210712 240145 210740 240244
rect 210698 240136 210754 240145
rect 210698 240071 210754 240080
rect 210344 238726 210464 238754
rect 209870 238368 209926 238377
rect 209870 238303 209926 238312
rect 209962 237416 210018 237425
rect 209962 237351 210018 237360
rect 209778 215248 209834 215257
rect 209778 215183 209834 215192
rect 209042 206272 209098 206281
rect 209042 206207 209098 206216
rect 209226 206272 209282 206281
rect 209226 206207 209282 206216
rect 209976 205465 210004 237351
rect 210436 234569 210464 238726
rect 210712 237425 210740 240071
rect 211264 238649 211292 240244
rect 211816 238754 211844 240244
rect 211448 238726 211844 238754
rect 211250 238640 211306 238649
rect 211250 238575 211306 238584
rect 211264 237425 211292 238575
rect 210698 237416 210754 237425
rect 210698 237351 210754 237360
rect 211250 237416 211306 237425
rect 211250 237351 211306 237360
rect 210422 234560 210478 234569
rect 210422 234495 210478 234504
rect 210436 220153 210464 234495
rect 211448 224330 211476 238726
rect 211804 229152 211856 229158
rect 211804 229094 211856 229100
rect 212184 229094 212212 240244
rect 212736 238754 212764 240244
rect 213104 240145 213132 240244
rect 213090 240136 213146 240145
rect 213090 240071 213146 240080
rect 211068 224324 211120 224330
rect 211068 224266 211120 224272
rect 211436 224324 211488 224330
rect 211436 224266 211488 224272
rect 210422 220144 210478 220153
rect 210422 220079 210478 220088
rect 210514 215248 210570 215257
rect 210514 215183 210570 215192
rect 209962 205456 210018 205465
rect 209962 205391 210018 205400
rect 210422 205456 210478 205465
rect 210422 205391 210478 205400
rect 209042 203552 209098 203561
rect 209042 203487 209098 203496
rect 207754 177440 207810 177449
rect 207664 177404 207716 177410
rect 207754 177375 207810 177384
rect 207664 177346 207716 177352
rect 206374 136776 206430 136785
rect 206374 136711 206430 136720
rect 206388 89622 206416 136711
rect 206468 133204 206520 133210
rect 206468 133146 206520 133152
rect 206480 91905 206508 133146
rect 206466 91896 206522 91905
rect 206466 91831 206522 91840
rect 206376 89616 206428 89622
rect 206376 89558 206428 89564
rect 206282 86320 206338 86329
rect 206282 86255 206338 86264
rect 207676 83502 207704 177346
rect 207756 113212 207808 113218
rect 207756 113154 207808 113160
rect 207768 85513 207796 113154
rect 207754 85504 207810 85513
rect 207754 85439 207810 85448
rect 207664 83496 207716 83502
rect 207664 83438 207716 83444
rect 206284 82136 206336 82142
rect 206284 82078 206336 82084
rect 205180 49700 205232 49706
rect 205180 49642 205232 49648
rect 204904 29708 204956 29714
rect 204904 29650 204956 29656
rect 202236 9036 202288 9042
rect 202236 8978 202288 8984
rect 206296 7682 206324 82078
rect 206284 7676 206336 7682
rect 206284 7618 206336 7624
rect 191104 6248 191156 6254
rect 191104 6190 191156 6196
rect 209056 3369 209084 203487
rect 209228 147688 209280 147694
rect 209228 147630 209280 147636
rect 209240 130422 209268 147630
rect 209228 130416 209280 130422
rect 209228 130358 209280 130364
rect 209136 129804 209188 129810
rect 209136 129746 209188 129752
rect 209148 59362 209176 129746
rect 209226 115152 209282 115161
rect 209226 115087 209282 115096
rect 209240 91089 209268 115087
rect 210436 96762 210464 205391
rect 210528 203561 210556 215183
rect 210514 203552 210570 203561
rect 210514 203487 210570 203496
rect 211080 202162 211108 224266
rect 211068 202156 211120 202162
rect 211068 202098 211120 202104
rect 211816 185745 211844 229094
rect 212000 229066 212212 229094
rect 212552 238726 212764 238754
rect 212000 219502 212028 229066
rect 212448 224256 212500 224262
rect 212448 224198 212500 224204
rect 212460 220726 212488 224198
rect 212448 220720 212500 220726
rect 212448 220662 212500 220668
rect 211988 219496 212040 219502
rect 211988 219438 212040 219444
rect 211896 208072 211948 208078
rect 211896 208014 211948 208020
rect 211802 185736 211858 185745
rect 211802 185671 211858 185680
rect 211908 182170 211936 208014
rect 212000 201482 212028 219438
rect 212552 213246 212580 238726
rect 213104 219434 213132 240071
rect 212736 219406 213132 219434
rect 212540 213240 212592 213246
rect 212540 213182 212592 213188
rect 212540 211064 212592 211070
rect 212540 211006 212592 211012
rect 212552 210458 212580 211006
rect 212540 210452 212592 210458
rect 212540 210394 212592 210400
rect 212552 209774 212580 210394
rect 212460 209746 212580 209774
rect 212736 209774 212764 219406
rect 213460 213920 213512 213926
rect 213460 213862 213512 213868
rect 213472 213246 213500 213862
rect 213460 213240 213512 213246
rect 213460 213182 213512 213188
rect 213656 211070 213684 240244
rect 214208 240145 214236 240244
rect 214194 240136 214250 240145
rect 214194 240071 214250 240080
rect 213826 239592 213882 239601
rect 213826 239527 213882 239536
rect 213840 238513 213868 239527
rect 213826 238504 213882 238513
rect 213826 238439 213882 238448
rect 214208 238377 214236 240071
rect 214194 238368 214250 238377
rect 214194 238303 214250 238312
rect 214208 237454 214236 238303
rect 214196 237448 214248 237454
rect 214196 237390 214248 237396
rect 213826 217424 213882 217433
rect 213826 217359 213882 217368
rect 213644 211064 213696 211070
rect 213840 211041 213868 217359
rect 214576 216578 214604 240244
rect 214656 237448 214708 237454
rect 214656 237390 214708 237396
rect 214564 216572 214616 216578
rect 214564 216514 214616 216520
rect 213644 211006 213696 211012
rect 213826 211032 213882 211041
rect 213826 210967 213882 210976
rect 212736 209746 213224 209774
rect 212460 207738 212488 209746
rect 213196 208321 213224 209746
rect 213182 208312 213238 208321
rect 213182 208247 213238 208256
rect 212448 207732 212500 207738
rect 212448 207674 212500 207680
rect 211988 201476 212040 201482
rect 211988 201418 212040 201424
rect 211896 182164 211948 182170
rect 211896 182106 211948 182112
rect 211804 180872 211856 180878
rect 211804 180814 211856 180820
rect 210514 174584 210570 174593
rect 210514 174519 210570 174528
rect 210528 171018 210556 174519
rect 211816 173806 211844 180814
rect 211804 173800 211856 173806
rect 211804 173742 211856 173748
rect 210516 171012 210568 171018
rect 210516 170954 210568 170960
rect 211896 153332 211948 153338
rect 211896 153274 211948 153280
rect 211804 132592 211856 132598
rect 211804 132534 211856 132540
rect 210514 131336 210570 131345
rect 210514 131271 210570 131280
rect 210424 96756 210476 96762
rect 210424 96698 210476 96704
rect 209226 91080 209282 91089
rect 209226 91015 209282 91024
rect 210528 60722 210556 131271
rect 210608 128376 210660 128382
rect 210608 128318 210660 128324
rect 210620 82793 210648 128318
rect 210606 82784 210662 82793
rect 210606 82719 210662 82728
rect 210516 60716 210568 60722
rect 210516 60658 210568 60664
rect 209136 59356 209188 59362
rect 209136 59298 209188 59304
rect 211816 57934 211844 132534
rect 211908 126274 211936 153274
rect 211988 152108 212040 152114
rect 211988 152050 212040 152056
rect 212000 131782 212028 152050
rect 211988 131776 212040 131782
rect 211988 131718 212040 131724
rect 211896 126268 211948 126274
rect 211896 126210 211948 126216
rect 213196 96014 213224 208247
rect 214472 206916 214524 206922
rect 214472 206858 214524 206864
rect 214484 205737 214512 206858
rect 214470 205728 214526 205737
rect 214470 205663 214472 205672
rect 214524 205663 214526 205672
rect 214472 205634 214524 205640
rect 214668 200802 214696 237390
rect 215128 234734 215156 240244
rect 215680 237454 215708 240244
rect 215668 237448 215720 237454
rect 215668 237390 215720 237396
rect 214748 234728 214800 234734
rect 214748 234670 214800 234676
rect 215116 234728 215168 234734
rect 215116 234670 215168 234676
rect 214760 230450 214788 234670
rect 214748 230444 214800 230450
rect 214748 230386 214800 230392
rect 215944 225616 215996 225622
rect 215944 225558 215996 225564
rect 215956 225049 215984 225558
rect 215942 225040 215998 225049
rect 215942 224975 215998 224984
rect 215298 216064 215354 216073
rect 215298 215999 215354 216008
rect 215312 214577 215340 215999
rect 215298 214568 215354 214577
rect 215298 214503 215354 214512
rect 215300 204332 215352 204338
rect 215300 204274 215352 204280
rect 215312 203590 215340 204274
rect 215300 203584 215352 203590
rect 215300 203526 215352 203532
rect 214656 200796 214708 200802
rect 214656 200738 214708 200744
rect 215300 185700 215352 185706
rect 215300 185642 215352 185648
rect 215312 185065 215340 185642
rect 215298 185056 215354 185065
rect 215298 184991 215354 185000
rect 215956 182850 215984 224975
rect 216048 206961 216076 240244
rect 216496 237448 216548 237454
rect 216600 237425 216628 240244
rect 216496 237390 216548 237396
rect 216586 237416 216642 237425
rect 216034 206952 216090 206961
rect 216034 206887 216090 206896
rect 216508 205698 216536 237390
rect 216586 237351 216642 237360
rect 216770 237416 216826 237425
rect 216770 237351 216826 237360
rect 216784 209778 216812 237351
rect 217152 220794 217180 240244
rect 217520 240145 217548 240244
rect 217506 240136 217562 240145
rect 217506 240071 217562 240080
rect 217520 237425 217548 240071
rect 217506 237416 217562 237425
rect 217506 237351 217562 237360
rect 217324 229764 217376 229770
rect 217324 229706 217376 229712
rect 217140 220788 217192 220794
rect 217140 220730 217192 220736
rect 217152 216073 217180 220730
rect 217336 219366 217364 229706
rect 218072 222057 218100 240244
rect 218150 234696 218206 234705
rect 218150 234631 218206 234640
rect 218164 234530 218192 234631
rect 218152 234524 218204 234530
rect 218152 234466 218204 234472
rect 218150 230344 218206 230353
rect 218150 230279 218206 230288
rect 218164 229129 218192 230279
rect 218150 229120 218206 229129
rect 218150 229055 218206 229064
rect 218164 228313 218192 229055
rect 218150 228304 218206 228313
rect 218150 228239 218206 228248
rect 218058 222048 218114 222057
rect 218058 221983 218114 221992
rect 217324 219360 217376 219366
rect 217324 219302 217376 219308
rect 218072 218657 218100 221983
rect 218058 218648 218114 218657
rect 218058 218583 218114 218592
rect 217138 216064 217194 216073
rect 217138 215999 217194 216008
rect 217416 214600 217468 214606
rect 217416 214542 217468 214548
rect 216772 209772 216824 209778
rect 216772 209714 216824 209720
rect 216036 205692 216088 205698
rect 216036 205634 216088 205640
rect 216128 205692 216180 205698
rect 216128 205634 216180 205640
rect 216496 205692 216548 205698
rect 216496 205634 216548 205640
rect 216048 199481 216076 205634
rect 216140 204270 216168 205634
rect 216128 204264 216180 204270
rect 216128 204206 216180 204212
rect 216784 200977 216812 209714
rect 217428 209098 217456 214542
rect 218440 211070 218468 240244
rect 218992 240145 219020 240244
rect 218978 240136 219034 240145
rect 218978 240071 219034 240080
rect 218992 230353 219020 240071
rect 219544 231713 219572 240244
rect 219912 238678 219940 240244
rect 220464 238754 220492 240244
rect 220728 240168 220780 240174
rect 220912 240168 220964 240174
rect 220728 240110 220780 240116
rect 220910 240136 220912 240145
rect 220964 240136 220966 240145
rect 220740 239873 220768 240110
rect 220910 240071 220966 240080
rect 220726 239864 220782 239873
rect 220726 239799 220782 239808
rect 220096 238726 220492 238754
rect 219900 238672 219952 238678
rect 219900 238614 219952 238620
rect 219912 234530 219940 238614
rect 219900 234524 219952 234530
rect 219900 234466 219952 234472
rect 219530 231704 219586 231713
rect 219530 231639 219586 231648
rect 218978 230344 219034 230353
rect 218978 230279 219034 230288
rect 220096 229022 220124 238726
rect 221016 233209 221044 240244
rect 221002 233200 221058 233209
rect 221002 233135 221058 233144
rect 220358 231704 220414 231713
rect 220358 231639 220414 231648
rect 220174 231296 220230 231305
rect 220174 231231 220230 231240
rect 220084 229016 220136 229022
rect 220084 228958 220136 228964
rect 218428 211064 218480 211070
rect 218428 211006 218480 211012
rect 218796 211064 218848 211070
rect 218796 211006 218848 211012
rect 217416 209092 217468 209098
rect 217416 209034 217468 209040
rect 216770 200968 216826 200977
rect 216770 200903 216826 200912
rect 218704 200864 218756 200870
rect 218704 200806 218756 200812
rect 216034 199472 216090 199481
rect 216034 199407 216090 199416
rect 217324 199436 217376 199442
rect 217324 199378 217376 199384
rect 217336 185881 217364 199378
rect 217322 185872 217378 185881
rect 217322 185807 217378 185816
rect 216036 185632 216088 185638
rect 216036 185574 216088 185580
rect 215116 182844 215168 182850
rect 215116 182786 215168 182792
rect 215944 182844 215996 182850
rect 215944 182786 215996 182792
rect 214196 179444 214248 179450
rect 214196 179386 214248 179392
rect 213920 176656 213972 176662
rect 213920 176598 213972 176604
rect 213932 175681 213960 176598
rect 213918 175672 213974 175681
rect 213918 175607 213974 175616
rect 214102 175536 214158 175545
rect 214102 175471 214158 175480
rect 214012 175228 214064 175234
rect 214012 175170 214064 175176
rect 213920 175160 213972 175166
rect 213920 175102 213972 175108
rect 213932 175001 213960 175102
rect 213918 174992 213974 175001
rect 213918 174927 213974 174936
rect 214024 174321 214052 175170
rect 214010 174312 214066 174321
rect 214010 174247 214066 174256
rect 213920 173868 213972 173874
rect 213920 173810 213972 173816
rect 213932 172961 213960 173810
rect 213918 172952 213974 172961
rect 213918 172887 213974 172896
rect 214116 171601 214144 175471
rect 214208 172281 214236 179386
rect 215128 178770 215156 182786
rect 215944 179444 215996 179450
rect 215944 179386 215996 179392
rect 215116 178764 215168 178770
rect 215116 178706 215168 178712
rect 214562 177168 214618 177177
rect 214562 177103 214618 177112
rect 214472 173800 214524 173806
rect 214472 173742 214524 173748
rect 214484 173641 214512 173742
rect 214470 173632 214526 173641
rect 214470 173567 214526 173576
rect 214194 172272 214250 172281
rect 214194 172207 214250 172216
rect 214102 171592 214158 171601
rect 214102 171527 214158 171536
rect 213920 171080 213972 171086
rect 213920 171022 213972 171028
rect 214010 171048 214066 171057
rect 213932 170377 213960 171022
rect 214010 170983 214012 170992
rect 214064 170983 214066 170992
rect 214012 170954 214064 170960
rect 213918 170368 213974 170377
rect 213918 170303 213974 170312
rect 214012 169720 214064 169726
rect 213918 169688 213974 169697
rect 214012 169662 214064 169668
rect 213918 169623 213920 169632
rect 213972 169623 213974 169632
rect 213920 169594 213972 169600
rect 214024 169017 214052 169662
rect 214010 169008 214066 169017
rect 214010 168943 214066 168952
rect 213920 168360 213972 168366
rect 213918 168328 213920 168337
rect 213972 168328 213974 168337
rect 213918 168263 213974 168272
rect 214012 168292 214064 168298
rect 214012 168234 214064 168240
rect 214024 167657 214052 168234
rect 214010 167648 214066 167657
rect 214010 167583 214066 167592
rect 214012 167000 214064 167006
rect 213918 166968 213974 166977
rect 214012 166942 214064 166948
rect 213918 166903 213920 166912
rect 213972 166903 213974 166912
rect 213920 166874 213972 166880
rect 214024 166433 214052 166942
rect 214010 166424 214066 166433
rect 214010 166359 214066 166368
rect 213920 165572 213972 165578
rect 213920 165514 213972 165520
rect 213932 165073 213960 165514
rect 213918 165064 213974 165073
rect 213918 164999 213974 165008
rect 214012 164212 214064 164218
rect 214012 164154 214064 164160
rect 213920 164144 213972 164150
rect 213920 164086 213972 164092
rect 213932 163713 213960 164086
rect 213918 163704 213974 163713
rect 213918 163639 213974 163648
rect 214024 163033 214052 164154
rect 214010 163024 214066 163033
rect 214010 162959 214066 162968
rect 213920 162852 213972 162858
rect 213920 162794 213972 162800
rect 213932 162353 213960 162794
rect 214012 162784 214064 162790
rect 214012 162726 214064 162732
rect 213918 162344 213974 162353
rect 213918 162279 213974 162288
rect 214024 161809 214052 162726
rect 214010 161800 214066 161809
rect 214010 161735 214066 161744
rect 214012 161424 214064 161430
rect 214012 161366 214064 161372
rect 213920 161356 213972 161362
rect 213920 161298 213972 161304
rect 213932 161129 213960 161298
rect 213918 161120 213974 161129
rect 213918 161055 213974 161064
rect 214024 160449 214052 161366
rect 214010 160440 214066 160449
rect 214010 160375 214066 160384
rect 213920 160064 213972 160070
rect 213920 160006 213972 160012
rect 213932 159769 213960 160006
rect 213918 159760 213974 159769
rect 213918 159695 213974 159704
rect 214576 159089 214604 177103
rect 215482 175944 215538 175953
rect 215482 175879 215538 175888
rect 215392 175296 215444 175302
rect 215392 175238 215444 175244
rect 215300 173936 215352 173942
rect 215404 173913 215432 175238
rect 215300 173878 215352 173884
rect 215390 173904 215446 173913
rect 215206 173224 215262 173233
rect 215206 173159 215262 173168
rect 215220 164393 215248 173159
rect 215312 172514 215340 173878
rect 215390 173839 215446 173848
rect 215300 172508 215352 172514
rect 215300 172450 215352 172456
rect 215496 172417 215524 175879
rect 215482 172408 215538 172417
rect 215482 172343 215538 172352
rect 215956 170921 215984 179386
rect 216048 177585 216076 185574
rect 216770 179480 216826 179489
rect 216770 179415 216826 179424
rect 216678 178120 216734 178129
rect 216678 178055 216734 178064
rect 216034 177576 216090 177585
rect 216034 177511 216090 177520
rect 216692 176633 216720 178055
rect 216678 176624 216734 176633
rect 216678 176559 216734 176568
rect 216784 172446 216812 179415
rect 218716 175982 218744 200806
rect 218808 198014 218836 211006
rect 218796 198008 218848 198014
rect 218796 197950 218848 197956
rect 218794 187776 218850 187785
rect 218794 187711 218850 187720
rect 218808 180810 218836 187711
rect 218796 180804 218848 180810
rect 218796 180746 218848 180752
rect 220096 180130 220124 228958
rect 220188 194546 220216 231231
rect 220372 198014 220400 231639
rect 221384 219366 221412 240244
rect 221936 238754 221964 240244
rect 221476 238726 221964 238754
rect 222304 238746 222332 240244
rect 222292 238740 222344 238746
rect 221476 237289 221504 238726
rect 222292 238682 222344 238688
rect 221462 237280 221518 237289
rect 221462 237215 221518 237224
rect 221372 219360 221424 219366
rect 221372 219302 221424 219308
rect 220360 198008 220412 198014
rect 220360 197950 220412 197956
rect 220176 194540 220228 194546
rect 220176 194482 220228 194488
rect 221476 191146 221504 237215
rect 222856 233238 222884 240244
rect 223304 240168 223356 240174
rect 223408 240122 223436 240244
rect 223356 240116 223436 240122
rect 223304 240110 223436 240116
rect 223316 240094 223436 240110
rect 223408 238754 223436 240094
rect 223408 238726 223528 238754
rect 222844 233232 222896 233238
rect 221646 233200 221702 233209
rect 223396 233232 223448 233238
rect 222844 233174 222896 233180
rect 223394 233200 223396 233209
rect 223448 233200 223450 233209
rect 221646 233135 221702 233144
rect 223394 233135 223450 233144
rect 221660 227662 221688 233135
rect 221648 227656 221700 227662
rect 221648 227598 221700 227604
rect 221556 227044 221608 227050
rect 221556 226986 221608 226992
rect 221568 196722 221596 226986
rect 221646 225720 221702 225729
rect 221646 225655 221702 225664
rect 221660 197334 221688 225655
rect 222384 215280 222436 215286
rect 222382 215248 222384 215257
rect 223396 215280 223448 215286
rect 222436 215248 222438 215257
rect 223396 215222 223448 215228
rect 222382 215183 222438 215192
rect 223408 213994 223436 215222
rect 223396 213988 223448 213994
rect 223396 213930 223448 213936
rect 223394 211168 223450 211177
rect 223394 211103 223450 211112
rect 223408 210361 223436 211103
rect 223394 210352 223450 210361
rect 223394 210287 223450 210296
rect 223408 209166 223436 210287
rect 223396 209160 223448 209166
rect 223396 209102 223448 209108
rect 221648 197328 221700 197334
rect 221648 197270 221700 197276
rect 221556 196716 221608 196722
rect 221556 196658 221608 196664
rect 223500 193934 223528 238726
rect 223776 235890 223804 240244
rect 224328 240145 224356 240244
rect 224314 240136 224370 240145
rect 224314 240071 224370 240080
rect 224328 237425 224356 240071
rect 224408 239420 224460 239426
rect 224408 239362 224460 239368
rect 224314 237416 224370 237425
rect 224314 237351 224370 237360
rect 223764 235884 223816 235890
rect 223764 235826 223816 235832
rect 223776 234666 223804 235826
rect 223764 234660 223816 234666
rect 223764 234602 223816 234608
rect 224224 234660 224276 234666
rect 224224 234602 224276 234608
rect 223488 193928 223540 193934
rect 223488 193870 223540 193876
rect 221464 191140 221516 191146
rect 221464 191082 221516 191088
rect 224236 190454 224264 234602
rect 224420 231810 224448 239362
rect 224774 238776 224830 238785
rect 224774 238711 224830 238720
rect 224788 238066 224816 238711
rect 224776 238060 224828 238066
rect 224776 238002 224828 238008
rect 224408 231804 224460 231810
rect 224408 231746 224460 231752
rect 224408 228404 224460 228410
rect 224408 228346 224460 228352
rect 224316 223576 224368 223582
rect 224316 223518 224368 223524
rect 224328 200870 224356 223518
rect 224420 215937 224448 228346
rect 224880 223582 224908 240244
rect 224868 223576 224920 223582
rect 224868 223518 224920 223524
rect 225248 217977 225276 240244
rect 225800 231169 225828 240244
rect 226168 234705 226196 240244
rect 226720 238513 226748 240244
rect 226706 238504 226762 238513
rect 226706 238439 226762 238448
rect 226720 237969 226748 238439
rect 226706 237960 226762 237969
rect 226706 237895 226762 237904
rect 226984 236020 227036 236026
rect 226984 235962 227036 235968
rect 226154 234696 226210 234705
rect 226154 234631 226210 234640
rect 226168 232558 226196 234631
rect 226156 232552 226208 232558
rect 226156 232494 226208 232500
rect 225786 231160 225842 231169
rect 225786 231095 225842 231104
rect 225800 219434 225828 231095
rect 225708 219406 225828 219434
rect 225234 217968 225290 217977
rect 225234 217903 225290 217912
rect 225248 215937 225276 217903
rect 225602 217424 225658 217433
rect 225602 217359 225658 217368
rect 224406 215928 224462 215937
rect 224406 215863 224462 215872
rect 225234 215928 225290 215937
rect 225234 215863 225290 215872
rect 224316 200864 224368 200870
rect 224316 200806 224368 200812
rect 225616 190466 225644 217359
rect 225708 209545 225736 219406
rect 225694 209536 225750 209545
rect 225694 209471 225750 209480
rect 225694 200968 225750 200977
rect 225694 200903 225750 200912
rect 225604 190460 225656 190466
rect 224236 190426 224356 190454
rect 224224 189100 224276 189106
rect 224224 189042 224276 189048
rect 224236 186318 224264 189042
rect 224224 186312 224276 186318
rect 224224 186254 224276 186260
rect 224328 182918 224356 190426
rect 225604 190402 225656 190408
rect 225708 184521 225736 200903
rect 226340 193248 226392 193254
rect 226340 193190 226392 193196
rect 226352 191826 226380 193190
rect 226340 191820 226392 191826
rect 226340 191762 226392 191768
rect 226340 185632 226392 185638
rect 226340 185574 226392 185580
rect 226352 184890 226380 185574
rect 226340 184884 226392 184890
rect 226340 184826 226392 184832
rect 225694 184512 225750 184521
rect 225694 184447 225750 184456
rect 224316 182912 224368 182918
rect 224316 182854 224368 182860
rect 226996 180878 227024 235962
rect 227272 229770 227300 240244
rect 227260 229764 227312 229770
rect 227260 229706 227312 229712
rect 227640 219337 227668 240244
rect 228192 222057 228220 240244
rect 228362 240136 228418 240145
rect 228744 240106 228772 240244
rect 228362 240071 228418 240080
rect 228732 240100 228784 240106
rect 228178 222048 228234 222057
rect 228178 221983 228234 221992
rect 227626 219328 227682 219337
rect 227626 219263 227682 219272
rect 227640 218113 227668 219263
rect 227074 218104 227130 218113
rect 227074 218039 227130 218048
rect 227626 218104 227682 218113
rect 227626 218039 227682 218048
rect 227088 203697 227116 218039
rect 227074 203688 227130 203697
rect 227074 203623 227130 203632
rect 227720 203652 227772 203658
rect 227720 203594 227772 203600
rect 227076 193860 227128 193866
rect 227076 193802 227128 193808
rect 226984 180872 227036 180878
rect 226984 180814 227036 180820
rect 227088 180305 227116 193802
rect 227074 180296 227130 180305
rect 227074 180231 227130 180240
rect 226338 180160 226394 180169
rect 220084 180124 220136 180130
rect 226338 180095 226394 180104
rect 220084 180066 220136 180072
rect 226352 177614 226380 180095
rect 226340 177608 226392 177614
rect 226340 177550 226392 177556
rect 226246 176760 226302 176769
rect 226246 176695 226302 176704
rect 218704 175976 218756 175982
rect 226260 175953 226288 176695
rect 227732 176225 227760 203594
rect 227812 185700 227864 185706
rect 227812 185642 227864 185648
rect 227824 185065 227852 185642
rect 227810 185056 227866 185065
rect 227810 184991 227866 185000
rect 227718 176216 227774 176225
rect 227718 176151 227774 176160
rect 228376 176050 228404 240071
rect 228732 240042 228784 240048
rect 228744 219434 228772 240042
rect 229112 238105 229140 240244
rect 229098 238096 229154 238105
rect 229098 238031 229154 238040
rect 228468 219406 228772 219434
rect 228468 215121 228496 219406
rect 228454 215112 228510 215121
rect 228454 215047 228510 215056
rect 229664 213897 229692 240244
rect 230216 234666 230244 240244
rect 230584 240145 230612 240244
rect 230570 240136 230626 240145
rect 230570 240071 230626 240080
rect 230478 238096 230534 238105
rect 230478 238031 230534 238040
rect 230204 234660 230256 234666
rect 230204 234602 230256 234608
rect 230388 229764 230440 229770
rect 230388 229706 230440 229712
rect 229650 213888 229706 213897
rect 229650 213823 229706 213832
rect 229192 207664 229244 207670
rect 229192 207606 229244 207612
rect 229204 180794 229232 207606
rect 230400 206825 230428 229706
rect 230492 213625 230520 238031
rect 230584 237425 230612 240071
rect 230570 237416 230626 237425
rect 230570 237351 230626 237360
rect 231136 229770 231164 240244
rect 231504 234569 231532 240244
rect 232056 240122 232084 240244
rect 232136 240168 232188 240174
rect 232056 240116 232136 240122
rect 232056 240110 232188 240116
rect 232502 240136 232558 240145
rect 232056 240094 232176 240110
rect 232056 239426 232084 240094
rect 232502 240071 232558 240080
rect 232044 239420 232096 239426
rect 232044 239362 232096 239368
rect 231766 237416 231822 237425
rect 231766 237351 231822 237360
rect 231490 234560 231546 234569
rect 231490 234495 231546 234504
rect 231124 229764 231176 229770
rect 231124 229706 231176 229712
rect 231504 219434 231532 234495
rect 231136 219406 231532 219434
rect 231136 218006 231164 219406
rect 231124 218000 231176 218006
rect 231124 217942 231176 217948
rect 230478 213616 230534 213625
rect 230478 213551 230534 213560
rect 230386 206816 230442 206825
rect 230386 206751 230442 206760
rect 230664 192500 230716 192506
rect 230664 192442 230716 192448
rect 229284 180872 229336 180878
rect 229284 180814 229336 180820
rect 229112 180766 229232 180794
rect 228364 176044 228416 176050
rect 228364 175986 228416 175992
rect 218704 175918 218756 175924
rect 226246 175944 226302 175953
rect 226246 175879 226302 175888
rect 229006 175944 229062 175953
rect 229006 175879 229062 175888
rect 229020 175302 229048 175879
rect 229008 175296 229060 175302
rect 229112 175273 229140 180766
rect 229190 176488 229246 176497
rect 229190 176423 229246 176432
rect 229008 175238 229060 175244
rect 229098 175264 229154 175273
rect 229098 175199 229154 175208
rect 229098 174720 229154 174729
rect 229020 174678 229098 174706
rect 229020 174010 229048 174678
rect 229098 174655 229154 174664
rect 229100 174616 229152 174622
rect 229100 174558 229152 174564
rect 229008 174004 229060 174010
rect 229008 173946 229060 173952
rect 216772 172440 216824 172446
rect 216772 172382 216824 172388
rect 215942 170912 215998 170921
rect 215942 170847 215998 170856
rect 215206 164384 215262 164393
rect 215206 164319 215262 164328
rect 214562 159080 214618 159089
rect 214562 159015 214618 159024
rect 213920 158704 213972 158710
rect 213920 158646 213972 158652
rect 213932 158409 213960 158646
rect 214012 158636 214064 158642
rect 214012 158578 214064 158584
rect 213918 158400 213974 158409
rect 213918 158335 213974 158344
rect 214024 157729 214052 158578
rect 214010 157720 214066 157729
rect 214010 157655 214066 157664
rect 213920 157344 213972 157350
rect 213920 157286 213972 157292
rect 213932 157185 213960 157286
rect 214012 157276 214064 157282
rect 214012 157218 214064 157224
rect 213918 157176 213974 157185
rect 213918 157111 213974 157120
rect 214024 156505 214052 157218
rect 214010 156496 214066 156505
rect 214010 156431 214066 156440
rect 214012 155916 214064 155922
rect 214012 155858 214064 155864
rect 213920 155848 213972 155854
rect 213918 155816 213920 155825
rect 213972 155816 213974 155825
rect 213918 155751 213974 155760
rect 214024 155145 214052 155858
rect 214010 155136 214066 155145
rect 214010 155071 214066 155080
rect 214010 154456 214066 154465
rect 214010 154391 214066 154400
rect 213918 153776 213974 153785
rect 213918 153711 213974 153720
rect 213932 153270 213960 153711
rect 214024 153338 214052 154391
rect 214012 153332 214064 153338
rect 214012 153274 214064 153280
rect 213920 153264 213972 153270
rect 213920 153206 213972 153212
rect 213918 153096 213974 153105
rect 213918 153031 213974 153040
rect 213932 151842 213960 153031
rect 214010 152552 214066 152561
rect 214010 152487 214066 152496
rect 214024 152114 214052 152487
rect 214012 152108 214064 152114
rect 214012 152050 214064 152056
rect 214562 151872 214618 151881
rect 213920 151836 213972 151842
rect 214562 151807 214618 151816
rect 213920 151778 213972 151784
rect 214010 151192 214066 151201
rect 214010 151127 214066 151136
rect 214024 150550 214052 151127
rect 214012 150544 214064 150550
rect 213918 150512 213974 150521
rect 214012 150486 214064 150492
rect 213918 150447 213920 150456
rect 213972 150447 213974 150456
rect 213920 150418 213972 150424
rect 214012 150408 214064 150414
rect 214012 150350 214064 150356
rect 213920 150340 213972 150346
rect 213920 150282 213972 150288
rect 213932 149841 213960 150282
rect 213918 149832 213974 149841
rect 213918 149767 213974 149776
rect 214024 149161 214052 150350
rect 214010 149152 214066 149161
rect 214010 149087 214066 149096
rect 213920 149048 213972 149054
rect 213920 148990 213972 148996
rect 213932 148481 213960 148990
rect 213918 148472 213974 148481
rect 213918 148407 213974 148416
rect 213918 147928 213974 147937
rect 213918 147863 213974 147872
rect 213932 147694 213960 147863
rect 213920 147688 213972 147694
rect 213920 147630 213972 147636
rect 214010 147248 214066 147257
rect 214010 147183 214066 147192
rect 213918 146568 213974 146577
rect 213918 146503 213974 146512
rect 213932 146334 213960 146503
rect 213920 146328 213972 146334
rect 213920 146270 213972 146276
rect 213918 145208 213974 145217
rect 213918 145143 213974 145152
rect 213932 144974 213960 145143
rect 213920 144968 213972 144974
rect 213920 144910 213972 144916
rect 214024 144226 214052 147183
rect 214194 144528 214250 144537
rect 214194 144463 214250 144472
rect 214012 144220 214064 144226
rect 214012 144162 214064 144168
rect 213918 143848 213974 143857
rect 213918 143783 213974 143792
rect 213932 143614 213960 143783
rect 213920 143608 213972 143614
rect 213920 143550 213972 143556
rect 214010 143304 214066 143313
rect 214010 143239 214066 143248
rect 213918 142624 213974 142633
rect 213918 142559 213974 142568
rect 213932 142186 213960 142559
rect 214024 142254 214052 143239
rect 214012 142248 214064 142254
rect 214012 142190 214064 142196
rect 213920 142180 213972 142186
rect 213920 142122 213972 142128
rect 214010 141944 214066 141953
rect 214010 141879 214066 141888
rect 213918 141264 213974 141273
rect 213918 141199 213974 141208
rect 213932 140894 213960 141199
rect 213920 140888 213972 140894
rect 213920 140830 213972 140836
rect 214024 140826 214052 141879
rect 214012 140820 214064 140826
rect 214012 140762 214064 140768
rect 213918 140584 213974 140593
rect 213918 140519 213974 140528
rect 213932 139466 213960 140519
rect 214208 140078 214236 144463
rect 214576 142154 214604 151807
rect 229112 148753 229140 174558
rect 229204 170921 229232 176423
rect 229296 174622 229324 180814
rect 230388 179376 230440 179382
rect 230386 179344 230388 179353
rect 230440 179344 230442 179353
rect 230386 179279 230442 179288
rect 229560 178696 229612 178702
rect 229560 178638 229612 178644
rect 229466 177304 229522 177313
rect 229466 177239 229522 177248
rect 229374 176352 229430 176361
rect 229374 176287 229430 176296
rect 229284 174616 229336 174622
rect 229284 174558 229336 174564
rect 229388 173369 229416 176287
rect 229480 174049 229508 177239
rect 229466 174040 229522 174049
rect 229466 173975 229522 173984
rect 229374 173360 229430 173369
rect 229374 173295 229430 173304
rect 229190 170912 229246 170921
rect 229190 170847 229246 170856
rect 229572 161945 229600 178638
rect 230572 177608 230624 177614
rect 230572 177550 230624 177556
rect 230018 176624 230074 176633
rect 230018 176559 230074 176568
rect 230032 174010 230060 176559
rect 230480 175228 230532 175234
rect 230480 175170 230532 175176
rect 230492 174729 230520 175170
rect 230478 174720 230534 174729
rect 230478 174655 230534 174664
rect 230020 174004 230072 174010
rect 230020 173946 230072 173952
rect 230584 173777 230612 177550
rect 230570 173768 230626 173777
rect 230570 173703 230626 173712
rect 229558 161936 229614 161945
rect 229558 161871 229614 161880
rect 229744 160132 229796 160138
rect 229744 160074 229796 160080
rect 229098 148744 229154 148753
rect 229098 148679 229154 148688
rect 229756 147257 229784 160074
rect 230572 159452 230624 159458
rect 230572 159394 230624 159400
rect 229834 157856 229890 157865
rect 229834 157791 229890 157800
rect 229742 147248 229798 147257
rect 229742 147183 229798 147192
rect 214392 142126 214604 142154
rect 214196 140072 214248 140078
rect 214196 140014 214248 140020
rect 213920 139460 213972 139466
rect 213920 139402 213972 139408
rect 213918 139224 213974 139233
rect 213918 139159 213974 139168
rect 213932 138038 213960 139159
rect 214102 138680 214158 138689
rect 214102 138615 214158 138624
rect 213920 138032 213972 138038
rect 213366 138000 213422 138009
rect 213920 137974 213972 137980
rect 213366 137935 213422 137944
rect 213274 103592 213330 103601
rect 213274 103527 213330 103536
rect 213184 96008 213236 96014
rect 213184 95950 213236 95956
rect 213184 91860 213236 91866
rect 213184 91802 213236 91808
rect 211804 57928 211856 57934
rect 211804 57870 211856 57876
rect 189722 3360 189778 3369
rect 189722 3295 189778 3304
rect 209042 3360 209098 3369
rect 209042 3295 209098 3304
rect 213196 2174 213224 91802
rect 213288 56574 213316 103527
rect 213380 91798 213408 137935
rect 214010 135960 214066 135969
rect 214010 135895 214066 135904
rect 213920 135380 213972 135386
rect 213920 135322 213972 135328
rect 213932 135289 213960 135322
rect 214024 135318 214052 135895
rect 214012 135312 214064 135318
rect 213918 135280 213974 135289
rect 214012 135254 214064 135260
rect 213918 135215 213974 135224
rect 213918 134600 213974 134609
rect 214116 134570 214144 138615
rect 214392 137290 214420 142126
rect 214562 139904 214618 139913
rect 214562 139839 214618 139848
rect 214380 137284 214432 137290
rect 214380 137226 214432 137232
rect 213918 134535 213974 134544
rect 214104 134564 214156 134570
rect 213932 133958 213960 134535
rect 214104 134506 214156 134512
rect 213920 133952 213972 133958
rect 213920 133894 213972 133900
rect 213918 133376 213974 133385
rect 213918 133311 213974 133320
rect 213932 132530 213960 133311
rect 214470 132696 214526 132705
rect 214470 132631 214526 132640
rect 214484 132598 214512 132631
rect 214472 132592 214524 132598
rect 214472 132534 214524 132540
rect 213920 132524 213972 132530
rect 213920 132466 213972 132472
rect 213918 132016 213974 132025
rect 213918 131951 213974 131960
rect 213932 131170 213960 131951
rect 213920 131164 213972 131170
rect 213920 131106 213972 131112
rect 213918 130656 213974 130665
rect 213918 130591 213974 130600
rect 213932 129810 213960 130591
rect 214472 130484 214524 130490
rect 214472 130426 214524 130432
rect 214010 129976 214066 129985
rect 214010 129911 214066 129920
rect 213920 129804 213972 129810
rect 213920 129746 213972 129752
rect 213918 129296 213974 129305
rect 213918 129231 213974 129240
rect 213932 128382 213960 129231
rect 213920 128376 213972 128382
rect 213920 128318 213972 128324
rect 213918 128072 213974 128081
rect 213918 128007 213974 128016
rect 213932 127022 213960 128007
rect 213920 127016 213972 127022
rect 213920 126958 213972 126964
rect 213918 126032 213974 126041
rect 213918 125967 213974 125976
rect 213932 125662 213960 125967
rect 213920 125656 213972 125662
rect 213920 125598 213972 125604
rect 213918 125352 213974 125361
rect 213918 125287 213974 125296
rect 213932 124234 213960 125287
rect 214024 124914 214052 129911
rect 214102 128752 214158 128761
rect 214102 128687 214158 128696
rect 214012 124908 214064 124914
rect 214012 124850 214064 124856
rect 213920 124228 213972 124234
rect 213920 124170 213972 124176
rect 214010 124128 214066 124137
rect 214010 124063 214066 124072
rect 213918 123448 213974 123457
rect 213918 123383 213974 123392
rect 213932 122874 213960 123383
rect 214024 122942 214052 124063
rect 214116 123593 214144 128687
rect 214102 123584 214158 123593
rect 214102 123519 214158 123528
rect 214012 122936 214064 122942
rect 214012 122878 214064 122884
rect 213920 122868 213972 122874
rect 213920 122810 213972 122816
rect 214484 122834 214512 130426
rect 214576 127634 214604 139839
rect 229744 136672 229796 136678
rect 215942 136640 215998 136649
rect 229744 136614 229796 136620
rect 215942 136575 215998 136584
rect 214564 127628 214616 127634
rect 214564 127570 214616 127576
rect 214746 126712 214802 126721
rect 214746 126647 214802 126656
rect 214484 122806 214604 122834
rect 214010 122768 214066 122777
rect 214010 122703 214066 122712
rect 213918 122088 213974 122097
rect 213918 122023 213974 122032
rect 213932 121582 213960 122023
rect 213920 121576 213972 121582
rect 213920 121518 213972 121524
rect 214024 121514 214052 122703
rect 214012 121508 214064 121514
rect 214012 121450 214064 121456
rect 214010 121408 214066 121417
rect 214010 121343 214066 121352
rect 213918 120728 213974 120737
rect 213918 120663 213974 120672
rect 213932 120154 213960 120663
rect 214024 120222 214052 121343
rect 214012 120216 214064 120222
rect 214012 120158 214064 120164
rect 213920 120148 213972 120154
rect 213920 120090 213972 120096
rect 214010 120048 214066 120057
rect 214010 119983 214066 119992
rect 213918 119504 213974 119513
rect 213918 119439 213974 119448
rect 213932 118794 213960 119439
rect 213920 118788 213972 118794
rect 213920 118730 213972 118736
rect 214024 118726 214052 119983
rect 214012 118720 214064 118726
rect 214012 118662 214064 118668
rect 214010 118144 214066 118153
rect 214010 118079 214066 118088
rect 213918 117464 213974 117473
rect 213918 117399 213920 117408
rect 213972 117399 213974 117408
rect 213920 117370 213972 117376
rect 214024 117366 214052 118079
rect 214012 117360 214064 117366
rect 214012 117302 214064 117308
rect 214010 116784 214066 116793
rect 214010 116719 214066 116728
rect 213918 116104 213974 116113
rect 213918 116039 213920 116048
rect 213972 116039 213974 116048
rect 213920 116010 213972 116016
rect 214024 116006 214052 116719
rect 214012 116000 214064 116006
rect 214012 115942 214064 115948
rect 214010 115424 214066 115433
rect 214010 115359 214066 115368
rect 213918 114880 213974 114889
rect 213918 114815 213974 114824
rect 213932 114646 213960 114815
rect 213920 114640 213972 114646
rect 213920 114582 213972 114588
rect 214024 114578 214052 115359
rect 214012 114572 214064 114578
rect 214012 114514 214064 114520
rect 213918 114200 213974 114209
rect 213918 114135 213974 114144
rect 213932 113218 213960 114135
rect 213920 113212 213972 113218
rect 213920 113154 213972 113160
rect 214010 112840 214066 112849
rect 214010 112775 214066 112784
rect 213918 112160 213974 112169
rect 213918 112095 213974 112104
rect 213932 111858 213960 112095
rect 214024 111926 214052 112775
rect 214012 111920 214064 111926
rect 214012 111862 214064 111868
rect 213920 111852 213972 111858
rect 213920 111794 213972 111800
rect 214010 111480 214066 111489
rect 214010 111415 214066 111424
rect 213918 110800 213974 110809
rect 213918 110735 213974 110744
rect 213932 110566 213960 110735
rect 213920 110560 213972 110566
rect 213920 110502 213972 110508
rect 214024 110498 214052 111415
rect 214012 110492 214064 110498
rect 214012 110434 214064 110440
rect 214010 110256 214066 110265
rect 214010 110191 214066 110200
rect 213918 109576 213974 109585
rect 213918 109511 213974 109520
rect 213932 109070 213960 109511
rect 214024 109138 214052 110191
rect 214012 109132 214064 109138
rect 214012 109074 214064 109080
rect 213920 109064 213972 109070
rect 213920 109006 213972 109012
rect 214010 108896 214066 108905
rect 214010 108831 214066 108840
rect 213918 108216 213974 108225
rect 213918 108151 213974 108160
rect 213932 107778 213960 108151
rect 213920 107772 213972 107778
rect 213920 107714 213972 107720
rect 214024 107710 214052 108831
rect 214012 107704 214064 107710
rect 214012 107646 214064 107652
rect 214010 107536 214066 107545
rect 214010 107471 214066 107480
rect 213918 106856 213974 106865
rect 213918 106791 213974 106800
rect 213932 106418 213960 106791
rect 213920 106412 213972 106418
rect 213920 106354 213972 106360
rect 214024 106350 214052 107471
rect 214012 106344 214064 106350
rect 214012 106286 214064 106292
rect 214010 106176 214066 106185
rect 214010 106111 214066 106120
rect 213918 105632 213974 105641
rect 213918 105567 213974 105576
rect 213932 104990 213960 105567
rect 213920 104984 213972 104990
rect 213920 104926 213972 104932
rect 214024 104922 214052 106111
rect 214012 104916 214064 104922
rect 214012 104858 214064 104864
rect 213918 102232 213974 102241
rect 213918 102167 213920 102176
rect 213972 102167 213974 102176
rect 213920 102138 213972 102144
rect 214010 101552 214066 101561
rect 214010 101487 214066 101496
rect 213918 101008 213974 101017
rect 213918 100943 213974 100952
rect 213932 100774 213960 100943
rect 214024 100842 214052 101487
rect 214012 100836 214064 100842
rect 214012 100778 214064 100784
rect 213920 100768 213972 100774
rect 213920 100710 213972 100716
rect 213918 99648 213974 99657
rect 213918 99583 213974 99592
rect 213932 99414 213960 99583
rect 213920 99408 213972 99414
rect 213920 99350 213972 99356
rect 214010 98968 214066 98977
rect 214010 98903 214066 98912
rect 213918 98288 213974 98297
rect 213918 98223 213974 98232
rect 213932 98122 213960 98223
rect 213920 98116 213972 98122
rect 213920 98058 213972 98064
rect 214024 98054 214052 98903
rect 214012 98048 214064 98054
rect 214012 97990 214064 97996
rect 213460 97300 213512 97306
rect 213460 97242 213512 97248
rect 213368 91792 213420 91798
rect 213368 91734 213420 91740
rect 213472 90438 213500 97242
rect 213918 96928 213974 96937
rect 213918 96863 213974 96872
rect 213932 96694 213960 96863
rect 213920 96688 213972 96694
rect 213920 96630 213972 96636
rect 213460 90432 213512 90438
rect 213460 90374 213512 90380
rect 214576 85542 214604 122806
rect 214760 113830 214788 126647
rect 215022 124672 215078 124681
rect 215022 124607 215078 124616
rect 214748 113824 214800 113830
rect 214748 113766 214800 113772
rect 215036 113174 215064 124607
rect 214668 113146 215064 113174
rect 214668 95946 214696 113146
rect 214746 104952 214802 104961
rect 214746 104887 214802 104896
rect 214656 95940 214708 95946
rect 214656 95882 214708 95888
rect 214564 85536 214616 85542
rect 214564 85478 214616 85484
rect 214656 80776 214708 80782
rect 214656 80718 214708 80724
rect 214564 79348 214616 79354
rect 214564 79290 214616 79296
rect 213276 56568 213328 56574
rect 213276 56510 213328 56516
rect 214576 15978 214604 79290
rect 214668 28422 214696 80718
rect 214760 75886 214788 104887
rect 214930 100328 214986 100337
rect 214930 100263 214986 100272
rect 214838 96384 214894 96393
rect 214838 96319 214894 96328
rect 214852 87718 214880 96319
rect 214944 93265 214972 100263
rect 215956 93945 215984 136575
rect 216126 133920 216182 133929
rect 216126 133855 216182 133864
rect 216034 95840 216090 95849
rect 216034 95775 216090 95784
rect 215942 93936 215998 93945
rect 215942 93871 215998 93880
rect 214930 93256 214986 93265
rect 216048 93226 216076 95775
rect 214930 93191 214986 93200
rect 216036 93220 216088 93226
rect 216036 93162 216088 93168
rect 215942 90400 215998 90409
rect 215942 90335 215998 90344
rect 214840 87712 214892 87718
rect 214840 87654 214892 87660
rect 214748 75880 214800 75886
rect 214748 75822 214800 75828
rect 214656 28416 214708 28422
rect 214656 28358 214708 28364
rect 215956 20058 215984 90335
rect 216140 89010 216168 133855
rect 216310 100056 216366 100065
rect 216310 99991 216366 100000
rect 217232 100020 217284 100026
rect 216220 94580 216272 94586
rect 216220 94522 216272 94528
rect 216128 89004 216180 89010
rect 216128 88946 216180 88952
rect 216232 84194 216260 94522
rect 216324 88262 216352 99991
rect 217232 99962 217284 99968
rect 216678 98696 216734 98705
rect 216678 98631 216734 98640
rect 216692 94518 216720 98631
rect 216680 94512 216732 94518
rect 216680 94454 216732 94460
rect 217244 92478 217272 99962
rect 219164 96076 219216 96082
rect 219164 96018 219216 96024
rect 219176 95985 219204 96018
rect 225604 96008 225656 96014
rect 219162 95976 219218 95985
rect 225604 95950 225656 95956
rect 219162 95911 219218 95920
rect 223488 94512 223540 94518
rect 223488 94454 223540 94460
rect 220084 93152 220136 93158
rect 220084 93094 220136 93100
rect 217232 92472 217284 92478
rect 217232 92414 217284 92420
rect 218704 90432 218756 90438
rect 218704 90374 218756 90380
rect 216312 88256 216364 88262
rect 216312 88198 216364 88204
rect 216048 84166 216260 84194
rect 216048 25566 216076 84166
rect 217324 82204 217376 82210
rect 217324 82146 217376 82152
rect 217336 47598 217364 82146
rect 217324 47592 217376 47598
rect 217324 47534 217376 47540
rect 216036 25560 216088 25566
rect 216036 25502 216088 25508
rect 215944 20052 215996 20058
rect 215944 19994 215996 20000
rect 214564 15972 214616 15978
rect 214564 15914 214616 15920
rect 218716 14482 218744 90374
rect 218704 14476 218756 14482
rect 218704 14418 218756 14424
rect 220096 3466 220124 93094
rect 223500 91050 223528 94454
rect 224314 93936 224370 93945
rect 224314 93871 224370 93880
rect 223488 91044 223540 91050
rect 223488 90986 223540 90992
rect 223028 90364 223080 90370
rect 223028 90306 223080 90312
rect 221464 89004 221516 89010
rect 221464 88946 221516 88952
rect 220176 83496 220228 83502
rect 220176 83438 220228 83444
rect 220188 57322 220216 83438
rect 220176 57316 220228 57322
rect 220176 57258 220228 57264
rect 221476 35290 221504 88946
rect 222844 86284 222896 86290
rect 222844 86226 222896 86232
rect 221464 35284 221516 35290
rect 221464 35226 221516 35232
rect 222856 18698 222884 86226
rect 222936 83496 222988 83502
rect 222936 83438 222988 83444
rect 222948 37942 222976 83438
rect 223040 82113 223068 90306
rect 224224 89072 224276 89078
rect 224224 89014 224276 89020
rect 223026 82104 223082 82113
rect 223026 82039 223082 82048
rect 222936 37936 222988 37942
rect 222936 37878 222988 37884
rect 222844 18692 222896 18698
rect 222844 18634 222896 18640
rect 224236 13122 224264 89014
rect 224328 35222 224356 93871
rect 225616 86902 225644 95950
rect 227076 95940 227128 95946
rect 227076 95882 227128 95888
rect 226984 94512 227036 94518
rect 226984 94454 227036 94460
rect 225604 86896 225656 86902
rect 225604 86838 225656 86844
rect 224316 35216 224368 35222
rect 224316 35158 224368 35164
rect 226996 33862 227024 94454
rect 227088 53174 227116 95882
rect 228454 95296 228510 95305
rect 228454 95231 228510 95240
rect 228362 87544 228418 87553
rect 228362 87479 228418 87488
rect 227076 53168 227128 53174
rect 227076 53110 227128 53116
rect 227076 47660 227128 47666
rect 227076 47602 227128 47608
rect 226984 33856 227036 33862
rect 226984 33798 227036 33804
rect 224224 13116 224276 13122
rect 224224 13058 224276 13064
rect 227088 11762 227116 47602
rect 228376 39370 228404 87479
rect 228468 79529 228496 95231
rect 228454 79520 228510 79529
rect 228454 79455 228510 79464
rect 229756 72554 229784 136614
rect 229848 117065 229876 157791
rect 230584 155281 230612 159394
rect 230676 157729 230704 192442
rect 231124 184204 231176 184210
rect 231124 184146 231176 184152
rect 230848 179444 230900 179450
rect 230848 179386 230900 179392
rect 230756 170672 230808 170678
rect 230756 170614 230808 170620
rect 230768 170513 230796 170614
rect 230754 170504 230810 170513
rect 230754 170439 230810 170448
rect 230860 169969 230888 179386
rect 231136 176730 231164 184146
rect 231780 178265 231808 237351
rect 231952 234660 232004 234666
rect 231952 234602 232004 234608
rect 231860 234592 231912 234598
rect 231860 234534 231912 234540
rect 231872 234161 231900 234534
rect 231858 234152 231914 234161
rect 231858 234087 231914 234096
rect 231964 217433 231992 234602
rect 231950 217424 232006 217433
rect 231950 217359 232006 217368
rect 232516 214441 232544 240071
rect 232608 240038 232636 240244
rect 232596 240032 232648 240038
rect 232596 239974 232648 239980
rect 232976 238754 233004 240244
rect 232976 238726 233096 238754
rect 232964 238060 233016 238066
rect 232964 238002 233016 238008
rect 232976 232626 233004 238002
rect 232964 232620 233016 232626
rect 232964 232562 233016 232568
rect 233068 230450 233096 238726
rect 233332 234728 233384 234734
rect 233528 234705 233556 240244
rect 234080 238785 234108 240244
rect 234066 238776 234122 238785
rect 234066 238711 234122 238720
rect 233332 234670 233384 234676
rect 233514 234696 233570 234705
rect 233056 230444 233108 230450
rect 233056 230386 233108 230392
rect 232502 214432 232558 214441
rect 232502 214367 232558 214376
rect 231952 213988 232004 213994
rect 231952 213930 232004 213936
rect 231766 178256 231822 178265
rect 231766 178191 231822 178200
rect 231124 176724 231176 176730
rect 231124 176666 231176 176672
rect 231860 176724 231912 176730
rect 231860 176666 231912 176672
rect 230940 174004 230992 174010
rect 230940 173946 230992 173952
rect 230846 169960 230902 169969
rect 230846 169895 230902 169904
rect 230952 168609 230980 173946
rect 231676 173188 231728 173194
rect 231676 173130 231728 173136
rect 231400 172508 231452 172514
rect 231400 172450 231452 172456
rect 231412 171873 231440 172450
rect 231688 172417 231716 173130
rect 231768 172440 231820 172446
rect 231674 172408 231730 172417
rect 231768 172382 231820 172388
rect 231674 172343 231730 172352
rect 231398 171864 231454 171873
rect 231398 171799 231454 171808
rect 231780 171465 231808 172382
rect 231766 171456 231822 171465
rect 231766 171391 231822 171400
rect 231124 170400 231176 170406
rect 231124 170342 231176 170348
rect 231674 170368 231730 170377
rect 230938 168600 230994 168609
rect 230938 168535 230994 168544
rect 230940 165164 230992 165170
rect 230940 165106 230992 165112
rect 230952 164393 230980 165106
rect 230938 164384 230994 164393
rect 230938 164319 230994 164328
rect 231032 164212 231084 164218
rect 231032 164154 231084 164160
rect 231044 163849 231072 164154
rect 231030 163840 231086 163849
rect 231030 163775 231086 163784
rect 231136 162897 231164 170342
rect 231674 170303 231730 170312
rect 231492 168360 231544 168366
rect 231492 168302 231544 168308
rect 231504 167657 231532 168302
rect 231490 167648 231546 167657
rect 231490 167583 231546 167592
rect 231308 166932 231360 166938
rect 231308 166874 231360 166880
rect 231320 166161 231348 166874
rect 231306 166152 231362 166161
rect 231306 166087 231362 166096
rect 231492 165232 231544 165238
rect 231490 165200 231492 165209
rect 231544 165200 231546 165209
rect 231490 165135 231546 165144
rect 231398 165064 231454 165073
rect 231398 164999 231454 165008
rect 231122 162888 231178 162897
rect 231122 162823 231178 162832
rect 231032 161084 231084 161090
rect 231032 161026 231084 161032
rect 231044 160585 231072 161026
rect 231030 160576 231086 160585
rect 231030 160511 231086 160520
rect 230662 157720 230718 157729
rect 230662 157655 230718 157664
rect 231214 156632 231270 156641
rect 231214 156567 231270 156576
rect 230570 155272 230626 155281
rect 230570 155207 230626 155216
rect 231228 154873 231256 156567
rect 231214 154864 231270 154873
rect 231214 154799 231270 154808
rect 231306 154456 231362 154465
rect 231306 154391 231362 154400
rect 230664 153876 230716 153882
rect 230664 153818 230716 153824
rect 230570 153096 230626 153105
rect 230570 153031 230626 153040
rect 230480 152516 230532 152522
rect 230480 152458 230532 152464
rect 230492 151858 230520 152458
rect 230584 152017 230612 153031
rect 230570 152008 230626 152017
rect 230570 151943 230626 151952
rect 230492 151830 230612 151858
rect 230480 151632 230532 151638
rect 230478 151600 230480 151609
rect 230532 151600 230534 151609
rect 230478 151535 230534 151544
rect 229928 151088 229980 151094
rect 229928 151030 229980 151036
rect 229834 117056 229890 117065
rect 229834 116991 229890 117000
rect 229834 114880 229890 114889
rect 229834 114815 229890 114824
rect 229744 72548 229796 72554
rect 229744 72490 229796 72496
rect 229848 57225 229876 114815
rect 229940 113257 229968 151030
rect 230584 147801 230612 151830
rect 230676 151065 230704 153818
rect 231216 153740 231268 153746
rect 231216 153682 231268 153688
rect 231228 153377 231256 153682
rect 231214 153368 231270 153377
rect 231214 153303 231270 153312
rect 230662 151056 230718 151065
rect 230662 150991 230718 151000
rect 231124 148368 231176 148374
rect 231124 148310 231176 148316
rect 230570 147792 230626 147801
rect 230570 147727 230626 147736
rect 230570 146296 230626 146305
rect 230570 146231 230626 146240
rect 230584 140185 230612 146231
rect 230570 140176 230626 140185
rect 230570 140111 230626 140120
rect 230756 135108 230808 135114
rect 230756 135050 230808 135056
rect 230768 126041 230796 135050
rect 231136 131209 231164 148310
rect 231320 142154 231348 154391
rect 231412 153921 231440 164999
rect 231688 164801 231716 170303
rect 231768 169584 231820 169590
rect 231766 169552 231768 169561
rect 231820 169552 231822 169561
rect 231766 169487 231822 169496
rect 231768 169176 231820 169182
rect 231768 169118 231820 169124
rect 231780 169017 231808 169118
rect 231766 169008 231822 169017
rect 231766 168943 231822 168952
rect 231766 168056 231822 168065
rect 231872 168042 231900 176666
rect 231822 168014 231900 168042
rect 231766 167991 231822 168000
rect 231768 166728 231820 166734
rect 231766 166696 231768 166705
rect 231820 166696 231822 166705
rect 231766 166631 231822 166640
rect 231674 164792 231730 164801
rect 231674 164727 231730 164736
rect 231676 162784 231728 162790
rect 231676 162726 231728 162732
rect 231688 161537 231716 162726
rect 231674 161528 231730 161537
rect 231674 161463 231730 161472
rect 231766 160712 231822 160721
rect 231766 160647 231822 160656
rect 231780 160041 231808 160647
rect 231964 160138 231992 213930
rect 232134 206816 232190 206825
rect 232134 206751 232190 206760
rect 232044 182912 232096 182918
rect 232044 182854 232096 182860
rect 231952 160132 232004 160138
rect 231952 160074 232004 160080
rect 231766 160032 231822 160041
rect 231766 159967 231822 159976
rect 231768 158704 231820 158710
rect 231766 158672 231768 158681
rect 231820 158672 231822 158681
rect 231492 158636 231544 158642
rect 231766 158607 231822 158616
rect 231492 158578 231544 158584
rect 231504 158137 231532 158578
rect 231490 158128 231546 158137
rect 231490 158063 231546 158072
rect 231674 157992 231730 158001
rect 231674 157927 231730 157936
rect 231688 157185 231716 157927
rect 231768 157344 231820 157350
rect 231768 157286 231820 157292
rect 231674 157176 231730 157185
rect 231674 157111 231730 157120
rect 231780 156777 231808 157286
rect 231766 156768 231822 156777
rect 231766 156703 231822 156712
rect 231768 155916 231820 155922
rect 231768 155858 231820 155864
rect 231780 155825 231808 155858
rect 231766 155816 231822 155825
rect 231766 155751 231822 155760
rect 231766 155272 231822 155281
rect 231766 155207 231822 155216
rect 231780 154329 231808 155207
rect 231766 154320 231822 154329
rect 231766 154255 231822 154264
rect 231398 153912 231454 153921
rect 231398 153847 231454 153856
rect 231766 153912 231822 153921
rect 231766 153847 231822 153856
rect 231780 152969 231808 153847
rect 231766 152960 231822 152969
rect 231766 152895 231822 152904
rect 232056 151814 232084 182854
rect 231872 151786 232084 151814
rect 231674 151056 231730 151065
rect 231674 150991 231730 151000
rect 231490 148336 231546 148345
rect 231490 148271 231546 148280
rect 231504 144945 231532 148271
rect 231490 144936 231546 144945
rect 231490 144871 231546 144880
rect 231688 143449 231716 150991
rect 231872 147098 231900 151786
rect 232148 151638 232176 206751
rect 233240 175976 233292 175982
rect 233240 175918 233292 175924
rect 233252 170678 233280 175918
rect 233240 170672 233292 170678
rect 233240 170614 233292 170620
rect 233344 165170 233372 234670
rect 233514 234631 233570 234640
rect 233528 231305 233556 234631
rect 233514 231296 233570 231305
rect 233514 231231 233570 231240
rect 233424 230444 233476 230450
rect 233424 230386 233476 230392
rect 233436 229770 233464 230386
rect 233424 229764 233476 229770
rect 233424 229706 233476 229712
rect 233436 220833 233464 229706
rect 234080 226273 234108 238711
rect 234066 226264 234122 226273
rect 234066 226199 234122 226208
rect 233422 220824 233478 220833
rect 233422 220759 233478 220768
rect 233516 216640 233568 216646
rect 233516 216582 233568 216588
rect 233528 216102 233556 216582
rect 234448 216102 234476 240244
rect 235000 231713 235028 240244
rect 234986 231704 235042 231713
rect 234986 231639 235042 231648
rect 235368 222193 235396 240244
rect 235354 222184 235410 222193
rect 235354 222119 235410 222128
rect 235368 217326 235396 222119
rect 235356 217320 235408 217326
rect 235356 217262 235408 217268
rect 233516 216096 233568 216102
rect 233516 216038 233568 216044
rect 234436 216096 234488 216102
rect 234436 216038 234488 216044
rect 233424 188420 233476 188426
rect 233424 188362 233476 188368
rect 233332 165164 233384 165170
rect 233332 165106 233384 165112
rect 232502 164928 232558 164937
rect 232502 164863 232558 164872
rect 232136 151632 232188 151638
rect 232136 151574 232188 151580
rect 231780 147070 231900 147098
rect 231780 146849 231808 147070
rect 231860 146940 231912 146946
rect 231860 146882 231912 146888
rect 231766 146840 231822 146849
rect 231766 146775 231822 146784
rect 231766 146160 231822 146169
rect 231872 146146 231900 146882
rect 231822 146118 231900 146146
rect 231766 146095 231822 146104
rect 231768 144900 231820 144906
rect 231768 144842 231820 144848
rect 231780 143993 231808 144842
rect 231766 143984 231822 143993
rect 231766 143919 231822 143928
rect 231674 143440 231730 143449
rect 231674 143375 231730 143384
rect 231768 142860 231820 142866
rect 231768 142802 231820 142808
rect 231780 142497 231808 142802
rect 231766 142488 231822 142497
rect 231766 142423 231822 142432
rect 231228 142126 231348 142154
rect 231228 141681 231256 142126
rect 231214 141672 231270 141681
rect 231214 141607 231270 141616
rect 231216 139528 231268 139534
rect 231216 139470 231268 139476
rect 231228 133113 231256 139470
rect 231400 139460 231452 139466
rect 231400 139402 231452 139408
rect 231308 138848 231360 138854
rect 231308 138790 231360 138796
rect 231320 135969 231348 138790
rect 231306 135960 231362 135969
rect 231306 135895 231362 135904
rect 231214 133104 231270 133113
rect 231214 133039 231270 133048
rect 231412 132494 231440 139402
rect 231768 139392 231820 139398
rect 231768 139334 231820 139340
rect 231780 138281 231808 139334
rect 231766 138272 231822 138281
rect 231766 138207 231822 138216
rect 231584 137964 231636 137970
rect 231584 137906 231636 137912
rect 231596 136921 231624 137906
rect 231582 136912 231638 136921
rect 231582 136847 231638 136856
rect 231492 136604 231544 136610
rect 231492 136546 231544 136552
rect 231504 135425 231532 136546
rect 231768 136536 231820 136542
rect 231768 136478 231820 136484
rect 231780 136377 231808 136478
rect 231766 136368 231822 136377
rect 231766 136303 231822 136312
rect 231490 135416 231546 135425
rect 231490 135351 231546 135360
rect 231492 135244 231544 135250
rect 231492 135186 231544 135192
rect 231504 134065 231532 135186
rect 231766 135144 231822 135153
rect 231766 135079 231822 135088
rect 231780 134473 231808 135079
rect 231766 134464 231822 134473
rect 231766 134399 231822 134408
rect 231490 134056 231546 134065
rect 231490 133991 231546 134000
rect 231676 133884 231728 133890
rect 231676 133826 231728 133832
rect 231688 132569 231716 133826
rect 231768 133816 231820 133822
rect 231768 133758 231820 133764
rect 231780 133521 231808 133758
rect 231766 133512 231822 133521
rect 231766 133447 231822 133456
rect 231674 132560 231730 132569
rect 231674 132495 231730 132504
rect 231320 132466 231440 132494
rect 231122 131200 231178 131209
rect 231122 131135 231178 131144
rect 231320 129849 231348 132466
rect 231768 132456 231820 132462
rect 231768 132398 231820 132404
rect 231676 131776 231728 131782
rect 231676 131718 231728 131724
rect 231400 131028 231452 131034
rect 231400 130970 231452 130976
rect 231412 130257 231440 130970
rect 231398 130248 231454 130257
rect 231398 130183 231454 130192
rect 231306 129840 231362 129849
rect 231306 129775 231362 129784
rect 231490 129840 231546 129849
rect 231490 129775 231546 129784
rect 231400 129668 231452 129674
rect 231400 129610 231452 129616
rect 231412 128897 231440 129610
rect 231398 128888 231454 128897
rect 231398 128823 231454 128832
rect 231308 128036 231360 128042
rect 231308 127978 231360 127984
rect 231320 127401 231348 127978
rect 231306 127392 231362 127401
rect 231306 127327 231362 127336
rect 230754 126032 230810 126041
rect 230754 125967 230810 125976
rect 230756 124976 230808 124982
rect 230756 124918 230808 124924
rect 230664 124908 230716 124914
rect 230664 124850 230716 124856
rect 230572 124092 230624 124098
rect 230572 124034 230624 124040
rect 230584 123593 230612 124034
rect 230570 123584 230626 123593
rect 230570 123519 230626 123528
rect 230018 122088 230074 122097
rect 230018 122023 230074 122032
rect 229926 113248 229982 113257
rect 229926 113183 229982 113192
rect 230032 89049 230060 122023
rect 230676 120329 230704 124850
rect 230662 120320 230718 120329
rect 230662 120255 230718 120264
rect 230768 116113 230796 124918
rect 231214 123448 231270 123457
rect 231214 123383 231270 123392
rect 230940 121916 230992 121922
rect 230940 121858 230992 121864
rect 230952 121689 230980 121858
rect 230938 121680 230994 121689
rect 230938 121615 230994 121624
rect 231122 120184 231178 120193
rect 231122 120119 231178 120128
rect 231032 119944 231084 119950
rect 231032 119886 231084 119892
rect 230940 118448 230992 118454
rect 230940 118390 230992 118396
rect 230952 118017 230980 118390
rect 230938 118008 230994 118017
rect 230938 117943 230994 117952
rect 231044 117473 231072 119886
rect 231030 117464 231086 117473
rect 231030 117399 231086 117408
rect 230754 116104 230810 116113
rect 230754 116039 230810 116048
rect 230664 114980 230716 114986
rect 230664 114922 230716 114928
rect 230676 114617 230704 114922
rect 230662 114608 230718 114617
rect 230662 114543 230718 114552
rect 230940 113076 230992 113082
rect 230940 113018 230992 113024
rect 230952 112713 230980 113018
rect 230938 112704 230994 112713
rect 230938 112639 230994 112648
rect 230756 110900 230808 110906
rect 230756 110842 230808 110848
rect 230768 110809 230796 110842
rect 230754 110800 230810 110809
rect 230754 110735 230810 110744
rect 230756 103488 230808 103494
rect 230756 103430 230808 103436
rect 230768 102377 230796 103430
rect 231136 103329 231164 120119
rect 231228 105233 231256 123383
rect 231504 122834 231532 129775
rect 231688 127945 231716 131718
rect 231780 131617 231808 132398
rect 231766 131608 231822 131617
rect 231766 131543 231822 131552
rect 231768 131096 231820 131102
rect 231768 131038 231820 131044
rect 231780 130665 231808 131038
rect 231766 130656 231822 130665
rect 231766 130591 231822 130600
rect 231768 129736 231820 129742
rect 231768 129678 231820 129684
rect 231780 129305 231808 129678
rect 231766 129296 231822 129305
rect 231766 129231 231822 129240
rect 231766 128344 231822 128353
rect 231766 128279 231768 128288
rect 231820 128279 231822 128288
rect 231768 128250 231820 128256
rect 231674 127936 231730 127945
rect 231674 127871 231730 127880
rect 231582 127664 231638 127673
rect 231582 127599 231638 127608
rect 231596 124137 231624 127599
rect 231766 126984 231822 126993
rect 231676 126948 231728 126954
rect 231766 126919 231822 126928
rect 231676 126890 231728 126896
rect 231688 126449 231716 126890
rect 231780 126886 231808 126919
rect 231768 126880 231820 126886
rect 231768 126822 231820 126828
rect 231674 126440 231730 126449
rect 231674 126375 231730 126384
rect 232516 125497 232544 164863
rect 232688 159384 232740 159390
rect 232688 159326 232740 159332
rect 232596 141432 232648 141438
rect 232596 141374 232648 141380
rect 232502 125488 232558 125497
rect 232502 125423 232558 125432
rect 231766 125352 231822 125361
rect 231766 125287 231822 125296
rect 231780 124545 231808 125287
rect 231766 124536 231822 124545
rect 231766 124471 231822 124480
rect 231768 124160 231820 124166
rect 231582 124128 231638 124137
rect 231768 124102 231820 124108
rect 231582 124063 231638 124072
rect 231780 123185 231808 124102
rect 231766 123176 231822 123185
rect 231766 123111 231822 123120
rect 231320 122806 231532 122834
rect 231320 119377 231348 122806
rect 231768 122800 231820 122806
rect 231768 122742 231820 122748
rect 231780 122233 231808 122742
rect 231766 122224 231822 122233
rect 231766 122159 231822 122168
rect 231676 121440 231728 121446
rect 231676 121382 231728 121388
rect 231688 120737 231716 121382
rect 231768 121372 231820 121378
rect 231768 121314 231820 121320
rect 231780 121281 231808 121314
rect 231766 121272 231822 121281
rect 231766 121207 231822 121216
rect 231674 120728 231730 120737
rect 231674 120663 231730 120672
rect 232502 120456 232558 120465
rect 232502 120391 232558 120400
rect 231768 120080 231820 120086
rect 231768 120022 231820 120028
rect 231306 119368 231362 119377
rect 231306 119303 231362 119312
rect 231780 118969 231808 120022
rect 231766 118960 231822 118969
rect 231766 118895 231822 118904
rect 231768 118652 231820 118658
rect 231768 118594 231820 118600
rect 231780 118425 231808 118594
rect 231766 118416 231822 118425
rect 231766 118351 231822 118360
rect 231582 118008 231638 118017
rect 231582 117943 231638 117952
rect 231492 117292 231544 117298
rect 231492 117234 231544 117240
rect 231504 116521 231532 117234
rect 231490 116512 231546 116521
rect 231490 116447 231546 116456
rect 231492 115932 231544 115938
rect 231492 115874 231544 115880
rect 231504 115161 231532 115874
rect 231490 115152 231546 115161
rect 231490 115087 231546 115096
rect 231398 113792 231454 113801
rect 231398 113727 231454 113736
rect 231308 108928 231360 108934
rect 231308 108870 231360 108876
rect 231320 107953 231348 108870
rect 231306 107944 231362 107953
rect 231306 107879 231362 107888
rect 231308 106276 231360 106282
rect 231308 106218 231360 106224
rect 231320 105641 231348 106218
rect 231306 105632 231362 105641
rect 231306 105567 231362 105576
rect 231214 105224 231270 105233
rect 231214 105159 231270 105168
rect 231216 105120 231268 105126
rect 231216 105062 231268 105068
rect 231122 103320 231178 103329
rect 231122 103255 231178 103264
rect 230754 102368 230810 102377
rect 230754 102303 230810 102312
rect 230572 101924 230624 101930
rect 230572 101866 230624 101872
rect 230584 101833 230612 101866
rect 230570 101824 230626 101833
rect 230570 101759 230626 101768
rect 230938 100736 230994 100745
rect 230938 100671 230994 100680
rect 230952 99521 230980 100671
rect 230938 99512 230994 99521
rect 230938 99447 230994 99456
rect 231122 98696 231178 98705
rect 231122 98631 231178 98640
rect 230570 96656 230626 96665
rect 230570 96591 230626 96600
rect 230478 96248 230534 96257
rect 230478 96183 230534 96192
rect 230492 96082 230520 96183
rect 230480 96076 230532 96082
rect 230480 96018 230532 96024
rect 230018 89040 230074 89049
rect 230018 88975 230074 88984
rect 230584 84194 230612 96591
rect 230492 84166 230612 84194
rect 229834 57216 229890 57225
rect 229834 57151 229890 57160
rect 230492 42158 230520 84166
rect 231136 53106 231164 98631
rect 231228 94489 231256 105062
rect 231308 102876 231360 102882
rect 231308 102818 231360 102824
rect 231320 102785 231348 102818
rect 231306 102776 231362 102785
rect 231306 102711 231362 102720
rect 231306 102232 231362 102241
rect 231306 102167 231362 102176
rect 231320 98569 231348 102167
rect 231412 101425 231440 113727
rect 231596 111761 231624 117943
rect 231768 114504 231820 114510
rect 231768 114446 231820 114452
rect 231676 114436 231728 114442
rect 231676 114378 231728 114384
rect 231688 113665 231716 114378
rect 231780 114209 231808 114446
rect 231766 114200 231822 114209
rect 231766 114135 231822 114144
rect 231674 113656 231730 113665
rect 231674 113591 231730 113600
rect 231768 113144 231820 113150
rect 231768 113086 231820 113092
rect 231780 112305 231808 113086
rect 231766 112296 231822 112305
rect 231766 112231 231822 112240
rect 231768 111784 231820 111790
rect 231582 111752 231638 111761
rect 231768 111726 231820 111732
rect 231582 111687 231638 111696
rect 231780 111353 231808 111726
rect 231766 111344 231822 111353
rect 231766 111279 231822 111288
rect 231490 111072 231546 111081
rect 231490 111007 231546 111016
rect 231504 105126 231532 111007
rect 231676 110424 231728 110430
rect 231676 110366 231728 110372
rect 231688 109857 231716 110366
rect 231768 110356 231820 110362
rect 231768 110298 231820 110304
rect 231674 109848 231730 109857
rect 231674 109783 231730 109792
rect 231780 109449 231808 110298
rect 231766 109440 231822 109449
rect 231766 109375 231822 109384
rect 231768 108996 231820 109002
rect 231768 108938 231820 108944
rect 231780 108497 231808 108938
rect 231766 108488 231822 108497
rect 231766 108423 231822 108432
rect 231768 107636 231820 107642
rect 231768 107578 231820 107584
rect 231676 107568 231728 107574
rect 231676 107510 231728 107516
rect 231688 106593 231716 107510
rect 231780 107137 231808 107578
rect 231766 107128 231822 107137
rect 231766 107063 231822 107072
rect 231674 106584 231730 106593
rect 231674 106519 231730 106528
rect 231584 106208 231636 106214
rect 231582 106176 231584 106185
rect 231636 106176 231638 106185
rect 231582 106111 231638 106120
rect 231492 105120 231544 105126
rect 231492 105062 231544 105068
rect 231768 104848 231820 104854
rect 231768 104790 231820 104796
rect 231676 104712 231728 104718
rect 231674 104680 231676 104689
rect 231728 104680 231730 104689
rect 231674 104615 231730 104624
rect 231780 103737 231808 104790
rect 231766 103728 231822 103737
rect 231766 103663 231822 103672
rect 231584 102060 231636 102066
rect 231584 102002 231636 102008
rect 231490 101552 231546 101561
rect 231490 101487 231546 101496
rect 231398 101416 231454 101425
rect 231398 101351 231454 101360
rect 231306 98560 231362 98569
rect 231306 98495 231362 98504
rect 231504 97617 231532 101487
rect 231596 100881 231624 102002
rect 231582 100872 231638 100881
rect 231582 100807 231638 100816
rect 231676 100700 231728 100706
rect 231676 100642 231728 100648
rect 231688 99929 231716 100642
rect 231768 100632 231820 100638
rect 231768 100574 231820 100580
rect 231780 100473 231808 100574
rect 231766 100464 231822 100473
rect 231766 100399 231822 100408
rect 231674 99920 231730 99929
rect 231674 99855 231730 99864
rect 231676 99340 231728 99346
rect 231676 99282 231728 99288
rect 231688 98025 231716 99282
rect 231768 99272 231820 99278
rect 231768 99214 231820 99220
rect 231780 98977 231808 99214
rect 231766 98968 231822 98977
rect 231766 98903 231822 98912
rect 231674 98016 231730 98025
rect 231674 97951 231730 97960
rect 231490 97608 231546 97617
rect 231490 97543 231546 97552
rect 231766 97064 231822 97073
rect 231766 96999 231822 97008
rect 231676 96688 231728 96694
rect 231674 96656 231676 96665
rect 231728 96656 231730 96665
rect 231674 96591 231730 96600
rect 231780 96529 231808 96999
rect 231766 96520 231822 96529
rect 231766 96455 231822 96464
rect 231214 94480 231270 94489
rect 231214 94415 231270 94424
rect 231124 53100 231176 53106
rect 231124 53042 231176 53048
rect 230480 42152 230532 42158
rect 230480 42094 230532 42100
rect 228364 39364 228416 39370
rect 228364 39306 228416 39312
rect 232516 26994 232544 120391
rect 232608 101930 232636 141374
rect 232700 124098 232728 159326
rect 233436 153746 233464 188362
rect 233528 161090 233556 216038
rect 235264 207732 235316 207738
rect 235264 207674 235316 207680
rect 234712 180124 234764 180130
rect 234712 180066 234764 180072
rect 234620 177336 234672 177342
rect 234620 177278 234672 177284
rect 233976 167068 234028 167074
rect 233976 167010 234028 167016
rect 233516 161084 233568 161090
rect 233516 161026 233568 161032
rect 233884 154624 233936 154630
rect 233884 154566 233936 154572
rect 233424 153740 233476 153746
rect 233424 153682 233476 153688
rect 232872 144968 232924 144974
rect 232872 144910 232924 144916
rect 232688 124092 232740 124098
rect 232688 124034 232740 124040
rect 232780 123480 232832 123486
rect 232780 123422 232832 123428
rect 232686 112160 232742 112169
rect 232686 112095 232742 112104
rect 232596 101924 232648 101930
rect 232596 101866 232648 101872
rect 232596 96076 232648 96082
rect 232596 96018 232648 96024
rect 232504 26988 232556 26994
rect 232504 26930 232556 26936
rect 227076 11756 227128 11762
rect 227076 11698 227128 11704
rect 232608 4214 232636 96018
rect 232700 82249 232728 112095
rect 232792 94586 232820 123422
rect 232884 120193 232912 144910
rect 232870 120184 232926 120193
rect 232870 120119 232926 120128
rect 233896 114986 233924 154566
rect 233988 128042 234016 167010
rect 234632 166938 234660 177278
rect 234724 169182 234752 180066
rect 235276 177342 235304 207674
rect 235920 206961 235948 240244
rect 236366 240000 236422 240009
rect 236366 239935 236422 239944
rect 236380 238754 236408 239935
rect 236472 239442 236500 240244
rect 236472 239414 236592 239442
rect 236380 238726 236500 238754
rect 236472 235657 236500 238726
rect 236564 235793 236592 239414
rect 236840 237522 236868 240244
rect 237392 238754 237420 240244
rect 237470 240136 237526 240145
rect 237470 240071 237526 240080
rect 237484 240038 237512 240071
rect 237472 240032 237524 240038
rect 237472 239974 237524 239980
rect 237392 238726 237512 238754
rect 237484 237590 237512 238726
rect 237472 237584 237524 237590
rect 237472 237526 237524 237532
rect 236828 237516 236880 237522
rect 236828 237458 236880 237464
rect 236644 236700 236696 236706
rect 236644 236642 236696 236648
rect 236550 235784 236606 235793
rect 236550 235719 236606 235728
rect 236458 235648 236514 235657
rect 236458 235583 236514 235592
rect 235906 206952 235962 206961
rect 235906 206887 235962 206896
rect 236000 200864 236052 200870
rect 236000 200806 236052 200812
rect 235356 186992 235408 186998
rect 235356 186934 235408 186940
rect 235264 177336 235316 177342
rect 235264 177278 235316 177284
rect 234804 176044 234856 176050
rect 234804 175986 234856 175992
rect 234712 169176 234764 169182
rect 234712 169118 234764 169124
rect 234816 168366 234844 175986
rect 235368 170513 235396 186934
rect 235354 170504 235410 170513
rect 235354 170439 235410 170448
rect 236012 169590 236040 200806
rect 236090 177576 236146 177585
rect 236090 177511 236146 177520
rect 236000 169584 236052 169590
rect 236000 169526 236052 169532
rect 235264 168428 235316 168434
rect 235264 168370 235316 168376
rect 234804 168360 234856 168366
rect 234804 168302 234856 168308
rect 234712 168020 234764 168026
rect 234712 167962 234764 167968
rect 234620 166932 234672 166938
rect 234620 166874 234672 166880
rect 234618 166832 234674 166841
rect 234618 166767 234674 166776
rect 234632 165238 234660 166767
rect 234724 166734 234752 167962
rect 234712 166728 234764 166734
rect 234712 166670 234764 166676
rect 234620 165232 234672 165238
rect 234620 165174 234672 165180
rect 234250 163432 234306 163441
rect 234250 163367 234306 163376
rect 234158 160440 234214 160449
rect 234158 160375 234214 160384
rect 234068 147688 234120 147694
rect 234068 147630 234120 147636
rect 233976 128036 234028 128042
rect 233976 127978 234028 127984
rect 233974 119096 234030 119105
rect 233974 119031 234030 119040
rect 233884 114980 233936 114986
rect 233884 114922 233936 114928
rect 233882 105224 233938 105233
rect 233882 105159 233938 105168
rect 232780 94580 232832 94586
rect 232780 94522 232832 94528
rect 232686 82240 232742 82249
rect 232686 82175 232742 82184
rect 233896 6186 233924 105159
rect 233988 76673 234016 119031
rect 234080 106214 234108 147630
rect 234172 119785 234200 160375
rect 234264 158642 234292 163367
rect 234252 158636 234304 158642
rect 234252 158578 234304 158584
rect 235276 139466 235304 168370
rect 235540 161492 235592 161498
rect 235540 161434 235592 161440
rect 235448 149116 235500 149122
rect 235448 149058 235500 149064
rect 235356 145036 235408 145042
rect 235356 144978 235408 144984
rect 235264 139460 235316 139466
rect 235264 139402 235316 139408
rect 235262 137048 235318 137057
rect 235262 136983 235318 136992
rect 234158 119776 234214 119785
rect 234158 119711 234214 119720
rect 234068 106208 234120 106214
rect 234068 106150 234120 106156
rect 233974 76664 234030 76673
rect 233974 76599 234030 76608
rect 235276 24138 235304 136983
rect 235368 102882 235396 144978
rect 235460 108934 235488 149058
rect 235552 121922 235580 161434
rect 236104 160993 236132 177511
rect 236090 160984 236146 160993
rect 236090 160919 236146 160928
rect 236656 146985 236684 236642
rect 237944 235521 237972 240244
rect 238024 237516 238076 237522
rect 238024 237458 238076 237464
rect 237378 235512 237434 235521
rect 237378 235447 237434 235456
rect 237930 235512 237986 235521
rect 237930 235447 237986 235456
rect 236920 172576 236972 172582
rect 236920 172518 236972 172524
rect 236734 156632 236790 156641
rect 236734 156567 236790 156576
rect 236642 146976 236698 146985
rect 236642 146911 236698 146920
rect 236642 138408 236698 138417
rect 236642 138343 236698 138352
rect 235540 121916 235592 121922
rect 235540 121858 235592 121864
rect 235540 116612 235592 116618
rect 235540 116554 235592 116560
rect 235448 108928 235500 108934
rect 235448 108870 235500 108876
rect 235356 102876 235408 102882
rect 235356 102818 235408 102824
rect 235552 80714 235580 116554
rect 235540 80708 235592 80714
rect 235540 80650 235592 80656
rect 236656 49026 236684 138343
rect 236748 118454 236776 156567
rect 236826 146704 236882 146713
rect 236826 146639 236882 146648
rect 236736 118448 236788 118454
rect 236736 118390 236788 118396
rect 236736 105596 236788 105602
rect 236736 105538 236788 105544
rect 236644 49020 236696 49026
rect 236644 48962 236696 48968
rect 235264 24132 235316 24138
rect 235264 24074 235316 24080
rect 236748 18630 236776 105538
rect 236840 104718 236868 146639
rect 236932 139534 236960 172518
rect 237392 168026 237420 235447
rect 238036 225622 238064 237458
rect 238312 237017 238340 240244
rect 238298 237008 238354 237017
rect 238298 236943 238354 236952
rect 238312 230353 238340 236943
rect 238298 230344 238354 230353
rect 238298 230279 238354 230288
rect 238864 229094 238892 240244
rect 239232 238202 239260 240244
rect 239220 238196 239272 238202
rect 239220 238138 239272 238144
rect 239404 237584 239456 237590
rect 239404 237526 239456 237532
rect 239416 236026 239444 237526
rect 239404 236020 239456 236026
rect 239404 235962 239456 235968
rect 238772 229066 238892 229094
rect 238024 225616 238076 225622
rect 238024 225558 238076 225564
rect 237562 210488 237618 210497
rect 237562 210423 237618 210432
rect 237472 209092 237524 209098
rect 237472 209034 237524 209040
rect 237380 168020 237432 168026
rect 237380 167962 237432 167968
rect 237012 165640 237064 165646
rect 237012 165582 237064 165588
rect 236920 139528 236972 139534
rect 236920 139470 236972 139476
rect 237024 135114 237052 165582
rect 237484 159633 237512 209034
rect 237576 162489 237604 210423
rect 238036 204241 238064 225558
rect 238772 220289 238800 229066
rect 239416 228585 239444 235962
rect 239402 228576 239458 228585
rect 239402 228511 239458 228520
rect 238758 220280 238814 220289
rect 238758 220215 238814 220224
rect 238772 220114 238800 220215
rect 238760 220108 238812 220114
rect 238760 220050 238812 220056
rect 239784 205601 239812 240244
rect 240336 238814 240364 240244
rect 240324 238808 240376 238814
rect 240324 238750 240376 238756
rect 240704 237289 240732 240244
rect 240876 238808 240928 238814
rect 240876 238750 240928 238756
rect 240690 237280 240746 237289
rect 240690 237215 240746 237224
rect 240046 233880 240102 233889
rect 240046 233815 240102 233824
rect 240060 231810 240088 233815
rect 240048 231804 240100 231810
rect 240048 231746 240100 231752
rect 240704 230489 240732 237215
rect 240784 234728 240836 234734
rect 240784 234670 240836 234676
rect 240690 230480 240746 230489
rect 240690 230415 240746 230424
rect 240796 212430 240824 234670
rect 240888 222154 240916 238750
rect 241256 233889 241284 240244
rect 241808 238678 241836 240244
rect 242176 240145 242204 240244
rect 242162 240136 242218 240145
rect 242162 240071 242218 240080
rect 242624 240100 242676 240106
rect 242624 240042 242676 240048
rect 241796 238672 241848 238678
rect 241796 238614 241848 238620
rect 241808 237425 241836 238614
rect 241794 237416 241850 237425
rect 241794 237351 241850 237360
rect 242636 236881 242664 240042
rect 242728 238754 242756 240244
rect 242728 238726 242848 238754
rect 242716 238196 242768 238202
rect 242716 238138 242768 238144
rect 242728 237153 242756 238138
rect 242820 237425 242848 238726
rect 242806 237416 242862 237425
rect 242806 237351 242862 237360
rect 242714 237144 242770 237153
rect 242714 237079 242770 237088
rect 242622 236872 242678 236881
rect 242622 236807 242678 236816
rect 241242 233880 241298 233889
rect 241242 233815 241298 233824
rect 242164 232620 242216 232626
rect 242164 232562 242216 232568
rect 240876 222148 240928 222154
rect 240876 222090 240928 222096
rect 240140 212424 240192 212430
rect 240140 212366 240192 212372
rect 240784 212424 240836 212430
rect 240784 212366 240836 212372
rect 239402 205592 239458 205601
rect 239402 205527 239458 205536
rect 239770 205592 239826 205601
rect 239770 205527 239826 205536
rect 238022 204232 238078 204241
rect 238022 204167 238078 204176
rect 239416 199442 239444 205527
rect 239404 199436 239456 199442
rect 239404 199378 239456 199384
rect 238760 193928 238812 193934
rect 238760 193870 238812 193876
rect 238208 173936 238260 173942
rect 238208 173878 238260 173884
rect 237562 162480 237618 162489
rect 237562 162415 237618 162424
rect 237470 159624 237526 159633
rect 237470 159559 237526 159568
rect 238116 151836 238168 151842
rect 238116 151778 238168 151784
rect 238024 138032 238076 138038
rect 238024 137974 238076 137980
rect 237012 135108 237064 135114
rect 237012 135050 237064 135056
rect 236920 117972 236972 117978
rect 236920 117914 236972 117920
rect 236828 104712 236880 104718
rect 236828 104654 236880 104660
rect 236932 91866 236960 117914
rect 236920 91860 236972 91866
rect 236920 91802 236972 91808
rect 238036 21486 238064 137974
rect 238128 110906 238156 151778
rect 238220 138854 238248 173878
rect 238300 157412 238352 157418
rect 238300 157354 238352 157360
rect 238208 138848 238260 138854
rect 238208 138790 238260 138796
rect 238206 129024 238262 129033
rect 238206 128959 238262 128968
rect 238116 110900 238168 110906
rect 238116 110842 238168 110848
rect 238116 103556 238168 103562
rect 238116 103498 238168 103504
rect 238024 21480 238076 21486
rect 238024 21422 238076 21428
rect 236736 18624 236788 18630
rect 236736 18566 236788 18572
rect 238128 10334 238156 103498
rect 238220 83502 238248 128959
rect 238312 119950 238340 157354
rect 238772 155922 238800 193870
rect 239404 192568 239456 192574
rect 239404 192510 239456 192516
rect 238850 180296 238906 180305
rect 238850 180231 238906 180240
rect 238760 155916 238812 155922
rect 238760 155858 238812 155864
rect 238864 152522 238892 180231
rect 239416 175982 239444 192510
rect 239404 175976 239456 175982
rect 239404 175918 239456 175924
rect 239496 175296 239548 175302
rect 239496 175238 239548 175244
rect 238852 152516 238904 152522
rect 238852 152458 238904 152464
rect 238392 151156 238444 151162
rect 238392 151098 238444 151104
rect 238404 129849 238432 151098
rect 239404 149728 239456 149734
rect 239404 149670 239456 149676
rect 238390 129840 238446 129849
rect 238390 129775 238446 129784
rect 239416 125361 239444 149670
rect 239402 125352 239458 125361
rect 239402 125287 239458 125296
rect 239402 123176 239458 123185
rect 239402 123111 239458 123120
rect 238300 119944 238352 119950
rect 238300 119886 238352 119892
rect 238298 110800 238354 110809
rect 238298 110735 238354 110744
rect 238208 83496 238260 83502
rect 238208 83438 238260 83444
rect 238312 77994 238340 110735
rect 238300 77988 238352 77994
rect 238300 77930 238352 77936
rect 239416 40798 239444 123111
rect 239508 99278 239536 175238
rect 239680 155236 239732 155242
rect 239680 155178 239732 155184
rect 239586 153232 239642 153241
rect 239586 153167 239642 153176
rect 239600 118017 239628 153167
rect 239692 131782 239720 155178
rect 240152 149161 240180 212366
rect 242176 209098 242204 232562
rect 242820 231849 242848 237351
rect 242806 231840 242862 231849
rect 242806 231775 242862 231784
rect 243280 209774 243308 240244
rect 243648 240009 243676 240244
rect 243634 240000 243690 240009
rect 243634 239935 243690 239944
rect 244016 238754 244044 244151
rect 243004 209746 243308 209774
rect 243924 238726 244044 238754
rect 243004 209681 243032 209746
rect 242990 209672 243046 209681
rect 242990 209607 243046 209616
rect 242164 209092 242216 209098
rect 242164 209034 242216 209040
rect 242900 206984 242952 206990
rect 242900 206926 242952 206932
rect 242912 206174 242940 206926
rect 242900 206168 242952 206174
rect 242900 206110 242952 206116
rect 240232 202156 240284 202162
rect 240232 202098 240284 202104
rect 240244 159458 240272 202098
rect 241612 195288 241664 195294
rect 241612 195230 241664 195236
rect 241520 182844 241572 182850
rect 241520 182786 241572 182792
rect 240324 178764 240376 178770
rect 240324 178706 240376 178712
rect 240336 170377 240364 178706
rect 240782 178120 240838 178129
rect 240782 178055 240838 178064
rect 240322 170368 240378 170377
rect 240322 170303 240378 170312
rect 240796 169833 240824 178055
rect 240782 169824 240838 169833
rect 240782 169759 240838 169768
rect 240876 169788 240928 169794
rect 240876 169730 240928 169736
rect 240782 168464 240838 168473
rect 240782 168399 240838 168408
rect 240232 159452 240284 159458
rect 240232 159394 240284 159400
rect 240138 149152 240194 149161
rect 240138 149087 240194 149096
rect 240796 144906 240824 168399
rect 240888 148374 240916 169730
rect 241060 158772 241112 158778
rect 241060 158714 241112 158720
rect 240876 148368 240928 148374
rect 240876 148310 240928 148316
rect 240968 147756 241020 147762
rect 240968 147698 241020 147704
rect 240876 146328 240928 146334
rect 240876 146270 240928 146276
rect 240784 144900 240836 144906
rect 240784 144842 240836 144848
rect 240782 143032 240838 143041
rect 240782 142967 240838 142976
rect 239680 131776 239732 131782
rect 239680 131718 239732 131724
rect 239678 124808 239734 124817
rect 239678 124743 239734 124752
rect 239586 118008 239642 118017
rect 239586 117943 239642 117952
rect 239586 102912 239642 102921
rect 239586 102847 239642 102856
rect 239496 99272 239548 99278
rect 239496 99214 239548 99220
rect 239600 82210 239628 102847
rect 239692 90438 239720 124743
rect 240796 121378 240824 142967
rect 240888 123457 240916 146270
rect 240874 123448 240930 123457
rect 240874 123383 240930 123392
rect 240784 121372 240836 121378
rect 240784 121314 240836 121320
rect 240876 119400 240928 119406
rect 240876 119342 240928 119348
rect 240784 118720 240836 118726
rect 240784 118662 240836 118668
rect 239680 90432 239732 90438
rect 239680 90374 239732 90380
rect 239588 82204 239640 82210
rect 239588 82146 239640 82152
rect 239404 40792 239456 40798
rect 239404 40734 239456 40740
rect 238116 10328 238168 10334
rect 238116 10270 238168 10276
rect 240796 7614 240824 118662
rect 240888 40730 240916 119342
rect 240980 106282 241008 147698
rect 241072 120086 241100 158714
rect 241532 150113 241560 182786
rect 241624 162790 241652 195230
rect 241702 174040 241758 174049
rect 241702 173975 241758 173984
rect 241612 162784 241664 162790
rect 241612 162726 241664 162732
rect 241716 158710 241744 173975
rect 242256 168496 242308 168502
rect 242256 168438 242308 168444
rect 241704 158704 241756 158710
rect 241704 158646 241756 158652
rect 242164 157480 242216 157486
rect 242164 157422 242216 157428
rect 241518 150104 241574 150113
rect 241518 150039 241574 150048
rect 241518 142896 241574 142905
rect 241518 142831 241520 142840
rect 241572 142831 241574 142840
rect 241520 142802 241572 142808
rect 241060 120080 241112 120086
rect 241060 120022 241112 120028
rect 242176 117298 242204 157422
rect 242268 129674 242296 168438
rect 242912 167113 242940 206110
rect 243004 172446 243032 209607
rect 243924 206174 243952 238726
rect 244280 229084 244332 229090
rect 244280 229026 244332 229032
rect 244292 228818 244320 229026
rect 244280 228812 244332 228818
rect 244280 228754 244332 228760
rect 243912 206168 243964 206174
rect 243912 206110 243964 206116
rect 243084 189100 243136 189106
rect 243084 189042 243136 189048
rect 242992 172440 243044 172446
rect 242992 172382 243044 172388
rect 242990 170504 243046 170513
rect 242990 170439 243046 170448
rect 242898 167104 242954 167113
rect 242898 167039 242954 167048
rect 242440 162852 242492 162858
rect 242440 162794 242492 162800
rect 242346 149696 242402 149705
rect 242346 149631 242402 149640
rect 242256 129668 242308 129674
rect 242256 129610 242308 129616
rect 242256 127016 242308 127022
rect 242256 126958 242308 126964
rect 242164 117292 242216 117298
rect 242164 117234 242216 117240
rect 242164 114572 242216 114578
rect 242164 114514 242216 114520
rect 241058 109440 241114 109449
rect 241058 109375 241114 109384
rect 240968 106276 241020 106282
rect 240968 106218 241020 106224
rect 241072 75313 241100 109375
rect 241058 75304 241114 75313
rect 241058 75239 241114 75248
rect 240876 40724 240928 40730
rect 240876 40666 240928 40672
rect 242176 17270 242204 114514
rect 242268 111081 242296 126958
rect 242254 111072 242310 111081
rect 242254 111007 242310 111016
rect 242360 109002 242388 149631
rect 242452 145897 242480 162794
rect 242438 145888 242494 145897
rect 242438 145823 242494 145832
rect 243004 136542 243032 170439
rect 243096 162858 243124 189042
rect 243176 177336 243228 177342
rect 243176 177278 243228 177284
rect 243084 162852 243136 162858
rect 243084 162794 243136 162800
rect 243188 155281 243216 177278
rect 243634 167104 243690 167113
rect 243634 167039 243690 167048
rect 243544 162852 243596 162858
rect 243544 162794 243596 162800
rect 243174 155272 243230 155281
rect 243174 155207 243230 155216
rect 243556 140729 243584 162794
rect 243542 140720 243598 140729
rect 243542 140655 243598 140664
rect 242992 136536 243044 136542
rect 242992 136478 243044 136484
rect 243544 135312 243596 135318
rect 243544 135254 243596 135260
rect 242438 113928 242494 113937
rect 242438 113863 242494 113872
rect 242348 108996 242400 109002
rect 242348 108938 242400 108944
rect 242254 107672 242310 107681
rect 242254 107607 242310 107616
rect 242268 60042 242296 107607
rect 242452 89078 242480 113863
rect 243452 93220 243504 93226
rect 243452 93162 243504 93168
rect 243464 90982 243492 93162
rect 243452 90976 243504 90982
rect 243452 90918 243504 90924
rect 242440 89072 242492 89078
rect 242440 89014 242492 89020
rect 242256 60036 242308 60042
rect 242256 59978 242308 59984
rect 243556 54534 243584 135254
rect 243648 126886 243676 167039
rect 244292 157350 244320 228754
rect 244384 210497 244412 261695
rect 244476 213858 244504 264415
rect 244464 213852 244516 213858
rect 244464 213794 244516 213800
rect 244370 210488 244426 210497
rect 244370 210423 244426 210432
rect 244372 196716 244424 196722
rect 244372 196658 244424 196664
rect 244384 171134 244412 196658
rect 244476 173194 244504 213794
rect 244936 175234 244964 273391
rect 245028 263022 245056 285738
rect 245672 273034 245700 294471
rect 245764 276729 245792 300154
rect 246316 290057 246344 322186
rect 246396 316056 246448 316062
rect 246396 315998 246448 316004
rect 246408 297430 246436 315998
rect 246396 297424 246448 297430
rect 246396 297366 246448 297372
rect 246302 290048 246358 290057
rect 246302 289983 246358 289992
rect 245844 287700 245896 287706
rect 245844 287642 245896 287648
rect 245856 287094 245884 287642
rect 245844 287088 245896 287094
rect 245844 287030 245896 287036
rect 245750 276720 245806 276729
rect 245750 276655 245752 276664
rect 245804 276655 245806 276664
rect 245752 276626 245804 276632
rect 245764 276595 245792 276626
rect 245856 274553 245884 287030
rect 247052 284594 247080 334591
rect 247132 296744 247184 296750
rect 247132 296686 247184 296692
rect 247144 291854 247172 296686
rect 248432 296041 248460 377590
rect 251376 374746 251404 377604
rect 252572 377590 253046 377618
rect 253952 377590 254702 377618
rect 255976 377590 256358 377618
rect 256712 377590 258014 377618
rect 259472 377590 259854 377618
rect 250444 374740 250496 374746
rect 250444 374682 250496 374688
rect 251364 374740 251416 374746
rect 251364 374682 251416 374688
rect 249064 345704 249116 345710
rect 249064 345646 249116 345652
rect 249076 345098 249104 345646
rect 249064 345092 249116 345098
rect 249064 345034 249116 345040
rect 248512 335368 248564 335374
rect 248512 335310 248564 335316
rect 248418 296032 248474 296041
rect 248418 295967 248474 295976
rect 247132 291848 247184 291854
rect 247132 291790 247184 291796
rect 247316 291304 247368 291310
rect 247316 291246 247368 291252
rect 247132 291236 247184 291242
rect 247132 291178 247184 291184
rect 246868 284566 247080 284594
rect 246868 283626 246896 284566
rect 247040 284436 247092 284442
rect 247040 284378 247092 284384
rect 247052 284322 247080 284378
rect 246960 284294 247080 284322
rect 246960 283801 246988 284294
rect 246946 283792 247002 283801
rect 246946 283727 247002 283736
rect 246304 283620 246356 283626
rect 246304 283562 246356 283568
rect 246856 283620 246908 283626
rect 246856 283562 246908 283568
rect 246316 283257 246344 283562
rect 246302 283248 246358 283257
rect 246302 283183 246358 283192
rect 245936 281716 245988 281722
rect 245936 281658 245988 281664
rect 245948 281625 245976 281658
rect 245934 281616 245990 281625
rect 245934 281551 245990 281560
rect 246118 281072 246174 281081
rect 246118 281007 246174 281016
rect 246132 280226 246160 281007
rect 246120 280220 246172 280226
rect 246120 280162 246172 280168
rect 245936 279540 245988 279546
rect 245936 279482 245988 279488
rect 245948 279449 245976 279482
rect 245934 279440 245990 279449
rect 245934 279375 245990 279384
rect 245936 278996 245988 279002
rect 245936 278938 245988 278944
rect 245948 278905 245976 278938
rect 245934 278896 245990 278905
rect 245934 278831 245990 278840
rect 245936 278044 245988 278050
rect 245936 277986 245988 277992
rect 245948 277545 245976 277986
rect 245934 277536 245990 277545
rect 245934 277471 245990 277480
rect 245936 276004 245988 276010
rect 245936 275946 245988 275952
rect 245948 275913 245976 275946
rect 245934 275904 245990 275913
rect 245934 275839 245990 275848
rect 245934 275360 245990 275369
rect 245934 275295 245936 275304
rect 245988 275295 245990 275304
rect 245936 275266 245988 275272
rect 245842 274544 245898 274553
rect 245842 274479 245898 274488
rect 245844 273216 245896 273222
rect 245842 273184 245844 273193
rect 245896 273184 245898 273193
rect 245842 273119 245898 273128
rect 245672 273006 245884 273034
rect 245856 271182 245884 273006
rect 245936 272536 245988 272542
rect 245936 272478 245988 272484
rect 245948 272377 245976 272478
rect 245934 272368 245990 272377
rect 245934 272303 245990 272312
rect 245934 271552 245990 271561
rect 245934 271487 245990 271496
rect 245948 271250 245976 271487
rect 245936 271244 245988 271250
rect 245936 271186 245988 271192
rect 245844 271176 245896 271182
rect 245844 271118 245896 271124
rect 245856 271017 245884 271118
rect 245842 271008 245898 271017
rect 245842 270943 245898 270952
rect 245948 270230 245976 270261
rect 245936 270224 245988 270230
rect 245934 270192 245936 270201
rect 245988 270192 245990 270201
rect 245934 270127 245990 270136
rect 245752 267708 245804 267714
rect 245752 267650 245804 267656
rect 245764 266665 245792 267650
rect 245750 266656 245806 266665
rect 245750 266591 245806 266600
rect 245842 265840 245898 265849
rect 245842 265775 245898 265784
rect 245856 265674 245884 265775
rect 245844 265668 245896 265674
rect 245844 265610 245896 265616
rect 245016 263016 245068 263022
rect 245016 262958 245068 262964
rect 245842 262304 245898 262313
rect 245842 262239 245844 262248
rect 245896 262239 245898 262248
rect 245844 262210 245896 262216
rect 245658 259584 245714 259593
rect 245658 259519 245714 259528
rect 245672 259486 245700 259519
rect 245660 259480 245712 259486
rect 245660 259422 245712 259428
rect 245844 259412 245896 259418
rect 245844 259354 245896 259360
rect 245658 258768 245714 258777
rect 245658 258703 245714 258712
rect 245672 258126 245700 258703
rect 245856 258233 245884 259354
rect 245842 258224 245898 258233
rect 245842 258159 245898 258168
rect 245660 258120 245712 258126
rect 245660 258062 245712 258068
rect 245844 258052 245896 258058
rect 245844 257994 245896 258000
rect 245856 257417 245884 257994
rect 245842 257408 245898 257417
rect 245842 257343 245898 257352
rect 245844 256692 245896 256698
rect 245844 256634 245896 256640
rect 245856 256601 245884 256634
rect 245842 256592 245898 256601
rect 245842 256527 245898 256536
rect 245844 256080 245896 256086
rect 245842 256048 245844 256057
rect 245896 256048 245898 256057
rect 245842 255983 245898 255992
rect 245842 255232 245898 255241
rect 245842 255167 245844 255176
rect 245896 255167 245898 255176
rect 245844 255138 245896 255144
rect 245658 253872 245714 253881
rect 245658 253807 245714 253816
rect 245672 252618 245700 253807
rect 245660 252612 245712 252618
rect 245660 252554 245712 252560
rect 245844 252272 245896 252278
rect 245842 252240 245844 252249
rect 245896 252240 245898 252249
rect 245842 252175 245898 252184
rect 245658 250880 245714 250889
rect 245658 250815 245714 250824
rect 245672 247110 245700 250815
rect 245842 247344 245898 247353
rect 245842 247279 245898 247288
rect 245856 247110 245884 247279
rect 245016 247104 245068 247110
rect 245016 247046 245068 247052
rect 245660 247104 245712 247110
rect 245660 247046 245712 247052
rect 245844 247104 245896 247110
rect 245844 247046 245896 247052
rect 245028 228818 245056 247046
rect 245660 246424 245712 246430
rect 245660 246366 245712 246372
rect 245672 245993 245700 246366
rect 245658 245984 245714 245993
rect 245658 245919 245714 245928
rect 245750 243808 245806 243817
rect 245750 243743 245806 243752
rect 245764 243030 245792 243743
rect 245752 243024 245804 243030
rect 245752 242966 245804 242972
rect 245658 241632 245714 241641
rect 245658 241567 245714 241576
rect 245672 240786 245700 241567
rect 245842 240816 245898 240825
rect 245660 240780 245712 240786
rect 245842 240751 245898 240760
rect 245660 240722 245712 240728
rect 245672 240242 245700 240722
rect 245660 240236 245712 240242
rect 245660 240178 245712 240184
rect 245016 228812 245068 228818
rect 245016 228754 245068 228760
rect 245750 214840 245806 214849
rect 245750 214775 245806 214784
rect 245658 178664 245714 178673
rect 245658 178599 245714 178608
rect 244924 175228 244976 175234
rect 244924 175170 244976 175176
rect 245016 174004 245068 174010
rect 245016 173946 245068 173952
rect 244464 173188 244516 173194
rect 244464 173130 244516 173136
rect 244384 171106 244504 171134
rect 244370 169824 244426 169833
rect 244370 169759 244426 169768
rect 244384 162858 244412 169759
rect 244476 165073 244504 171106
rect 244462 165064 244518 165073
rect 244462 164999 244518 165008
rect 244372 162852 244424 162858
rect 244372 162794 244424 162800
rect 244280 157344 244332 157350
rect 244280 157286 244332 157292
rect 243818 154864 243874 154873
rect 243818 154799 243874 154808
rect 243636 126880 243688 126886
rect 243636 126822 243688 126828
rect 243728 126268 243780 126274
rect 243728 126210 243780 126216
rect 243634 117600 243690 117609
rect 243634 117535 243690 117544
rect 243544 54528 243596 54534
rect 243544 54470 243596 54476
rect 243648 50289 243676 117535
rect 243740 84862 243768 126210
rect 243832 114442 243860 154799
rect 244922 150920 244978 150929
rect 244922 150855 244978 150864
rect 244280 142860 244332 142866
rect 244280 142802 244332 142808
rect 244292 142497 244320 142802
rect 244278 142488 244334 142497
rect 244278 142423 244334 142432
rect 243820 114436 243872 114442
rect 243820 114378 243872 114384
rect 244936 110362 244964 150855
rect 245028 136610 245056 173946
rect 245108 163532 245160 163538
rect 245108 163474 245160 163480
rect 245016 136604 245068 136610
rect 245016 136546 245068 136552
rect 245120 128314 245148 163474
rect 245200 160132 245252 160138
rect 245200 160074 245252 160080
rect 245108 128308 245160 128314
rect 245108 128250 245160 128256
rect 245212 124914 245240 160074
rect 245672 138825 245700 178599
rect 245764 148209 245792 214775
rect 245856 207670 245884 240751
rect 245844 207664 245896 207670
rect 245844 207606 245896 207612
rect 245844 205692 245896 205698
rect 245844 205634 245896 205640
rect 245856 153882 245884 205634
rect 245948 172825 245976 270127
rect 246302 269648 246358 269657
rect 246302 269583 246358 269592
rect 246028 266348 246080 266354
rect 246028 266290 246080 266296
rect 246040 265305 246068 266290
rect 246026 265296 246082 265305
rect 246026 265231 246082 265240
rect 246028 260840 246080 260846
rect 246028 260782 246080 260788
rect 246040 260137 246068 260782
rect 246026 260128 246082 260137
rect 246026 260063 246082 260072
rect 246028 255264 246080 255270
rect 246028 255206 246080 255212
rect 246040 254425 246068 255206
rect 246026 254416 246082 254425
rect 246026 254351 246082 254360
rect 246028 253904 246080 253910
rect 246028 253846 246080 253852
rect 246040 253065 246068 253846
rect 246026 253056 246082 253065
rect 246026 252991 246082 253000
rect 246028 252544 246080 252550
rect 246028 252486 246080 252492
rect 246040 251705 246068 252486
rect 246026 251696 246082 251705
rect 246026 251631 246082 251640
rect 246028 249756 246080 249762
rect 246028 249698 246080 249704
rect 246040 249529 246068 249698
rect 246026 249520 246082 249529
rect 246026 249455 246082 249464
rect 246316 246362 246344 269583
rect 246396 263016 246448 263022
rect 246396 262958 246448 262964
rect 246304 246356 246356 246362
rect 246304 246298 246356 246304
rect 246026 245168 246082 245177
rect 246026 245103 246082 245112
rect 246040 234734 246068 245103
rect 246408 244254 246436 262958
rect 247144 260953 247172 291178
rect 247222 282432 247278 282441
rect 247222 282367 247278 282376
rect 247130 260944 247186 260953
rect 247130 260879 247186 260888
rect 247040 253972 247092 253978
rect 247040 253914 247092 253920
rect 246396 244248 246448 244254
rect 246396 244190 246448 244196
rect 246118 242448 246174 242457
rect 246118 242383 246174 242392
rect 246132 241534 246160 242383
rect 246120 241528 246172 241534
rect 246120 241470 246172 241476
rect 246028 234728 246080 234734
rect 246028 234670 246080 234676
rect 246132 224262 246160 241470
rect 246120 224256 246172 224262
rect 246120 224198 246172 224204
rect 245934 172816 245990 172825
rect 245934 172751 245990 172760
rect 246302 171728 246358 171737
rect 246302 171663 246358 171672
rect 246316 158001 246344 171663
rect 247052 170406 247080 253914
rect 247130 248704 247186 248713
rect 247130 248639 247186 248648
rect 247144 226302 247172 248639
rect 247132 226296 247184 226302
rect 247132 226238 247184 226244
rect 247040 170400 247092 170406
rect 247040 170342 247092 170348
rect 246302 157992 246358 158001
rect 246302 157927 246358 157936
rect 246304 155984 246356 155990
rect 246304 155926 246356 155932
rect 245844 153876 245896 153882
rect 245844 153818 245896 153824
rect 245750 148200 245806 148209
rect 245750 148135 245806 148144
rect 245658 138816 245714 138825
rect 245658 138751 245714 138760
rect 245200 124908 245252 124914
rect 245200 124850 245252 124856
rect 245292 124908 245344 124914
rect 245292 124850 245344 124856
rect 245108 113212 245160 113218
rect 245108 113154 245160 113160
rect 244924 110356 244976 110362
rect 244924 110298 244976 110304
rect 245014 99512 245070 99521
rect 245014 99447 245070 99456
rect 243728 84856 243780 84862
rect 243728 84798 243780 84804
rect 244924 75880 244976 75886
rect 244924 75822 244976 75828
rect 243634 50280 243690 50289
rect 243634 50215 243690 50224
rect 242164 17264 242216 17270
rect 242164 17206 242216 17212
rect 243544 17264 243596 17270
rect 243544 17206 243596 17212
rect 242164 11756 242216 11762
rect 242164 11698 242216 11704
rect 240784 7608 240836 7614
rect 240784 7550 240836 7556
rect 233884 6180 233936 6186
rect 233884 6122 233936 6128
rect 232596 4208 232648 4214
rect 232596 4150 232648 4156
rect 235816 4208 235868 4214
rect 235816 4150 235868 4156
rect 220084 3460 220136 3466
rect 220084 3402 220136 3408
rect 213184 2168 213236 2174
rect 213184 2110 213236 2116
rect 177394 2000 177450 2009
rect 177394 1935 177450 1944
rect 235828 480 235856 4150
rect 240508 3392 240560 3398
rect 240508 3334 240560 3340
rect 239312 2168 239364 2174
rect 239312 2110 239364 2116
rect 239324 480 239352 2110
rect 240520 480 240548 3334
rect 241704 3324 241756 3330
rect 241704 3266 241756 3272
rect 241716 480 241744 3266
rect 242176 2106 242204 11698
rect 243556 9654 243584 17206
rect 242900 9648 242952 9654
rect 242900 9590 242952 9596
rect 243544 9648 243596 9654
rect 243544 9590 243596 9596
rect 242164 2100 242216 2106
rect 242164 2042 242216 2048
rect 242912 480 242940 9590
rect 244094 4992 244150 5001
rect 244094 4927 244150 4936
rect 244108 480 244136 4927
rect 244936 3330 244964 75822
rect 245028 43450 245056 99447
rect 245120 64161 245148 113154
rect 245200 104916 245252 104922
rect 245200 104858 245252 104864
rect 245212 68377 245240 104858
rect 245304 100638 245332 124850
rect 246316 115569 246344 155926
rect 246486 153776 246542 153785
rect 246486 153711 246542 153720
rect 246394 132832 246450 132841
rect 246394 132767 246450 132776
rect 246302 115560 246358 115569
rect 246302 115495 246358 115504
rect 245292 100632 245344 100638
rect 245292 100574 245344 100580
rect 246304 98660 246356 98666
rect 246304 98602 246356 98608
rect 245198 68368 245254 68377
rect 245198 68303 245254 68312
rect 245106 64152 245162 64161
rect 245106 64087 245162 64096
rect 245016 43444 245068 43450
rect 245016 43386 245068 43392
rect 246316 31074 246344 98602
rect 246408 71097 246436 132767
rect 246500 115938 246528 153711
rect 247144 151065 247172 226238
rect 247236 223553 247264 282367
rect 247328 255202 247356 291246
rect 248420 289944 248472 289950
rect 248420 289886 248472 289892
rect 247500 288448 247552 288454
rect 247500 288390 247552 288396
rect 247512 282198 247540 288390
rect 247682 285152 247738 285161
rect 247682 285087 247738 285096
rect 247696 284442 247724 285087
rect 247684 284436 247736 284442
rect 247684 284378 247736 284384
rect 247500 282192 247552 282198
rect 247500 282134 247552 282140
rect 247316 255196 247368 255202
rect 247316 255138 247368 255144
rect 247328 253978 247356 255138
rect 247316 253972 247368 253978
rect 247316 253914 247368 253920
rect 247314 250336 247370 250345
rect 247314 250271 247370 250280
rect 247328 249830 247356 250271
rect 247316 249824 247368 249830
rect 247316 249766 247368 249772
rect 247328 239873 247356 249766
rect 247314 239864 247370 239873
rect 247314 239799 247370 239808
rect 247222 223544 247278 223553
rect 247222 223479 247278 223488
rect 247236 159089 247264 223479
rect 247684 169856 247736 169862
rect 247684 169798 247736 169804
rect 247222 159080 247278 159089
rect 247222 159015 247278 159024
rect 247130 151056 247186 151065
rect 247130 150991 247186 151000
rect 246578 137184 246634 137193
rect 246578 137119 246634 137128
rect 246488 115932 246540 115938
rect 246488 115874 246540 115880
rect 246592 105602 246620 137119
rect 247696 131034 247724 169798
rect 247776 164280 247828 164286
rect 247776 164222 247828 164228
rect 247788 143177 247816 164222
rect 248432 164218 248460 289886
rect 248524 270230 248552 335310
rect 248604 273216 248656 273222
rect 248602 273184 248604 273193
rect 248656 273184 248658 273193
rect 248602 273119 248658 273128
rect 248604 271244 248656 271250
rect 248604 271186 248656 271192
rect 248512 270224 248564 270230
rect 248512 270166 248564 270172
rect 248512 262268 248564 262274
rect 248512 262210 248564 262216
rect 248524 202774 248552 262210
rect 248616 236706 248644 271186
rect 248604 236700 248656 236706
rect 248604 236642 248656 236648
rect 249076 219434 249104 345034
rect 249800 331900 249852 331906
rect 249800 331842 249852 331848
rect 249154 310040 249210 310049
rect 249154 309975 249210 309984
rect 249168 299538 249196 309975
rect 249156 299532 249208 299538
rect 249156 299474 249208 299480
rect 249168 279002 249196 299474
rect 249156 278996 249208 279002
rect 249156 278938 249208 278944
rect 249812 252278 249840 331842
rect 249892 278044 249944 278050
rect 249892 277986 249944 277992
rect 249800 252272 249852 252278
rect 249800 252214 249852 252220
rect 249904 232665 249932 277986
rect 249984 244248 250036 244254
rect 249984 244190 250036 244196
rect 249890 232656 249946 232665
rect 249890 232591 249946 232600
rect 249800 229832 249852 229838
rect 249800 229774 249852 229780
rect 249812 225690 249840 229774
rect 249800 225684 249852 225690
rect 249800 225626 249852 225632
rect 248984 219406 249104 219434
rect 248984 216578 249012 219406
rect 248972 216572 249024 216578
rect 248972 216514 249024 216520
rect 249708 216572 249760 216578
rect 249708 216514 249760 216520
rect 249720 215966 249748 216514
rect 249708 215960 249760 215966
rect 249708 215902 249760 215908
rect 248512 202768 248564 202774
rect 248512 202710 248564 202716
rect 248524 200114 248552 202710
rect 248524 200086 248644 200114
rect 248510 187776 248566 187785
rect 248510 187711 248566 187720
rect 248420 164212 248472 164218
rect 248420 164154 248472 164160
rect 248524 146946 248552 187711
rect 248616 172514 248644 200086
rect 249996 190454 250024 244190
rect 250456 196654 250484 374682
rect 252572 369918 252600 377590
rect 253952 370530 253980 377590
rect 253940 370524 253992 370530
rect 253940 370466 253992 370472
rect 252560 369912 252612 369918
rect 252560 369854 252612 369860
rect 253296 369912 253348 369918
rect 253296 369854 253348 369860
rect 253204 369164 253256 369170
rect 253204 369106 253256 369112
rect 251914 353424 251970 353433
rect 251914 353359 251970 353368
rect 251824 348492 251876 348498
rect 251824 348434 251876 348440
rect 251272 318096 251324 318102
rect 251272 318038 251324 318044
rect 250626 302424 250682 302433
rect 250626 302359 250682 302368
rect 250534 285832 250590 285841
rect 250534 285767 250590 285776
rect 250548 257378 250576 285767
rect 250640 281518 250668 302359
rect 251180 283620 251232 283626
rect 251180 283562 251232 283568
rect 251086 282840 251142 282849
rect 251086 282775 251142 282784
rect 251100 281722 251128 282775
rect 251088 281716 251140 281722
rect 251088 281658 251140 281664
rect 250628 281512 250680 281518
rect 250628 281454 250680 281460
rect 250536 257372 250588 257378
rect 250536 257314 250588 257320
rect 251088 252272 251140 252278
rect 251088 252214 251140 252220
rect 251100 251841 251128 252214
rect 251086 251832 251142 251841
rect 251086 251767 251142 251776
rect 250534 213208 250590 213217
rect 250534 213143 250590 213152
rect 250548 207670 250576 213143
rect 250536 207664 250588 207670
rect 250536 207606 250588 207612
rect 250444 196648 250496 196654
rect 250444 196590 250496 196596
rect 249904 190426 250024 190454
rect 249800 188352 249852 188358
rect 249800 188294 249852 188300
rect 248604 172508 248656 172514
rect 248604 172450 248656 172456
rect 249340 171148 249392 171154
rect 249340 171090 249392 171096
rect 249064 165708 249116 165714
rect 249064 165650 249116 165656
rect 248512 146940 248564 146946
rect 248512 146882 248564 146888
rect 247868 144220 247920 144226
rect 247868 144162 247920 144168
rect 247774 143168 247830 143177
rect 247774 143103 247830 143112
rect 247684 131028 247736 131034
rect 247684 130970 247736 130976
rect 247774 124672 247830 124681
rect 247774 124607 247830 124616
rect 247684 110492 247736 110498
rect 247684 110434 247736 110440
rect 246580 105596 246632 105602
rect 246580 105538 246632 105544
rect 246488 96688 246540 96694
rect 246488 96630 246540 96636
rect 246500 86970 246528 96630
rect 246488 86964 246540 86970
rect 246488 86906 246540 86912
rect 247038 86320 247094 86329
rect 247038 86255 247094 86264
rect 247052 75886 247080 86255
rect 247040 75880 247092 75886
rect 247040 75822 247092 75828
rect 246394 71088 246450 71097
rect 246394 71023 246450 71032
rect 247696 58682 247724 110434
rect 247788 80782 247816 124607
rect 247880 104854 247908 144162
rect 247960 141500 248012 141506
rect 247960 141442 248012 141448
rect 247972 110401 248000 141442
rect 248052 139460 248104 139466
rect 248052 139402 248104 139408
rect 248064 123486 248092 139402
rect 249076 126954 249104 165650
rect 249248 151904 249300 151910
rect 249248 151846 249300 151852
rect 249156 143608 249208 143614
rect 249156 143550 249208 143556
rect 249064 126948 249116 126954
rect 249064 126890 249116 126896
rect 248052 123480 248104 123486
rect 248052 123422 248104 123428
rect 248418 123448 248474 123457
rect 248418 123383 248474 123392
rect 248432 117978 248460 123383
rect 249064 121508 249116 121514
rect 249064 121450 249116 121456
rect 248420 117972 248472 117978
rect 248420 117914 248472 117920
rect 247958 110392 248014 110401
rect 247958 110327 248014 110336
rect 247958 108080 248014 108089
rect 247958 108015 248014 108024
rect 247868 104848 247920 104854
rect 247868 104790 247920 104796
rect 247972 94518 248000 108015
rect 247960 94512 248012 94518
rect 247960 94454 248012 94460
rect 247776 80776 247828 80782
rect 247776 80718 247828 80724
rect 247684 58676 247736 58682
rect 247684 58618 247736 58624
rect 248328 58676 248380 58682
rect 248328 58618 248380 58624
rect 246396 43444 246448 43450
rect 246396 43386 246448 43392
rect 246304 31068 246356 31074
rect 246304 31010 246356 31016
rect 245660 18692 245712 18698
rect 245660 18634 245712 18640
rect 245672 16574 245700 18634
rect 245672 16546 245976 16574
rect 245658 3904 245714 3913
rect 245658 3839 245714 3848
rect 245672 3466 245700 3839
rect 245660 3460 245712 3466
rect 245660 3402 245712 3408
rect 244924 3324 244976 3330
rect 244924 3266 244976 3272
rect 245200 2984 245252 2990
rect 245200 2926 245252 2932
rect 245212 480 245240 2926
rect 245948 490 245976 16546
rect 246408 3398 246436 43386
rect 248340 36718 248368 58618
rect 247040 36712 247092 36718
rect 247040 36654 247092 36660
rect 248328 36712 248380 36718
rect 248328 36654 248380 36660
rect 246396 3392 246448 3398
rect 246396 3334 246448 3340
rect 247052 2990 247080 36654
rect 249076 19990 249104 121450
rect 249168 103494 249196 143550
rect 249260 111790 249288 151846
rect 249352 132462 249380 171090
rect 249708 160744 249760 160750
rect 249708 160686 249760 160692
rect 249720 155242 249748 160686
rect 249708 155236 249760 155242
rect 249708 155178 249760 155184
rect 249812 137970 249840 188294
rect 249904 185638 249932 190426
rect 249892 185632 249944 185638
rect 249892 185574 249944 185580
rect 249904 185473 249932 185574
rect 249890 185464 249946 185473
rect 249890 185399 249946 185408
rect 250536 172644 250588 172650
rect 250536 172586 250588 172592
rect 250444 154692 250496 154698
rect 250444 154634 250496 154640
rect 249800 137964 249852 137970
rect 249800 137906 249852 137912
rect 249340 132456 249392 132462
rect 249340 132398 249392 132404
rect 250456 114510 250484 154634
rect 250548 135250 250576 172586
rect 250628 156052 250680 156058
rect 250628 155994 250680 156000
rect 250536 135244 250588 135250
rect 250536 135186 250588 135192
rect 250640 124982 250668 155994
rect 251192 144129 251220 283562
rect 251284 273222 251312 318038
rect 251364 301572 251416 301578
rect 251364 301514 251416 301520
rect 251272 273216 251324 273222
rect 251272 273158 251324 273164
rect 251270 273048 251326 273057
rect 251270 272983 251326 272992
rect 251284 272542 251312 272983
rect 251272 272536 251324 272542
rect 251272 272478 251324 272484
rect 251270 270464 251326 270473
rect 251270 270399 251326 270408
rect 251284 205057 251312 270399
rect 251376 255270 251404 301514
rect 251364 255264 251416 255270
rect 251364 255206 251416 255212
rect 251836 249762 251864 348434
rect 251928 340882 251956 353359
rect 253216 349897 253244 369106
rect 253308 355337 253336 369854
rect 255976 369170 256004 377590
rect 256056 369232 256108 369238
rect 256056 369174 256108 369180
rect 255964 369164 256016 369170
rect 255964 369106 256016 369112
rect 254582 356688 254638 356697
rect 254582 356623 254638 356632
rect 253294 355328 253350 355337
rect 253294 355263 253350 355272
rect 253202 349888 253258 349897
rect 253202 349823 253258 349832
rect 252560 340944 252612 340950
rect 252560 340886 252612 340892
rect 251916 340876 251968 340882
rect 251916 340818 251968 340824
rect 251916 334688 251968 334694
rect 251916 334630 251968 334636
rect 251928 324970 251956 334630
rect 251916 324964 251968 324970
rect 251916 324906 251968 324912
rect 252468 272536 252520 272542
rect 252468 272478 252520 272484
rect 252480 271930 252508 272478
rect 252468 271924 252520 271930
rect 252468 271866 252520 271872
rect 252572 265674 252600 340886
rect 252652 338156 252704 338162
rect 252652 338098 252704 338104
rect 252560 265668 252612 265674
rect 252560 265610 252612 265616
rect 252468 255264 252520 255270
rect 252468 255206 252520 255212
rect 252480 254658 252508 255206
rect 252468 254652 252520 254658
rect 252468 254594 252520 254600
rect 252468 249892 252520 249898
rect 252468 249834 252520 249840
rect 252480 249762 252508 249834
rect 251824 249756 251876 249762
rect 251824 249698 251876 249704
rect 252468 249756 252520 249762
rect 252468 249698 252520 249704
rect 251822 247072 251878 247081
rect 251822 247007 251878 247016
rect 251836 225729 251864 247007
rect 251822 225720 251878 225729
rect 251822 225655 251878 225664
rect 251916 209092 251968 209098
rect 251916 209034 251968 209040
rect 251822 207632 251878 207641
rect 251822 207567 251878 207576
rect 251270 205048 251326 205057
rect 251270 204983 251326 204992
rect 251178 144120 251234 144129
rect 251178 144055 251234 144064
rect 250812 135380 250864 135386
rect 250812 135322 250864 135328
rect 250720 134564 250772 134570
rect 250720 134506 250772 134512
rect 250628 124976 250680 124982
rect 250628 124918 250680 124924
rect 250536 114640 250588 114646
rect 250536 114582 250588 114588
rect 250444 114504 250496 114510
rect 250444 114446 250496 114452
rect 249248 111784 249300 111790
rect 249248 111726 249300 111732
rect 249156 103488 249208 103494
rect 249156 103430 249208 103436
rect 249248 102196 249300 102202
rect 249248 102138 249300 102144
rect 249154 75168 249210 75177
rect 249154 75103 249210 75112
rect 249064 19984 249116 19990
rect 249064 19926 249116 19932
rect 249168 16590 249196 75103
rect 249260 69698 249288 102138
rect 250442 98424 250498 98433
rect 250442 98359 250498 98368
rect 249248 69692 249300 69698
rect 249248 69634 249300 69640
rect 250456 42090 250484 98359
rect 250548 58585 250576 114582
rect 250626 109304 250682 109313
rect 250626 109239 250682 109248
rect 250640 62937 250668 109239
rect 250732 99346 250760 134506
rect 250824 124817 250852 135322
rect 250810 124808 250866 124817
rect 250810 124743 250866 124752
rect 250812 122868 250864 122874
rect 250812 122810 250864 122816
rect 250720 99340 250772 99346
rect 250720 99282 250772 99288
rect 250824 89010 250852 122810
rect 250812 89004 250864 89010
rect 250812 88946 250864 88952
rect 250626 62928 250682 62937
rect 250626 62863 250682 62872
rect 250534 58576 250590 58585
rect 250534 58511 250590 58520
rect 250536 51808 250588 51814
rect 250536 51750 250588 51756
rect 250444 42084 250496 42090
rect 250444 42026 250496 42032
rect 250444 19984 250496 19990
rect 250444 19926 250496 19932
rect 249156 16584 249208 16590
rect 250456 16574 250484 19926
rect 249156 16526 249208 16532
rect 249996 16546 250484 16574
rect 249168 15230 249196 16526
rect 248420 15224 248472 15230
rect 248420 15166 248472 15172
rect 249156 15224 249208 15230
rect 249996 15201 250024 16546
rect 249156 15166 249208 15172
rect 249982 15192 250038 15201
rect 247776 4140 247828 4146
rect 247776 4082 247828 4088
rect 247788 3369 247816 4082
rect 247590 3360 247646 3369
rect 247590 3295 247646 3304
rect 247774 3360 247830 3369
rect 247774 3295 247830 3304
rect 247040 2984 247092 2990
rect 247040 2926 247092 2932
rect 246224 598 246436 626
rect 246224 490 246252 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 462 246252 490
rect 246408 480 246436 598
rect 247604 480 247632 3295
rect 248432 490 248460 15166
rect 249982 15127 250038 15136
rect 248616 598 248828 626
rect 248616 490 248644 598
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 462 248644 490
rect 248800 480 248828 598
rect 249996 480 250024 15127
rect 250548 4146 250576 51750
rect 250536 4140 250588 4146
rect 250536 4082 250588 4088
rect 251836 3641 251864 207567
rect 251928 196654 251956 209034
rect 251916 196648 251968 196654
rect 251916 196590 251968 196596
rect 252098 169008 252154 169017
rect 252098 168943 252154 168952
rect 252008 131164 252060 131170
rect 252008 131106 252060 131112
rect 251916 128376 251968 128382
rect 251916 128318 251968 128324
rect 251928 47569 251956 128318
rect 252020 59945 252048 131106
rect 252112 129742 252140 168943
rect 252192 162920 252244 162926
rect 252192 162862 252244 162868
rect 252100 129736 252152 129742
rect 252100 129678 252152 129684
rect 252204 124166 252232 162862
rect 252572 153105 252600 265610
rect 252664 238678 252692 338098
rect 254596 298081 254624 356623
rect 255962 349888 256018 349897
rect 255962 349823 256018 349832
rect 254676 321632 254728 321638
rect 254676 321574 254728 321580
rect 254688 311234 254716 321574
rect 255504 314696 255556 314702
rect 255504 314638 255556 314644
rect 254676 311228 254728 311234
rect 254676 311170 254728 311176
rect 255410 311128 255466 311137
rect 255410 311063 255466 311072
rect 254676 298784 254728 298790
rect 254676 298726 254728 298732
rect 254030 298072 254086 298081
rect 254030 298007 254086 298016
rect 254582 298072 254638 298081
rect 254582 298007 254638 298016
rect 254044 297401 254072 298007
rect 254030 297392 254086 297401
rect 254030 297327 254086 297336
rect 253204 292664 253256 292670
rect 253204 292606 253256 292612
rect 253216 286385 253244 292606
rect 253940 291848 253992 291854
rect 253940 291790 253992 291796
rect 253846 288552 253902 288561
rect 253846 288487 253902 288496
rect 253202 286376 253258 286385
rect 253202 286311 253258 286320
rect 253294 285016 253350 285025
rect 253294 284951 253350 284960
rect 253204 281716 253256 281722
rect 253204 281658 253256 281664
rect 252834 275768 252890 275777
rect 252834 275703 252890 275712
rect 252848 275330 252876 275703
rect 252836 275324 252888 275330
rect 252836 275266 252888 275272
rect 252848 274718 252876 275266
rect 252836 274712 252888 274718
rect 252836 274654 252888 274660
rect 253112 246424 253164 246430
rect 253112 246366 253164 246372
rect 253124 245857 253152 246366
rect 253110 245848 253166 245857
rect 253110 245783 253166 245792
rect 252652 238672 252704 238678
rect 252652 238614 252704 238620
rect 253216 156777 253244 281658
rect 253308 269249 253336 284951
rect 253860 282169 253888 288487
rect 253846 282160 253902 282169
rect 253846 282095 253902 282104
rect 253294 269240 253350 269249
rect 253294 269175 253350 269184
rect 253294 172816 253350 172825
rect 253294 172751 253350 172760
rect 253202 156768 253258 156777
rect 253202 156703 253258 156712
rect 253204 153264 253256 153270
rect 253204 153206 253256 153212
rect 252558 153096 252614 153105
rect 252558 153031 252614 153040
rect 252192 124160 252244 124166
rect 252192 124102 252244 124108
rect 252100 122936 252152 122942
rect 252100 122878 252152 122884
rect 252112 78033 252140 122878
rect 253216 113082 253244 153206
rect 253308 133822 253336 172751
rect 253386 148336 253442 148345
rect 253386 148271 253442 148280
rect 253296 133816 253348 133822
rect 253296 133758 253348 133764
rect 253296 116000 253348 116006
rect 253296 115942 253348 115948
rect 253204 113076 253256 113082
rect 253204 113018 253256 113024
rect 253204 107704 253256 107710
rect 253204 107646 253256 107652
rect 252098 78024 252154 78033
rect 252098 77959 252154 77968
rect 252006 59936 252062 59945
rect 252006 59871 252062 59880
rect 251914 47560 251970 47569
rect 251914 47495 251970 47504
rect 253216 44878 253244 107646
rect 253308 65521 253336 115942
rect 253400 109041 253428 148271
rect 253952 139777 253980 291790
rect 254044 213897 254072 297327
rect 254122 287736 254178 287745
rect 254122 287671 254178 287680
rect 254136 256698 254164 287671
rect 254688 284986 254716 298726
rect 255320 289876 255372 289882
rect 255320 289818 255372 289824
rect 254676 284980 254728 284986
rect 254676 284922 254728 284928
rect 254584 284436 254636 284442
rect 254584 284378 254636 284384
rect 254596 261594 254624 284378
rect 254584 261588 254636 261594
rect 254584 261530 254636 261536
rect 254124 256692 254176 256698
rect 254124 256634 254176 256640
rect 254136 256018 254164 256634
rect 254124 256012 254176 256018
rect 254124 255954 254176 255960
rect 254030 213888 254086 213897
rect 254030 213823 254086 213832
rect 254044 213246 254072 213823
rect 254032 213240 254084 213246
rect 254032 213182 254084 213188
rect 255332 171737 255360 289818
rect 255424 240281 255452 311063
rect 255516 281722 255544 314638
rect 255504 281716 255556 281722
rect 255504 281658 255556 281664
rect 255504 281512 255556 281518
rect 255504 281454 255556 281460
rect 255516 260846 255544 281454
rect 255504 260840 255556 260846
rect 255504 260782 255556 260788
rect 255410 240272 255466 240281
rect 255410 240207 255466 240216
rect 255410 179480 255466 179489
rect 255410 179415 255466 179424
rect 255318 171728 255374 171737
rect 255318 171663 255374 171672
rect 254584 171216 254636 171222
rect 254584 171158 254636 171164
rect 253938 139768 253994 139777
rect 253938 139703 253994 139712
rect 254596 133890 254624 171158
rect 255424 139398 255452 179415
rect 255412 139392 255464 139398
rect 255412 139334 255464 139340
rect 254584 133884 254636 133890
rect 254584 133826 254636 133832
rect 253572 132524 253624 132530
rect 253572 132466 253624 132472
rect 253480 117360 253532 117366
rect 253480 117302 253532 117308
rect 253386 109032 253442 109041
rect 253386 108967 253442 108976
rect 253492 87650 253520 117302
rect 253584 116618 253612 132466
rect 254582 126032 254638 126041
rect 254582 125967 254638 125976
rect 253572 116612 253624 116618
rect 253572 116554 253624 116560
rect 253480 87644 253532 87650
rect 253480 87586 253532 87592
rect 253294 65512 253350 65521
rect 253294 65447 253350 65456
rect 254596 55865 254624 125967
rect 254768 124228 254820 124234
rect 254768 124170 254820 124176
rect 254676 99408 254728 99414
rect 254676 99350 254728 99356
rect 254582 55856 254638 55865
rect 254582 55791 254638 55800
rect 254688 51746 254716 99350
rect 254780 79354 254808 124170
rect 255976 102241 256004 349823
rect 256068 291854 256096 369174
rect 256712 306374 256740 377590
rect 258724 375352 258776 375358
rect 258724 375294 258776 375300
rect 258736 356726 258764 375294
rect 259472 364334 259500 377590
rect 261496 375358 261524 377604
rect 262232 377590 263166 377618
rect 264256 377590 264822 377618
rect 266372 377590 266478 377618
rect 261484 375352 261536 375358
rect 261484 375294 261536 375300
rect 260838 367840 260894 367849
rect 260838 367775 260894 367784
rect 259472 364306 259592 364334
rect 259564 359514 259592 364306
rect 259552 359508 259604 359514
rect 259552 359450 259604 359456
rect 258724 356720 258776 356726
rect 258724 356662 258776 356668
rect 258736 354674 258764 356662
rect 258736 354646 258948 354674
rect 258816 340196 258868 340202
rect 258816 340138 258868 340144
rect 258722 329080 258778 329089
rect 258722 329015 258778 329024
rect 257342 313304 257398 313313
rect 257342 313239 257398 313248
rect 256712 306346 256832 306374
rect 256804 300121 256832 306346
rect 256790 300112 256846 300121
rect 256790 300047 256846 300056
rect 256700 297424 256752 297430
rect 256700 297366 256752 297372
rect 256056 291848 256108 291854
rect 256056 291790 256108 291796
rect 256712 258058 256740 297366
rect 256804 266422 256832 300047
rect 257356 277545 257384 313239
rect 258170 301472 258226 301481
rect 258170 301407 258226 301416
rect 257526 283656 257582 283665
rect 257526 283591 257582 283600
rect 257342 277536 257398 277545
rect 257342 277471 257398 277480
rect 257356 276010 257384 277471
rect 257344 276004 257396 276010
rect 257344 275946 257396 275952
rect 256792 266416 256844 266422
rect 256792 266358 256844 266364
rect 257540 264897 257568 283591
rect 257526 264888 257582 264897
rect 257526 264823 257582 264832
rect 258078 264888 258134 264897
rect 258078 264823 258134 264832
rect 257436 264308 257488 264314
rect 257436 264250 257488 264256
rect 256700 258052 256752 258058
rect 256700 257994 256752 258000
rect 256712 256766 256740 257994
rect 256700 256760 256752 256766
rect 256700 256702 256752 256708
rect 257344 246424 257396 246430
rect 257344 246366 257396 246372
rect 257356 174321 257384 246366
rect 257448 231169 257476 264250
rect 257528 255332 257580 255338
rect 257528 255274 257580 255280
rect 257540 239970 257568 255274
rect 257528 239964 257580 239970
rect 257528 239906 257580 239912
rect 257434 231160 257490 231169
rect 257434 231095 257490 231104
rect 257448 184210 257476 231095
rect 257436 184204 257488 184210
rect 257436 184146 257488 184152
rect 258092 179382 258120 264823
rect 258184 256086 258212 301407
rect 258172 256080 258224 256086
rect 258172 256022 258224 256028
rect 258184 254590 258212 256022
rect 258172 254584 258224 254590
rect 258172 254526 258224 254532
rect 258736 243545 258764 329015
rect 258828 264761 258856 340138
rect 258920 289882 258948 354646
rect 259092 340876 259144 340882
rect 259092 340818 259144 340824
rect 259104 340202 259132 340818
rect 259092 340196 259144 340202
rect 259092 340138 259144 340144
rect 259458 322144 259514 322153
rect 259458 322079 259514 322088
rect 258908 289876 258960 289882
rect 258908 289818 258960 289824
rect 258920 289134 258948 289818
rect 258908 289128 258960 289134
rect 258908 289070 258960 289076
rect 258906 288688 258962 288697
rect 258906 288623 258962 288632
rect 258814 264752 258870 264761
rect 258814 264687 258870 264696
rect 258920 262274 258948 288623
rect 259366 264752 259422 264761
rect 259366 264687 259422 264696
rect 259380 264246 259408 264687
rect 259368 264240 259420 264246
rect 259368 264182 259420 264188
rect 258908 262268 258960 262274
rect 258908 262210 258960 262216
rect 258920 258074 258948 262210
rect 258828 258046 258948 258074
rect 258722 243536 258778 243545
rect 258722 243471 258778 243480
rect 258828 234433 258856 258046
rect 259368 238128 259420 238134
rect 259368 238070 259420 238076
rect 259380 237969 259408 238070
rect 259366 237960 259422 237969
rect 259366 237895 259422 237904
rect 258814 234424 258870 234433
rect 258814 234359 258870 234368
rect 258080 179376 258132 179382
rect 258080 179318 258132 179324
rect 259276 179376 259328 179382
rect 259276 179318 259328 179324
rect 259288 178673 259316 179318
rect 259274 178664 259330 178673
rect 259274 178599 259330 178608
rect 257342 174312 257398 174321
rect 257342 174247 257398 174256
rect 258722 169824 258778 169833
rect 258722 169759 258778 169768
rect 257344 164348 257396 164354
rect 257344 164290 257396 164296
rect 256148 162172 256200 162178
rect 256148 162114 256200 162120
rect 256056 129804 256108 129810
rect 256056 129746 256108 129752
rect 255962 102232 256018 102241
rect 255962 102167 256018 102176
rect 255964 100768 256016 100774
rect 255964 100710 256016 100716
rect 254768 79348 254820 79354
rect 254768 79290 254820 79296
rect 255976 72457 256004 100710
rect 255962 72448 256018 72457
rect 255962 72383 256018 72392
rect 256068 66881 256096 129746
rect 256160 122806 256188 162114
rect 256700 131776 256752 131782
rect 256700 131718 256752 131724
rect 256712 126274 256740 131718
rect 257356 127673 257384 164290
rect 257620 142180 257672 142186
rect 257620 142122 257672 142128
rect 257528 128444 257580 128450
rect 257528 128386 257580 128392
rect 257342 127664 257398 127673
rect 257342 127599 257398 127608
rect 256700 126268 256752 126274
rect 256700 126210 256752 126216
rect 257436 125656 257488 125662
rect 257436 125598 257488 125604
rect 256148 122800 256200 122806
rect 256148 122742 256200 122748
rect 256240 110560 256292 110566
rect 256240 110502 256292 110508
rect 256148 102808 256200 102814
rect 256148 102750 256200 102756
rect 256054 66872 256110 66881
rect 256054 66807 256110 66816
rect 254676 51740 254728 51746
rect 254676 51682 254728 51688
rect 256160 48929 256188 102750
rect 256252 76809 256280 110502
rect 257342 102232 257398 102241
rect 257342 102167 257398 102176
rect 256238 76800 256294 76809
rect 256238 76735 256294 76744
rect 256146 48920 256202 48929
rect 256146 48855 256202 48864
rect 257356 44878 257384 102167
rect 257448 73953 257476 125598
rect 257540 86193 257568 128386
rect 257632 102066 257660 142122
rect 258736 132433 258764 169759
rect 258814 142624 258870 142633
rect 258814 142559 258870 142568
rect 258722 132424 258778 132433
rect 258722 132359 258778 132368
rect 258724 118788 258776 118794
rect 258724 118730 258776 118736
rect 258078 109712 258134 109721
rect 258078 109647 258134 109656
rect 258092 109313 258120 109647
rect 258078 109304 258134 109313
rect 258078 109239 258134 109248
rect 257620 102060 257672 102066
rect 257620 102002 257672 102008
rect 257526 86184 257582 86193
rect 257526 86119 257582 86128
rect 257434 73944 257490 73953
rect 257434 73879 257490 73888
rect 258736 46238 258764 118730
rect 258828 100706 258856 142559
rect 258906 130248 258962 130257
rect 258906 130183 258962 130192
rect 258920 119406 258948 130183
rect 258908 119400 258960 119406
rect 258908 119342 258960 119348
rect 258906 107128 258962 107137
rect 258906 107063 258962 107072
rect 258816 100700 258868 100706
rect 258816 100642 258868 100648
rect 258816 92540 258868 92546
rect 258816 92482 258868 92488
rect 258828 82142 258856 92482
rect 258816 82136 258868 82142
rect 258816 82078 258868 82084
rect 258920 65657 258948 107063
rect 259380 95198 259408 237895
rect 259472 211138 259500 322079
rect 259564 288250 259592 359450
rect 259644 322312 259696 322318
rect 259644 322254 259696 322260
rect 259552 288244 259604 288250
rect 259552 288186 259604 288192
rect 259656 267714 259684 322254
rect 259736 294024 259788 294030
rect 259736 293966 259788 293972
rect 259644 267708 259696 267714
rect 259644 267650 259696 267656
rect 259656 267034 259684 267650
rect 259644 267028 259696 267034
rect 259644 266970 259696 266976
rect 259748 245857 259776 293966
rect 260104 288244 260156 288250
rect 260104 288186 260156 288192
rect 260116 287162 260144 288186
rect 260104 287156 260156 287162
rect 260104 287098 260156 287104
rect 260116 269822 260144 287098
rect 260104 269816 260156 269822
rect 260104 269758 260156 269764
rect 260104 256760 260156 256766
rect 260104 256702 260156 256708
rect 259734 245848 259790 245857
rect 259734 245783 259790 245792
rect 259460 211132 259512 211138
rect 259460 211074 259512 211080
rect 260116 180198 260144 256702
rect 260746 245848 260802 245857
rect 260746 245783 260802 245792
rect 260760 245002 260788 245783
rect 260748 244996 260800 245002
rect 260748 244938 260800 244944
rect 260748 211132 260800 211138
rect 260748 211074 260800 211080
rect 260760 210458 260788 211074
rect 260748 210452 260800 210458
rect 260748 210394 260800 210400
rect 260852 196761 260880 367775
rect 261484 342916 261536 342922
rect 261484 342858 261536 342864
rect 260930 291408 260986 291417
rect 260930 291343 260986 291352
rect 260944 259418 260972 291343
rect 261496 266393 261524 342858
rect 262126 312624 262182 312633
rect 262126 312559 262182 312568
rect 262140 309806 262168 312559
rect 262128 309800 262180 309806
rect 262128 309742 262180 309748
rect 262232 301617 262260 377590
rect 264256 374105 264284 377590
rect 264242 374096 264298 374105
rect 264242 374031 264298 374040
rect 262864 370524 262916 370530
rect 262864 370466 262916 370472
rect 262310 331800 262366 331809
rect 262310 331735 262366 331744
rect 262218 301608 262274 301617
rect 262218 301543 262274 301552
rect 261576 284980 261628 284986
rect 261576 284922 261628 284928
rect 261482 266384 261538 266393
rect 261482 266319 261538 266328
rect 261496 263537 261524 266319
rect 261482 263528 261538 263537
rect 261482 263463 261538 263472
rect 260932 259412 260984 259418
rect 260932 259354 260984 259360
rect 261588 237969 261616 284922
rect 262128 259412 262180 259418
rect 262128 259354 262180 259360
rect 262140 258806 262168 259354
rect 262128 258800 262180 258806
rect 262128 258742 262180 258748
rect 262128 243432 262180 243438
rect 262128 243374 262180 243380
rect 262140 243030 262168 243374
rect 262128 243024 262180 243030
rect 262128 242966 262180 242972
rect 261574 237960 261630 237969
rect 261574 237895 261630 237904
rect 260838 196752 260894 196761
rect 260838 196687 260894 196696
rect 260104 180192 260156 180198
rect 260104 180134 260156 180140
rect 262140 178702 262168 242966
rect 262324 231169 262352 331735
rect 262876 317422 262904 370466
rect 263690 351112 263746 351121
rect 263690 351047 263746 351056
rect 262404 317416 262456 317422
rect 262404 317358 262456 317364
rect 262864 317416 262916 317422
rect 262864 317358 262916 317364
rect 262416 316130 262444 317358
rect 262404 316124 262456 316130
rect 262404 316066 262456 316072
rect 262416 243438 262444 316066
rect 262956 301572 263008 301578
rect 262956 301514 263008 301520
rect 262862 292768 262918 292777
rect 262862 292703 262918 292712
rect 262770 247072 262826 247081
rect 262770 247007 262826 247016
rect 262404 243432 262456 243438
rect 262404 243374 262456 243380
rect 262784 242962 262812 247007
rect 262772 242956 262824 242962
rect 262772 242898 262824 242904
rect 262310 231160 262366 231169
rect 262310 231095 262366 231104
rect 262876 180130 262904 292703
rect 262968 238134 262996 301514
rect 263600 282940 263652 282946
rect 263600 282882 263652 282888
rect 263612 282849 263640 282882
rect 263598 282840 263654 282849
rect 263598 282775 263654 282784
rect 263600 282192 263652 282198
rect 263600 282134 263652 282140
rect 262956 238128 263008 238134
rect 262956 238070 263008 238076
rect 262864 180124 262916 180130
rect 262864 180066 262916 180072
rect 262128 178696 262180 178702
rect 262128 178638 262180 178644
rect 261482 174448 261538 174457
rect 261482 174383 261538 174392
rect 260102 170232 260158 170241
rect 260102 170167 260158 170176
rect 260116 131102 260144 170167
rect 260286 159080 260342 159089
rect 260286 159015 260342 159024
rect 260196 133952 260248 133958
rect 260196 133894 260248 133900
rect 260104 131096 260156 131102
rect 260104 131038 260156 131044
rect 260104 120216 260156 120222
rect 260104 120158 260156 120164
rect 259368 95192 259420 95198
rect 259368 95134 259420 95140
rect 258906 65648 258962 65657
rect 258906 65583 258962 65592
rect 259460 57316 259512 57322
rect 259460 57258 259512 57264
rect 258724 46232 258776 46238
rect 258724 46174 258776 46180
rect 253204 44872 253256 44878
rect 253204 44814 253256 44820
rect 257344 44872 257396 44878
rect 257344 44814 257396 44820
rect 252560 31068 252612 31074
rect 252560 31010 252612 31016
rect 252572 30297 252600 31010
rect 252558 30288 252614 30297
rect 252558 30223 252614 30232
rect 251916 21412 251968 21418
rect 251916 21354 251968 21360
rect 251928 9489 251956 21354
rect 252572 16574 252600 30223
rect 255964 22840 256016 22846
rect 255964 22782 256016 22788
rect 255976 16574 256004 22782
rect 252572 16546 253520 16574
rect 251914 9480 251970 9489
rect 251914 9415 251970 9424
rect 251822 3632 251878 3641
rect 251822 3567 251878 3576
rect 251928 3534 251956 9415
rect 252374 3632 252430 3641
rect 252374 3567 252430 3576
rect 251180 3528 251232 3534
rect 251180 3470 251232 3476
rect 251916 3528 251968 3534
rect 251916 3470 251968 3476
rect 251192 480 251220 3470
rect 252388 480 252416 3567
rect 253492 480 253520 16546
rect 255884 16546 256004 16574
rect 255884 15162 255912 16546
rect 255872 15156 255924 15162
rect 255872 15098 255924 15104
rect 254676 3800 254728 3806
rect 254676 3742 254728 3748
rect 254688 480 254716 3742
rect 255884 480 255912 15098
rect 257356 9654 257384 44814
rect 258080 39364 258132 39370
rect 258080 39306 258132 39312
rect 257436 21412 257488 21418
rect 257436 21354 257488 21360
rect 257344 9648 257396 9654
rect 257344 9590 257396 9596
rect 257448 6914 257476 21354
rect 257080 6886 257476 6914
rect 257080 3466 257108 6886
rect 258092 3806 258120 39306
rect 258724 9648 258776 9654
rect 258724 9590 258776 9596
rect 258080 3800 258132 3806
rect 258080 3742 258132 3748
rect 258736 3534 258764 9590
rect 258264 3528 258316 3534
rect 258264 3470 258316 3476
rect 258724 3528 258776 3534
rect 258724 3470 258776 3476
rect 257068 3460 257120 3466
rect 257068 3402 257120 3408
rect 257080 480 257108 3402
rect 258276 480 258304 3470
rect 259472 480 259500 57258
rect 260116 32502 260144 120158
rect 260208 69601 260236 133894
rect 260300 121446 260328 159015
rect 261496 142769 261524 174383
rect 262126 167240 262182 167249
rect 262126 167175 262182 167184
rect 261482 142760 261538 142769
rect 261482 142695 261538 142704
rect 261666 140856 261722 140865
rect 261666 140791 261722 140800
rect 261484 127084 261536 127090
rect 261484 127026 261536 127032
rect 260380 126268 260432 126274
rect 260380 126210 260432 126216
rect 260288 121440 260340 121446
rect 260288 121382 260340 121388
rect 260288 109064 260340 109070
rect 260288 109006 260340 109012
rect 260194 69592 260250 69601
rect 260194 69527 260250 69536
rect 260300 57254 260328 109006
rect 260392 92546 260420 126210
rect 260380 92540 260432 92546
rect 260380 92482 260432 92488
rect 260288 57248 260340 57254
rect 260288 57190 260340 57196
rect 260104 32496 260156 32502
rect 260104 32438 260156 32444
rect 259552 22840 259604 22846
rect 259552 22782 259604 22788
rect 259564 19417 259592 22782
rect 261496 22778 261524 127026
rect 261576 111852 261628 111858
rect 261576 111794 261628 111800
rect 261588 72486 261616 111794
rect 261680 101561 261708 140791
rect 261666 101552 261722 101561
rect 261666 101487 261722 101496
rect 261668 98048 261720 98054
rect 261668 97990 261720 97996
rect 261680 79393 261708 97990
rect 262140 93226 262168 167175
rect 262956 167136 263008 167142
rect 262956 167078 263008 167084
rect 262862 163296 262918 163305
rect 262862 163231 262918 163240
rect 262876 122777 262904 163231
rect 262968 160750 262996 167078
rect 263612 163441 263640 282134
rect 263704 252550 263732 351047
rect 264256 344321 264284 374031
rect 266372 365022 266400 377590
rect 267648 374128 267700 374134
rect 267648 374070 267700 374076
rect 267004 374060 267056 374066
rect 267004 374002 267056 374008
rect 266360 365016 266412 365022
rect 266360 364958 266412 364964
rect 265624 364404 265676 364410
rect 265624 364346 265676 364352
rect 264336 360256 264388 360262
rect 264336 360198 264388 360204
rect 264242 344312 264298 344321
rect 264242 344247 264298 344256
rect 264348 343602 264376 360198
rect 265636 354686 265664 364346
rect 265624 354680 265676 354686
rect 265624 354622 265676 354628
rect 264336 343596 264388 343602
rect 264336 343538 264388 343544
rect 264348 342854 264376 343538
rect 264336 342848 264388 342854
rect 264336 342790 264388 342796
rect 264888 342848 264940 342854
rect 264888 342790 264940 342796
rect 264242 318880 264298 318889
rect 264242 318815 264298 318824
rect 263784 291848 263836 291854
rect 263784 291790 263836 291796
rect 263692 252544 263744 252550
rect 263692 252486 263744 252492
rect 263704 251870 263732 252486
rect 263692 251864 263744 251870
rect 263692 251806 263744 251812
rect 263796 219366 263824 291790
rect 263784 219360 263836 219366
rect 263784 219302 263836 219308
rect 263796 218657 263824 219302
rect 263782 218648 263838 218657
rect 263782 218583 263838 218592
rect 264256 189786 264284 318815
rect 264900 282946 264928 342790
rect 264980 337476 265032 337482
rect 264980 337418 265032 337424
rect 264888 282940 264940 282946
rect 264888 282882 264940 282888
rect 264992 206961 265020 337418
rect 264978 206952 265034 206961
rect 264978 206887 265034 206896
rect 264992 206310 265020 206887
rect 264980 206304 265032 206310
rect 264980 206246 265032 206252
rect 264244 189780 264296 189786
rect 264244 189722 264296 189728
rect 264978 175672 265034 175681
rect 264978 175607 265034 175616
rect 264992 175302 265020 175607
rect 264980 175296 265032 175302
rect 264980 175238 265032 175244
rect 265070 175264 265126 175273
rect 265070 175199 265126 175208
rect 264978 174856 265034 174865
rect 264978 174791 265034 174800
rect 264992 174010 265020 174791
rect 264980 174004 265032 174010
rect 264980 173946 265032 173952
rect 265084 173942 265112 175199
rect 265254 174040 265310 174049
rect 265254 173975 265310 173984
rect 265072 173936 265124 173942
rect 265072 173878 265124 173884
rect 265070 173632 265126 173641
rect 265070 173567 265126 173576
rect 264978 172680 265034 172689
rect 265084 172650 265112 173567
rect 264978 172615 265034 172624
rect 265072 172644 265124 172650
rect 264992 172582 265020 172615
rect 265072 172586 265124 172592
rect 264980 172576 265032 172582
rect 264980 172518 265032 172524
rect 265268 172417 265296 173975
rect 264242 172408 264298 172417
rect 264242 172343 264298 172352
rect 265254 172408 265310 172417
rect 265254 172343 265310 172352
rect 263598 163432 263654 163441
rect 263598 163367 263654 163376
rect 262956 160744 263008 160750
rect 262956 160686 263008 160692
rect 263048 160200 263100 160206
rect 263048 160142 263100 160148
rect 263060 151162 263088 160142
rect 263048 151156 263100 151162
rect 263048 151098 263100 151104
rect 262956 150476 263008 150482
rect 262956 150418 263008 150424
rect 262862 122768 262918 122777
rect 262862 122703 262918 122712
rect 262772 120148 262824 120154
rect 262772 120090 262824 120096
rect 262784 113174 262812 120090
rect 262862 116920 262918 116929
rect 262862 116855 262918 116864
rect 262876 116113 262904 116855
rect 262862 116104 262918 116113
rect 262862 116039 262918 116048
rect 262784 113146 262904 113174
rect 262772 100836 262824 100842
rect 262772 100778 262824 100784
rect 262784 95946 262812 100778
rect 262772 95940 262824 95946
rect 262772 95882 262824 95888
rect 262128 93220 262180 93226
rect 262128 93162 262180 93168
rect 261666 79384 261722 79393
rect 261666 79319 261722 79328
rect 261576 72480 261628 72486
rect 261576 72422 261628 72428
rect 262876 31142 262904 113146
rect 262968 110430 262996 150418
rect 263048 146396 263100 146402
rect 263048 146338 263100 146344
rect 262956 110424 263008 110430
rect 262956 110366 263008 110372
rect 263060 107574 263088 146338
rect 263140 138100 263192 138106
rect 263140 138042 263192 138048
rect 263152 126274 263180 138042
rect 264256 135153 264284 172343
rect 265070 172272 265126 172281
rect 265070 172207 265126 172216
rect 264978 171456 265034 171465
rect 264978 171391 265034 171400
rect 264992 171154 265020 171391
rect 265084 171222 265112 172207
rect 265162 171864 265218 171873
rect 265162 171799 265218 171808
rect 265072 171216 265124 171222
rect 265072 171158 265124 171164
rect 264980 171148 265032 171154
rect 264980 171090 265032 171096
rect 265070 171048 265126 171057
rect 265070 170983 265126 170992
rect 264978 170096 265034 170105
rect 264978 170031 265034 170040
rect 264992 169862 265020 170031
rect 264980 169856 265032 169862
rect 264980 169798 265032 169804
rect 265084 169794 265112 170983
rect 265176 169833 265204 171799
rect 265162 169824 265218 169833
rect 265072 169788 265124 169794
rect 265162 169759 265218 169768
rect 265072 169730 265124 169736
rect 265070 169688 265126 169697
rect 265070 169623 265126 169632
rect 264978 168872 265034 168881
rect 264978 168807 265034 168816
rect 264992 168502 265020 168807
rect 264980 168496 265032 168502
rect 264980 168438 265032 168444
rect 265084 168434 265112 169623
rect 265438 168464 265494 168473
rect 265072 168428 265124 168434
rect 265438 168399 265494 168408
rect 265072 168370 265124 168376
rect 265346 167920 265402 167929
rect 265346 167855 265402 167864
rect 264978 167512 265034 167521
rect 264978 167447 265034 167456
rect 264992 167074 265020 167447
rect 265360 167142 265388 167855
rect 265348 167136 265400 167142
rect 265348 167078 265400 167084
rect 264980 167068 265032 167074
rect 264980 167010 265032 167016
rect 265070 166696 265126 166705
rect 265070 166631 265126 166640
rect 264978 166288 265034 166297
rect 264978 166223 265034 166232
rect 264992 165646 265020 166223
rect 265084 165714 265112 166631
rect 265162 165880 265218 165889
rect 265162 165815 265218 165824
rect 265072 165708 265124 165714
rect 265072 165650 265124 165656
rect 264980 165640 265032 165646
rect 264980 165582 265032 165588
rect 265070 165336 265126 165345
rect 265070 165271 265126 165280
rect 264978 164520 265034 164529
rect 264978 164455 265034 164464
rect 264992 164354 265020 164455
rect 264980 164348 265032 164354
rect 264980 164290 265032 164296
rect 265084 164286 265112 165271
rect 265176 164937 265204 165815
rect 265162 164928 265218 164937
rect 265162 164863 265218 164872
rect 265072 164280 265124 164286
rect 265072 164222 265124 164228
rect 265254 164112 265310 164121
rect 265254 164047 265310 164056
rect 265070 163704 265126 163713
rect 265070 163639 265126 163648
rect 265084 162926 265112 163639
rect 265072 162920 265124 162926
rect 264978 162888 265034 162897
rect 265072 162862 265124 162868
rect 264978 162823 265034 162832
rect 264992 162178 265020 162823
rect 265070 162344 265126 162353
rect 265070 162279 265126 162288
rect 264980 162172 265032 162178
rect 264980 162114 265032 162120
rect 265084 161498 265112 162279
rect 265162 161528 265218 161537
rect 265072 161492 265124 161498
rect 265162 161463 265218 161472
rect 265072 161434 265124 161440
rect 264978 161120 265034 161129
rect 264978 161055 265034 161064
rect 264992 160138 265020 161055
rect 264980 160132 265032 160138
rect 264980 160074 265032 160080
rect 264978 159760 265034 159769
rect 264978 159695 265034 159704
rect 264992 158778 265020 159695
rect 265176 159089 265204 161463
rect 265268 159390 265296 164047
rect 265452 163538 265480 168399
rect 265636 167249 265664 354622
rect 267016 305697 267044 374002
rect 267096 306400 267148 306406
rect 267096 306342 267148 306348
rect 267002 305688 267058 305697
rect 267002 305623 267058 305632
rect 265714 290456 265770 290465
rect 265714 290391 265770 290400
rect 265728 249082 265756 290391
rect 267004 285728 267056 285734
rect 267004 285670 267056 285676
rect 265716 249076 265768 249082
rect 265716 249018 265768 249024
rect 266360 231124 266412 231130
rect 266360 231066 266412 231072
rect 266372 229838 266400 231066
rect 266360 229832 266412 229838
rect 266360 229774 266412 229780
rect 267016 185638 267044 285670
rect 267108 218754 267136 306342
rect 267186 299568 267242 299577
rect 267186 299503 267242 299512
rect 267200 274038 267228 299503
rect 267188 274032 267240 274038
rect 267188 273974 267240 273980
rect 267660 234598 267688 374070
rect 268120 374066 268148 377604
rect 269776 374134 269804 377604
rect 270512 377590 271446 377618
rect 272720 377590 273102 377618
rect 269856 375352 269908 375358
rect 269856 375294 269908 375300
rect 269764 374128 269816 374134
rect 269764 374070 269816 374076
rect 268108 374060 268160 374066
rect 268108 374002 268160 374008
rect 269764 357468 269816 357474
rect 269764 357410 269816 357416
rect 269120 325712 269172 325718
rect 269120 325654 269172 325660
rect 267738 320784 267794 320793
rect 267738 320719 267794 320728
rect 267648 234592 267700 234598
rect 267648 234534 267700 234540
rect 267752 222057 267780 320719
rect 267832 305108 267884 305114
rect 267832 305050 267884 305056
rect 267844 253910 267872 305050
rect 268382 284200 268438 284209
rect 268382 284135 268438 284144
rect 268396 276010 268424 284135
rect 268384 276004 268436 276010
rect 268384 275946 268436 275952
rect 267832 253904 267884 253910
rect 267832 253846 267884 253852
rect 267832 247104 267884 247110
rect 267832 247046 267884 247052
rect 267738 222048 267794 222057
rect 267738 221983 267794 221992
rect 267844 219201 267872 247046
rect 268396 227730 268424 275946
rect 269028 253904 269080 253910
rect 269028 253846 269080 253852
rect 269040 253230 269068 253846
rect 269028 253224 269080 253230
rect 269028 253166 269080 253172
rect 269132 246430 269160 325654
rect 269120 246424 269172 246430
rect 269120 246366 269172 246372
rect 269776 235929 269804 357410
rect 269868 345710 269896 375294
rect 270408 358080 270460 358086
rect 270408 358022 270460 358028
rect 270420 357474 270448 358022
rect 270408 357468 270460 357474
rect 270408 357410 270460 357416
rect 270408 352572 270460 352578
rect 270408 352514 270460 352520
rect 270420 352073 270448 352514
rect 270406 352064 270462 352073
rect 270406 351999 270462 352008
rect 269856 345704 269908 345710
rect 269856 345646 269908 345652
rect 269854 296984 269910 296993
rect 269854 296919 269910 296928
rect 269762 235920 269818 235929
rect 269762 235855 269818 235864
rect 269764 234592 269816 234598
rect 269764 234534 269816 234540
rect 268384 227724 268436 227730
rect 268384 227666 268436 227672
rect 267830 219192 267886 219201
rect 267830 219127 267886 219136
rect 267096 218748 267148 218754
rect 267096 218690 267148 218696
rect 268396 188358 268424 227666
rect 269026 222048 269082 222057
rect 269026 221983 269082 221992
rect 269040 221542 269068 221983
rect 269028 221536 269080 221542
rect 269028 221478 269080 221484
rect 268384 188352 268436 188358
rect 268384 188294 268436 188300
rect 269776 186425 269804 234534
rect 269762 186416 269818 186425
rect 269762 186351 269818 186360
rect 267004 185632 267056 185638
rect 267004 185574 267056 185580
rect 269868 181558 269896 296919
rect 270420 244934 270448 351999
rect 270408 244928 270460 244934
rect 270408 244870 270460 244876
rect 270420 244322 270448 244870
rect 269948 244316 270000 244322
rect 269948 244258 270000 244264
rect 270408 244316 270460 244322
rect 270408 244258 270460 244264
rect 269960 237153 269988 244258
rect 269946 237144 270002 237153
rect 269946 237079 270002 237088
rect 270406 235920 270462 235929
rect 270406 235855 270462 235864
rect 270420 235278 270448 235855
rect 270408 235272 270460 235278
rect 270408 235214 270460 235220
rect 270408 230444 270460 230450
rect 270408 230386 270460 230392
rect 270420 229838 270448 230386
rect 270408 229832 270460 229838
rect 270408 229774 270460 229780
rect 270420 195294 270448 229774
rect 270512 219434 270540 377590
rect 272720 376961 272748 377590
rect 272706 376952 272762 376961
rect 272706 376887 272762 376896
rect 274744 375358 274772 377604
rect 276032 377590 276414 377618
rect 274732 375352 274784 375358
rect 274732 375294 274784 375300
rect 274086 374640 274142 374649
rect 274086 374575 274142 374584
rect 273902 374096 273958 374105
rect 271144 374060 271196 374066
rect 273902 374031 273958 374040
rect 271144 374002 271196 374008
rect 271156 230450 271184 374002
rect 272524 348424 272576 348430
rect 272524 348366 272576 348372
rect 272536 336705 272564 348366
rect 271878 336696 271934 336705
rect 271878 336631 271934 336640
rect 272522 336696 272578 336705
rect 272522 336631 272578 336640
rect 271892 335481 271920 336631
rect 271878 335472 271934 335481
rect 271878 335407 271934 335416
rect 271234 317656 271290 317665
rect 271234 317591 271290 317600
rect 271144 230444 271196 230450
rect 271144 230386 271196 230392
rect 270500 219428 270552 219434
rect 270500 219370 270552 219376
rect 270512 218074 270540 219370
rect 270500 218068 270552 218074
rect 270500 218010 270552 218016
rect 271144 218068 271196 218074
rect 271144 218010 271196 218016
rect 270408 195288 270460 195294
rect 270408 195230 270460 195236
rect 270314 184512 270370 184521
rect 270314 184447 270370 184456
rect 270328 182850 270356 184447
rect 270316 182844 270368 182850
rect 270316 182786 270368 182792
rect 269856 181552 269908 181558
rect 269856 181494 269908 181500
rect 271156 178770 271184 218010
rect 271248 184890 271276 317591
rect 271892 313410 271920 335407
rect 272616 327752 272668 327758
rect 272616 327694 272668 327700
rect 272628 327146 272656 327694
rect 272616 327140 272668 327146
rect 272616 327082 272668 327088
rect 271880 313404 271932 313410
rect 271880 313346 271932 313352
rect 272524 313404 272576 313410
rect 272524 313346 272576 313352
rect 272430 266384 272486 266393
rect 272430 266319 272486 266328
rect 272444 262857 272472 266319
rect 272430 262848 272486 262857
rect 272430 262783 272486 262792
rect 272432 184952 272484 184958
rect 272432 184894 272484 184900
rect 271236 184884 271288 184890
rect 271236 184826 271288 184832
rect 272444 182170 272472 184894
rect 272432 182164 272484 182170
rect 272432 182106 272484 182112
rect 271144 178764 271196 178770
rect 271144 178706 271196 178712
rect 272536 177585 272564 313346
rect 272628 216617 272656 327082
rect 273168 295452 273220 295458
rect 273168 295394 273220 295400
rect 273180 238882 273208 295394
rect 273916 257446 273944 374031
rect 274100 339561 274128 374575
rect 274640 365016 274692 365022
rect 274640 364958 274692 364964
rect 274086 339552 274142 339561
rect 274086 339487 274142 339496
rect 274100 335354 274128 339487
rect 274008 335326 274128 335354
rect 274008 322250 274036 335326
rect 273996 322244 274048 322250
rect 273996 322186 274048 322192
rect 273994 306640 274050 306649
rect 273994 306575 274050 306584
rect 273904 257440 273956 257446
rect 273904 257382 273956 257388
rect 273168 238876 273220 238882
rect 273168 238818 273220 238824
rect 273180 238746 273208 238818
rect 273168 238740 273220 238746
rect 273168 238682 273220 238688
rect 273904 221468 273956 221474
rect 273904 221410 273956 221416
rect 272708 220108 272760 220114
rect 272708 220050 272760 220056
rect 272614 216608 272670 216617
rect 272614 216543 272670 216552
rect 272628 215393 272656 216543
rect 272614 215384 272670 215393
rect 272614 215319 272670 215328
rect 272720 209098 272748 220050
rect 272708 209092 272760 209098
rect 272708 209034 272760 209040
rect 273916 181490 273944 221410
rect 274008 201822 274036 306575
rect 274088 302320 274140 302326
rect 274088 302262 274140 302268
rect 274100 246430 274128 302262
rect 274088 246424 274140 246430
rect 274088 246366 274140 246372
rect 274086 215384 274142 215393
rect 274086 215319 274142 215328
rect 273996 201816 274048 201822
rect 273996 201758 274048 201764
rect 273904 181484 273956 181490
rect 273904 181426 273956 181432
rect 274100 180169 274128 215319
rect 274652 211070 274680 364958
rect 275282 303784 275338 303793
rect 275282 303719 275338 303728
rect 274640 211064 274692 211070
rect 274640 211006 274692 211012
rect 274652 210526 274680 211006
rect 274640 210520 274692 210526
rect 274640 210462 274692 210468
rect 274086 180160 274142 180169
rect 274086 180095 274142 180104
rect 274638 178664 274694 178673
rect 274638 178599 274694 178608
rect 272522 177576 272578 177585
rect 272522 177511 272578 177520
rect 274652 177313 274680 178599
rect 275296 178129 275324 303719
rect 276032 227662 276060 377590
rect 278056 374066 278084 377604
rect 279516 375352 279568 375358
rect 279516 375294 279568 375300
rect 278228 375148 278280 375154
rect 278228 375090 278280 375096
rect 278044 374060 278096 374066
rect 278044 374002 278096 374008
rect 276664 324352 276716 324358
rect 276664 324294 276716 324300
rect 276020 227656 276072 227662
rect 276020 227598 276072 227604
rect 276032 227050 276060 227598
rect 276020 227044 276072 227050
rect 276020 226986 276072 226992
rect 275376 218748 275428 218754
rect 275376 218690 275428 218696
rect 275388 190454 275416 218690
rect 275388 190426 275508 190454
rect 275282 178120 275338 178129
rect 275282 178055 275338 178064
rect 275480 178022 275508 190426
rect 276676 178809 276704 324294
rect 278042 296848 278098 296857
rect 278042 296783 278098 296792
rect 276754 295488 276810 295497
rect 276754 295423 276810 295432
rect 276768 265674 276796 295423
rect 277398 267064 277454 267073
rect 277398 266999 277454 267008
rect 276756 265668 276808 265674
rect 276756 265610 276808 265616
rect 277412 220862 277440 266999
rect 276756 220856 276808 220862
rect 276756 220798 276808 220804
rect 277400 220856 277452 220862
rect 277400 220798 277452 220804
rect 276768 211041 276796 220798
rect 276754 211032 276810 211041
rect 276754 210967 276810 210976
rect 276662 178800 276718 178809
rect 276662 178735 276718 178744
rect 275468 178016 275520 178022
rect 275468 177958 275520 177964
rect 276768 177342 276796 210967
rect 278056 186425 278084 296783
rect 278240 295458 278268 375090
rect 279424 309188 279476 309194
rect 279424 309130 279476 309136
rect 278228 295452 278280 295458
rect 278228 295394 278280 295400
rect 278134 295352 278190 295361
rect 278134 295287 278190 295296
rect 278042 186416 278098 186425
rect 278042 186351 278098 186360
rect 278148 185745 278176 295287
rect 279056 280628 279108 280634
rect 279056 280570 279108 280576
rect 278228 201816 278280 201822
rect 278228 201758 278280 201764
rect 278134 185736 278190 185745
rect 278134 185671 278190 185680
rect 276756 177336 276808 177342
rect 274638 177304 274694 177313
rect 276756 177278 276808 177284
rect 274638 177239 274694 177248
rect 278240 175846 278268 201758
rect 278318 189952 278374 189961
rect 278318 189887 278374 189896
rect 278332 178673 278360 189887
rect 278318 178664 278374 178673
rect 278318 178599 278374 178608
rect 278228 175840 278280 175846
rect 278228 175782 278280 175788
rect 279068 170490 279096 280570
rect 279436 194585 279464 309130
rect 279528 298761 279556 375294
rect 279712 375154 279740 377604
rect 281368 376825 281396 377604
rect 283038 377590 283604 377618
rect 281354 376816 281410 376825
rect 281354 376751 281410 376760
rect 280158 376680 280214 376689
rect 280158 376615 280214 376624
rect 280172 375358 280200 376615
rect 280160 375352 280212 375358
rect 280160 375294 280212 375300
rect 279700 375148 279752 375154
rect 279700 375090 279752 375096
rect 283576 359553 283604 377590
rect 284312 377590 284694 377618
rect 285692 377590 286350 377618
rect 283562 359544 283618 359553
rect 282184 359508 282236 359514
rect 283562 359479 283618 359488
rect 282184 359450 282236 359456
rect 280894 338736 280950 338745
rect 280894 338671 280950 338680
rect 280804 322992 280856 322998
rect 280804 322934 280856 322940
rect 279514 298752 279570 298761
rect 279514 298687 279570 298696
rect 280160 225684 280212 225690
rect 280160 225626 280212 225632
rect 279422 194576 279478 194585
rect 279422 194511 279478 194520
rect 279148 185632 279200 185638
rect 279148 185574 279200 185580
rect 279160 173894 279188 185574
rect 279608 184884 279660 184890
rect 279608 184826 279660 184832
rect 279620 178129 279648 184826
rect 279974 178800 280030 178809
rect 279974 178735 280030 178744
rect 279606 178120 279662 178129
rect 279606 178055 279662 178064
rect 279988 176654 280016 178735
rect 279988 176626 280108 176654
rect 279332 175840 279384 175846
rect 279332 175782 279384 175788
rect 279422 175808 279478 175817
rect 279160 173866 279280 173894
rect 279252 173618 279280 173866
rect 279344 173777 279372 175782
rect 279422 175743 279478 175752
rect 279330 173768 279386 173777
rect 279330 173703 279386 173712
rect 279252 173590 279372 173618
rect 279344 170762 279372 173590
rect 279436 172281 279464 175743
rect 279422 172272 279478 172281
rect 279422 172207 279478 172216
rect 280080 171057 280108 176626
rect 280066 171048 280122 171057
rect 280066 170983 280122 170992
rect 280068 170944 280120 170950
rect 280068 170886 280120 170892
rect 279344 170734 279464 170762
rect 279330 170504 279386 170513
rect 279068 170462 279330 170490
rect 279330 170439 279386 170448
rect 265622 167240 265678 167249
rect 265622 167175 265678 167184
rect 265622 164928 265678 164937
rect 265622 164863 265678 164872
rect 265440 163532 265492 163538
rect 265440 163474 265492 163480
rect 265438 160304 265494 160313
rect 265438 160239 265494 160248
rect 265452 160206 265480 160239
rect 265440 160200 265492 160206
rect 265440 160142 265492 160148
rect 265256 159384 265308 159390
rect 265256 159326 265308 159332
rect 265162 159080 265218 159089
rect 265162 159015 265218 159024
rect 265162 158944 265218 158953
rect 265162 158879 265218 158888
rect 264980 158772 265032 158778
rect 264980 158714 265032 158720
rect 265070 158536 265126 158545
rect 265070 158471 265126 158480
rect 264978 157720 265034 157729
rect 264978 157655 265034 157664
rect 264992 157486 265020 157655
rect 264980 157480 265032 157486
rect 264980 157422 265032 157428
rect 265084 157418 265112 158471
rect 265072 157412 265124 157418
rect 265072 157354 265124 157360
rect 265070 157176 265126 157185
rect 265070 157111 265126 157120
rect 264978 156768 265034 156777
rect 264978 156703 265034 156712
rect 264992 155990 265020 156703
rect 265084 156058 265112 157111
rect 265176 156641 265204 158879
rect 265162 156632 265218 156641
rect 265162 156567 265218 156576
rect 265162 156360 265218 156369
rect 265162 156295 265218 156304
rect 265072 156052 265124 156058
rect 265072 155994 265124 156000
rect 264980 155984 265032 155990
rect 264980 155926 265032 155932
rect 265070 155952 265126 155961
rect 265070 155887 265126 155896
rect 264978 155544 265034 155553
rect 264978 155479 265034 155488
rect 264992 154698 265020 155479
rect 264980 154692 265032 154698
rect 264980 154634 265032 154640
rect 265084 154630 265112 155887
rect 265072 154624 265124 154630
rect 265072 154566 265124 154572
rect 264978 154184 265034 154193
rect 264978 154119 265034 154128
rect 264426 153504 264482 153513
rect 264426 153439 264482 153448
rect 264242 135144 264298 135153
rect 264242 135079 264298 135088
rect 263140 126268 263192 126274
rect 263140 126210 263192 126216
rect 264334 118144 264390 118153
rect 264334 118079 264390 118088
rect 264242 112024 264298 112033
rect 264242 111959 264298 111968
rect 263048 107568 263100 107574
rect 263048 107510 263100 107516
rect 262956 106344 263008 106350
rect 262956 106286 263008 106292
rect 262968 67017 262996 106286
rect 263324 104984 263376 104990
rect 263324 104926 263376 104932
rect 263048 104168 263100 104174
rect 263048 104110 263100 104116
rect 262954 67008 263010 67017
rect 262954 66943 263010 66952
rect 262956 61464 263008 61470
rect 262956 61406 263008 61412
rect 262864 31136 262916 31142
rect 262864 31078 262916 31084
rect 261484 22772 261536 22778
rect 261484 22714 261536 22720
rect 259550 19408 259606 19417
rect 259550 19343 259606 19352
rect 260102 19408 260158 19417
rect 260102 19343 260158 19352
rect 260116 3505 260144 19343
rect 262968 19281 262996 61406
rect 263060 61402 263088 104110
rect 263336 102814 263364 104926
rect 263324 102808 263376 102814
rect 263324 102750 263376 102756
rect 263048 61396 263100 61402
rect 263048 61338 263100 61344
rect 262218 19272 262274 19281
rect 262218 19207 262274 19216
rect 262954 19272 263010 19281
rect 262954 19207 263010 19216
rect 262232 16574 262260 19207
rect 262232 16546 262536 16574
rect 261760 10328 261812 10334
rect 261758 10296 261760 10305
rect 261812 10296 261814 10305
rect 261758 10231 261814 10240
rect 260102 3496 260158 3505
rect 260102 3431 260158 3440
rect 260654 3496 260710 3505
rect 260654 3431 260710 3440
rect 260668 480 260696 3431
rect 261772 480 261800 10231
rect 262508 490 262536 16546
rect 264256 11762 264284 111959
rect 264348 29646 264376 118079
rect 264440 113150 264468 153439
rect 264992 153270 265020 154119
rect 265176 153785 265204 156295
rect 265162 153776 265218 153785
rect 265162 153711 265218 153720
rect 264980 153264 265032 153270
rect 264980 153206 265032 153212
rect 265070 152960 265126 152969
rect 265070 152895 265126 152904
rect 264978 152552 265034 152561
rect 264978 152487 265034 152496
rect 264992 151842 265020 152487
rect 265084 151910 265112 152895
rect 265072 151904 265124 151910
rect 265072 151846 265124 151852
rect 264980 151836 265032 151842
rect 264980 151778 265032 151784
rect 265346 151600 265402 151609
rect 265346 151535 265402 151544
rect 265070 150784 265126 150793
rect 265070 150719 265126 150728
rect 264978 149968 265034 149977
rect 264978 149903 265034 149912
rect 264992 149122 265020 149903
rect 264980 149116 265032 149122
rect 264980 149058 265032 149064
rect 265084 148345 265112 150719
rect 265360 150482 265388 151535
rect 265348 150476 265400 150482
rect 265348 150418 265400 150424
rect 265636 149734 265664 164863
rect 279436 164234 279464 170734
rect 279160 164206 279464 164234
rect 267278 159352 267334 159361
rect 267278 159287 267334 159296
rect 265714 154592 265770 154601
rect 265714 154527 265770 154536
rect 265728 151094 265756 154527
rect 265806 152008 265862 152017
rect 265806 151943 265862 151952
rect 265716 151088 265768 151094
rect 265716 151030 265768 151036
rect 265624 149728 265676 149734
rect 265624 149670 265676 149676
rect 265622 149016 265678 149025
rect 265622 148951 265678 148960
rect 265162 148608 265218 148617
rect 265162 148543 265218 148552
rect 265070 148336 265126 148345
rect 265070 148271 265126 148280
rect 265070 148200 265126 148209
rect 265070 148135 265126 148144
rect 264978 147792 265034 147801
rect 264978 147727 264980 147736
rect 265032 147727 265034 147736
rect 264980 147698 265032 147704
rect 265084 147694 265112 148135
rect 265072 147688 265124 147694
rect 265072 147630 265124 147636
rect 265070 147384 265126 147393
rect 265070 147319 265126 147328
rect 264978 146432 265034 146441
rect 264978 146367 265034 146376
rect 264992 145761 265020 146367
rect 265084 146334 265112 147319
rect 265176 146402 265204 148543
rect 265164 146396 265216 146402
rect 265164 146338 265216 146344
rect 265072 146328 265124 146334
rect 265072 146270 265124 146276
rect 265162 146024 265218 146033
rect 265162 145959 265218 145968
rect 264978 145752 265034 145761
rect 264978 145687 265034 145696
rect 265070 145616 265126 145625
rect 265070 145551 265126 145560
rect 264978 145208 265034 145217
rect 264978 145143 265034 145152
rect 264992 145042 265020 145143
rect 264980 145036 265032 145042
rect 264980 144978 265032 144984
rect 265084 144974 265112 145551
rect 265072 144968 265124 144974
rect 265072 144910 265124 144916
rect 264978 144800 265034 144809
rect 264978 144735 265034 144744
rect 264610 143848 264666 143857
rect 264610 143783 264666 143792
rect 264520 137284 264572 137290
rect 264520 137226 264572 137232
rect 264428 113144 264480 113150
rect 264428 113086 264480 113092
rect 264426 108624 264482 108633
rect 264426 108559 264482 108568
rect 264440 55894 264468 108559
rect 264532 107642 264560 137226
rect 264624 113801 264652 143783
rect 264992 143614 265020 144735
rect 265176 144226 265204 145959
rect 265254 144392 265310 144401
rect 265254 144327 265310 144336
rect 265164 144220 265216 144226
rect 265164 144162 265216 144168
rect 264980 143608 265032 143614
rect 264980 143550 265032 143556
rect 265070 143440 265126 143449
rect 265070 143375 265126 143384
rect 264980 142860 265032 142866
rect 264980 142802 265032 142808
rect 264992 142225 265020 142802
rect 264978 142216 265034 142225
rect 265084 142186 265112 143375
rect 264978 142151 265034 142160
rect 265072 142180 265124 142186
rect 265268 142154 265296 144327
rect 265072 142122 265124 142128
rect 265176 142126 265296 142154
rect 265176 141438 265204 142126
rect 265164 141432 265216 141438
rect 265164 141374 265216 141380
rect 265254 141264 265310 141273
rect 265254 141199 265310 141208
rect 264978 140040 265034 140049
rect 264978 139975 265034 139984
rect 264992 139466 265020 139975
rect 264980 139460 265032 139466
rect 264980 139402 265032 139408
rect 265070 139224 265126 139233
rect 265070 139159 265126 139168
rect 264978 138272 265034 138281
rect 264978 138207 265034 138216
rect 264992 138038 265020 138207
rect 265084 138106 265112 139159
rect 265072 138100 265124 138106
rect 265072 138042 265124 138048
rect 264980 138032 265032 138038
rect 264980 137974 265032 137980
rect 264978 137864 265034 137873
rect 264978 137799 265034 137808
rect 264992 136678 265020 137799
rect 264980 136672 265032 136678
rect 264980 136614 265032 136620
rect 265070 136640 265126 136649
rect 265070 136575 265126 136584
rect 264978 135688 265034 135697
rect 264978 135623 265034 135632
rect 264992 135318 265020 135623
rect 265084 135386 265112 136575
rect 265072 135380 265124 135386
rect 265072 135322 265124 135328
rect 264980 135312 265032 135318
rect 264980 135254 265032 135260
rect 265070 135280 265126 135289
rect 265070 135215 265126 135224
rect 265084 134473 265112 135215
rect 265162 134872 265218 134881
rect 265162 134807 265218 134816
rect 265070 134464 265126 134473
rect 265070 134399 265126 134408
rect 264978 134056 265034 134065
rect 264978 133991 265034 134000
rect 264992 133958 265020 133991
rect 264980 133952 265032 133958
rect 264980 133894 265032 133900
rect 264978 133648 265034 133657
rect 264978 133583 265034 133592
rect 264992 132530 265020 133583
rect 264980 132524 265032 132530
rect 264980 132466 265032 132472
rect 264978 131880 265034 131889
rect 264978 131815 265034 131824
rect 264992 131170 265020 131815
rect 265176 131782 265204 134807
rect 265268 134570 265296 141199
rect 265636 137290 265664 148951
rect 265714 143032 265770 143041
rect 265714 142967 265770 142976
rect 265624 137284 265676 137290
rect 265624 137226 265676 137232
rect 265256 134564 265308 134570
rect 265256 134506 265308 134512
rect 265622 134192 265678 134201
rect 265622 134127 265678 134136
rect 265164 131776 265216 131782
rect 265164 131718 265216 131724
rect 264980 131164 265032 131170
rect 264980 131106 265032 131112
rect 264978 131064 265034 131073
rect 264978 130999 265034 131008
rect 264992 129810 265020 130999
rect 264980 129804 265032 129810
rect 264980 129746 265032 129752
rect 265070 129296 265126 129305
rect 265070 129231 265126 129240
rect 264978 128888 265034 128897
rect 264978 128823 265034 128832
rect 264992 128382 265020 128823
rect 265084 128450 265112 129231
rect 265072 128444 265124 128450
rect 265072 128386 265124 128392
rect 264980 128376 265032 128382
rect 264980 128318 265032 128324
rect 264978 127936 265034 127945
rect 264978 127871 265034 127880
rect 264992 127022 265020 127871
rect 265070 127528 265126 127537
rect 265070 127463 265126 127472
rect 265084 127090 265112 127463
rect 265072 127084 265124 127090
rect 265072 127026 265124 127032
rect 264980 127016 265032 127022
rect 264980 126958 265032 126964
rect 264978 125896 265034 125905
rect 264978 125831 265034 125840
rect 264992 125662 265020 125831
rect 264980 125656 265032 125662
rect 264980 125598 265032 125604
rect 264978 124536 265034 124545
rect 264978 124471 265034 124480
rect 264992 124234 265020 124471
rect 264980 124228 265032 124234
rect 264980 124170 265032 124176
rect 265070 124128 265126 124137
rect 265070 124063 265126 124072
rect 264980 122936 265032 122942
rect 264978 122904 264980 122913
rect 265032 122904 265034 122913
rect 265084 122874 265112 124063
rect 264978 122839 265034 122848
rect 265072 122868 265124 122874
rect 265072 122810 265124 122816
rect 264978 121952 265034 121961
rect 264978 121887 265034 121896
rect 264992 121514 265020 121887
rect 264980 121508 265032 121514
rect 264980 121450 265032 121456
rect 264978 120728 265034 120737
rect 264978 120663 265034 120672
rect 264992 120154 265020 120663
rect 265070 120320 265126 120329
rect 265070 120255 265126 120264
rect 265084 120222 265112 120255
rect 265072 120216 265124 120222
rect 265072 120158 265124 120164
rect 264980 120148 265032 120154
rect 264980 120090 265032 120096
rect 264978 119368 265034 119377
rect 264978 119303 265034 119312
rect 264992 118726 265020 119303
rect 265070 118960 265126 118969
rect 265070 118895 265126 118904
rect 265084 118794 265112 118895
rect 265072 118788 265124 118794
rect 265072 118730 265124 118736
rect 264980 118720 265032 118726
rect 264980 118662 265032 118668
rect 264978 118552 265034 118561
rect 264978 118487 265034 118496
rect 264992 117366 265020 118487
rect 264980 117360 265032 117366
rect 264980 117302 265032 117308
rect 265162 116784 265218 116793
rect 265162 116719 265218 116728
rect 264980 116000 265032 116006
rect 264978 115968 264980 115977
rect 265032 115968 265034 115977
rect 264978 115903 265034 115912
rect 265070 115152 265126 115161
rect 265070 115087 265126 115096
rect 265084 114646 265112 115087
rect 265072 114640 265124 114646
rect 264978 114608 265034 114617
rect 265072 114582 265124 114588
rect 264978 114543 264980 114552
rect 265032 114543 265034 114552
rect 264980 114514 265032 114520
rect 264978 114200 265034 114209
rect 264978 114135 265034 114144
rect 264610 113792 264666 113801
rect 264610 113727 264666 113736
rect 264992 113218 265020 114135
rect 265176 113937 265204 116719
rect 265162 113928 265218 113937
rect 265162 113863 265218 113872
rect 264980 113212 265032 113218
rect 264980 113154 265032 113160
rect 264978 112568 265034 112577
rect 264978 112503 265034 112512
rect 264992 111858 265020 112503
rect 264980 111852 265032 111858
rect 264980 111794 265032 111800
rect 265070 111616 265126 111625
rect 265070 111551 265126 111560
rect 264978 111208 265034 111217
rect 264978 111143 265034 111152
rect 264992 110566 265020 111143
rect 264980 110560 265032 110566
rect 264980 110502 265032 110508
rect 265084 110498 265112 111551
rect 265072 110492 265124 110498
rect 265072 110434 265124 110440
rect 265070 110392 265126 110401
rect 265070 110327 265126 110336
rect 265084 109070 265112 110327
rect 265072 109064 265124 109070
rect 264978 109032 265034 109041
rect 265072 109006 265124 109012
rect 264978 108967 265034 108976
rect 264992 107710 265020 108967
rect 264980 107704 265032 107710
rect 264980 107646 265032 107652
rect 264520 107636 264572 107642
rect 264520 107578 264572 107584
rect 265254 106992 265310 107001
rect 265254 106927 265310 106936
rect 265268 106350 265296 106927
rect 265256 106344 265308 106350
rect 265256 106286 265308 106292
rect 264978 106040 265034 106049
rect 264978 105975 265034 105984
rect 264992 104922 265020 105975
rect 265162 105632 265218 105641
rect 265162 105567 265218 105576
rect 265176 104990 265204 105567
rect 265164 104984 265216 104990
rect 265164 104926 265216 104932
rect 264980 104916 265032 104922
rect 264980 104858 265032 104864
rect 265070 104816 265126 104825
rect 265070 104751 265126 104760
rect 264978 104408 265034 104417
rect 264978 104343 265034 104352
rect 264518 103864 264574 103873
rect 264518 103799 264574 103808
rect 264532 98666 264560 103799
rect 264992 103562 265020 104343
rect 265084 104174 265112 104751
rect 265072 104168 265124 104174
rect 265072 104110 265124 104116
rect 264980 103556 265032 103562
rect 264980 103498 265032 103504
rect 264978 103456 265034 103465
rect 264978 103391 265034 103400
rect 264992 102202 265020 103391
rect 265070 102640 265126 102649
rect 265070 102575 265126 102584
rect 264980 102196 265032 102202
rect 264980 102138 265032 102144
rect 264978 101280 265034 101289
rect 264978 101215 265034 101224
rect 264992 100774 265020 101215
rect 264980 100768 265032 100774
rect 264980 100710 265032 100716
rect 264978 100056 265034 100065
rect 264978 99991 265034 100000
rect 264992 99414 265020 99991
rect 264980 99408 265032 99414
rect 264980 99350 265032 99356
rect 265084 98977 265112 102575
rect 265162 100872 265218 100881
rect 265162 100807 265164 100816
rect 265216 100807 265218 100816
rect 265164 100778 265216 100784
rect 265070 98968 265126 98977
rect 265070 98903 265126 98912
rect 264978 98696 265034 98705
rect 264520 98660 264572 98666
rect 264978 98631 265034 98640
rect 264520 98602 264572 98608
rect 264992 98054 265020 98631
rect 264980 98048 265032 98054
rect 264980 97990 265032 97996
rect 264978 97880 265034 97889
rect 264978 97815 265034 97824
rect 264518 97472 264574 97481
rect 264518 97407 264574 97416
rect 264532 80753 264560 97407
rect 264992 97306 265020 97815
rect 264980 97300 265032 97306
rect 264980 97242 265032 97248
rect 264518 80744 264574 80753
rect 264518 80679 264574 80688
rect 265636 61441 265664 134127
rect 265728 124914 265756 142967
rect 265820 141506 265848 151943
rect 265808 141500 265860 141506
rect 265808 141442 265860 141448
rect 265806 139632 265862 139641
rect 265806 139567 265862 139576
rect 265716 124908 265768 124914
rect 265716 124850 265768 124856
rect 265714 98288 265770 98297
rect 265714 98223 265770 98232
rect 265622 61432 265678 61441
rect 265622 61367 265678 61376
rect 264428 55888 264480 55894
rect 264428 55830 264480 55836
rect 265728 36582 265756 98223
rect 265820 91769 265848 139567
rect 267094 131472 267150 131481
rect 267094 131407 267150 131416
rect 265898 126304 265954 126313
rect 265898 126239 265954 126248
rect 265912 93158 265940 126239
rect 267002 121544 267058 121553
rect 267002 121479 267058 121488
rect 265900 93152 265952 93158
rect 265900 93094 265952 93100
rect 265806 91760 265862 91769
rect 265806 91695 265862 91704
rect 266360 62824 266412 62830
rect 266360 62766 266412 62772
rect 265716 36576 265768 36582
rect 265716 36518 265768 36524
rect 264336 29640 264388 29646
rect 264336 29582 264388 29588
rect 264336 24132 264388 24138
rect 264336 24074 264388 24080
rect 264348 13802 264376 24074
rect 266372 16574 266400 62766
rect 267016 46306 267044 121479
rect 267108 68241 267136 131407
rect 267186 125352 267242 125361
rect 267186 125287 267242 125296
rect 267200 83609 267228 125287
rect 267292 118658 267320 159287
rect 267280 118652 267332 118658
rect 267280 118594 267332 118600
rect 279160 113174 279188 164206
rect 280080 161474 280108 170886
rect 279252 161446 280108 161474
rect 279252 151814 279280 161446
rect 279252 151786 279372 151814
rect 279344 136921 279372 151786
rect 279330 136912 279386 136921
rect 279330 136847 279386 136856
rect 280172 118425 280200 225626
rect 280816 195362 280844 322934
rect 280908 272542 280936 338671
rect 282196 326369 282224 359450
rect 283564 338768 283616 338774
rect 283564 338710 283616 338716
rect 282182 326360 282238 326369
rect 282182 326295 282238 326304
rect 283576 319462 283604 338710
rect 283564 319456 283616 319462
rect 283564 319398 283616 319404
rect 282920 311908 282972 311914
rect 282920 311850 282972 311856
rect 282932 310457 282960 311850
rect 282918 310448 282974 310457
rect 282918 310383 282974 310392
rect 283562 310448 283618 310457
rect 283562 310383 283618 310392
rect 282184 307896 282236 307902
rect 282184 307838 282236 307844
rect 280988 304360 281040 304366
rect 280988 304302 281040 304308
rect 281000 283014 281028 304302
rect 280988 283008 281040 283014
rect 280988 282950 281040 282956
rect 281724 283008 281776 283014
rect 281724 282950 281776 282956
rect 280896 272536 280948 272542
rect 280896 272478 280948 272484
rect 280896 204944 280948 204950
rect 280896 204886 280948 204892
rect 280804 195356 280856 195362
rect 280804 195298 280856 195304
rect 280434 194032 280490 194041
rect 280434 193967 280490 193976
rect 280252 184204 280304 184210
rect 280252 184146 280304 184152
rect 280158 118416 280214 118425
rect 280158 118351 280214 118360
rect 279160 113146 279464 113174
rect 267278 106448 267334 106457
rect 267278 106383 267334 106392
rect 267186 83600 267242 83609
rect 267186 83535 267242 83544
rect 267292 73817 267320 106383
rect 279330 105768 279386 105777
rect 279330 105703 279386 105712
rect 279344 103514 279372 105703
rect 279436 104961 279464 113146
rect 280264 105505 280292 184146
rect 280344 178696 280396 178702
rect 280344 178638 280396 178644
rect 280356 151881 280384 178638
rect 280448 174729 280476 193967
rect 280908 178702 280936 204886
rect 281632 189780 281684 189786
rect 281632 189722 281684 189728
rect 280896 178696 280948 178702
rect 280896 178638 280948 178644
rect 280804 177336 280856 177342
rect 280804 177278 280856 177284
rect 280434 174720 280490 174729
rect 280434 174655 280490 174664
rect 280342 151872 280398 151881
rect 280342 151807 280398 151816
rect 280342 145072 280398 145081
rect 280342 145007 280398 145016
rect 280250 105496 280306 105505
rect 280250 105431 280306 105440
rect 279422 104952 279478 104961
rect 279422 104887 279478 104896
rect 279068 103486 279372 103514
rect 267830 96656 267886 96665
rect 267830 96591 267886 96600
rect 267738 95840 267794 95849
rect 267738 95775 267794 95784
rect 267752 93838 267780 95775
rect 267844 95130 267872 96591
rect 267832 95124 267884 95130
rect 267832 95066 267884 95072
rect 269120 95124 269172 95130
rect 269120 95066 269172 95072
rect 267740 93832 267792 93838
rect 267740 93774 267792 93780
rect 267278 73808 267334 73817
rect 267278 73743 267334 73752
rect 267094 68232 267150 68241
rect 267094 68167 267150 68176
rect 269132 47666 269160 95066
rect 273350 94480 273406 94489
rect 273350 94415 273406 94424
rect 270592 93220 270644 93226
rect 270592 93162 270644 93168
rect 269120 47660 269172 47666
rect 269120 47602 269172 47608
rect 268384 47592 268436 47598
rect 268384 47534 268436 47540
rect 267004 46300 267056 46306
rect 267004 46242 267056 46248
rect 266372 16546 266584 16574
rect 264336 13796 264388 13802
rect 264336 13738 264388 13744
rect 264244 11756 264296 11762
rect 264244 11698 264296 11704
rect 264348 6914 264376 13738
rect 264164 6886 264376 6914
rect 262784 598 262996 626
rect 262784 490 262812 598
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 462 262812 490
rect 262968 480 262996 598
rect 264164 480 264192 6886
rect 265348 4140 265400 4146
rect 265348 4082 265400 4088
rect 265360 480 265388 4082
rect 266556 480 266584 16546
rect 267740 11960 267792 11966
rect 267740 11902 267792 11908
rect 267752 480 267780 11902
rect 268396 6905 268424 47534
rect 269764 46232 269816 46238
rect 269764 46174 269816 46180
rect 269118 29608 269174 29617
rect 269118 29543 269174 29552
rect 268476 25628 268528 25634
rect 268476 25570 268528 25576
rect 268488 12374 268516 25570
rect 269132 16574 269160 29543
rect 269132 16546 269712 16574
rect 268476 12368 268528 12374
rect 268476 12310 268528 12316
rect 268488 11966 268516 12310
rect 268476 11960 268528 11966
rect 268476 11902 268528 11908
rect 268382 6896 268438 6905
rect 268382 6831 268438 6840
rect 268396 4078 268424 6831
rect 268384 4072 268436 4078
rect 268384 4014 268436 4020
rect 268844 4072 268896 4078
rect 268844 4014 268896 4020
rect 268856 480 268884 4014
rect 269684 3482 269712 16546
rect 269776 4146 269804 46174
rect 270500 28280 270552 28286
rect 270500 28222 270552 28228
rect 270512 26246 270540 28222
rect 270500 26240 270552 26246
rect 270500 26182 270552 26188
rect 269764 4140 269816 4146
rect 269764 4082 269816 4088
rect 269684 3454 270080 3482
rect 270052 480 270080 3454
rect 270512 626 270540 26182
rect 270604 2174 270632 93162
rect 273166 66872 273222 66881
rect 273166 66807 273222 66816
rect 273180 6914 273208 66807
rect 273364 35193 273392 94415
rect 274008 93838 274036 96084
rect 273996 93832 274048 93838
rect 273996 93774 274048 93780
rect 276018 91896 276074 91905
rect 276018 91831 276074 91840
rect 276032 88330 276060 91831
rect 276020 88324 276072 88330
rect 276020 88266 276072 88272
rect 273902 38040 273958 38049
rect 273902 37975 273958 37984
rect 273350 35184 273406 35193
rect 273350 35119 273406 35128
rect 273916 12345 273944 37975
rect 274640 32428 274692 32434
rect 274640 32370 274692 32376
rect 274652 27606 274680 32370
rect 274640 27600 274692 27606
rect 274640 27542 274692 27548
rect 274652 16574 274680 27542
rect 274652 16546 274864 16574
rect 273902 12336 273958 12345
rect 273902 12271 273958 12280
rect 274546 12336 274602 12345
rect 274546 12271 274602 12280
rect 273180 6886 273300 6914
rect 273272 3534 273300 6886
rect 274560 3534 274588 12271
rect 272432 3528 272484 3534
rect 272432 3470 272484 3476
rect 273260 3528 273312 3534
rect 273260 3470 273312 3476
rect 273628 3528 273680 3534
rect 273628 3470 273680 3476
rect 274548 3528 274600 3534
rect 274548 3470 274600 3476
rect 271788 2780 271840 2786
rect 271788 2722 271840 2728
rect 271800 2174 271828 2722
rect 270592 2168 270644 2174
rect 270592 2110 270644 2116
rect 271788 2168 271840 2174
rect 271788 2110 271840 2116
rect 270512 598 270816 626
rect 270788 490 270816 598
rect 271064 598 271276 626
rect 271064 490 271092 598
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 462 271092 490
rect 271248 480 271276 598
rect 272444 480 272472 3470
rect 273640 480 273668 3470
rect 274836 480 274864 16546
rect 276032 480 276060 88266
rect 279068 84153 279096 103486
rect 279422 99648 279478 99657
rect 279422 99583 279478 99592
rect 279330 96656 279386 96665
rect 279330 96591 279386 96600
rect 279344 95033 279372 96591
rect 279436 95198 279464 99583
rect 280158 98560 280214 98569
rect 280158 98495 280214 98504
rect 280066 95840 280122 95849
rect 280066 95775 280122 95784
rect 279424 95192 279476 95198
rect 279424 95134 279476 95140
rect 279330 95024 279386 95033
rect 279330 94959 279386 94968
rect 280080 93809 280108 95775
rect 280172 95169 280200 98495
rect 280158 95160 280214 95169
rect 280158 95095 280214 95104
rect 280066 93800 280122 93809
rect 280066 93735 280122 93744
rect 280356 91050 280384 145007
rect 280816 143585 280844 177278
rect 281538 175536 281594 175545
rect 281538 175471 281594 175480
rect 281552 175302 281580 175471
rect 281540 175296 281592 175302
rect 281540 175238 281592 175244
rect 281540 169720 281592 169726
rect 281540 169662 281592 169668
rect 281552 168745 281580 169662
rect 281538 168736 281594 168745
rect 281538 168671 281594 168680
rect 281644 165617 281672 189722
rect 281630 165608 281686 165617
rect 281630 165543 281686 165552
rect 281632 162852 281684 162858
rect 281632 162794 281684 162800
rect 281644 162625 281672 162794
rect 281630 162616 281686 162625
rect 281630 162551 281686 162560
rect 281540 157412 281592 157418
rect 281540 157354 281592 157360
rect 281552 155689 281580 157354
rect 281736 157321 281764 282950
rect 282196 246265 282224 307838
rect 283576 280634 283604 310383
rect 283564 280628 283616 280634
rect 283564 280570 283616 280576
rect 283564 246356 283616 246362
rect 283564 246298 283616 246304
rect 282182 246256 282238 246265
rect 282182 246191 282238 246200
rect 283196 238876 283248 238882
rect 283196 238818 283248 238824
rect 282182 237960 282238 237969
rect 282182 237895 282238 237904
rect 282196 187202 282224 237895
rect 282276 209160 282328 209166
rect 282276 209102 282328 209108
rect 282184 187196 282236 187202
rect 282184 187138 282236 187144
rect 282288 177954 282316 209102
rect 283104 181552 283156 181558
rect 283104 181494 283156 181500
rect 283012 178764 283064 178770
rect 283012 178706 283064 178712
rect 282276 177948 282328 177954
rect 282276 177890 282328 177896
rect 281908 175976 281960 175982
rect 281908 175918 281960 175924
rect 281816 175228 281868 175234
rect 281816 175170 281868 175176
rect 281828 174049 281856 175170
rect 281814 174040 281870 174049
rect 281814 173975 281870 173984
rect 281920 169425 281948 175918
rect 281906 169416 281962 169425
rect 281906 169351 281962 169360
rect 281908 167000 281960 167006
rect 281908 166942 281960 166948
rect 281920 166433 281948 166942
rect 281906 166424 281962 166433
rect 281906 166359 281962 166368
rect 282184 164960 282236 164966
rect 282184 164902 282236 164908
rect 282826 164928 282882 164937
rect 281816 163532 281868 163538
rect 281816 163474 281868 163480
rect 281828 158817 281856 163474
rect 281908 161832 281960 161838
rect 281906 161800 281908 161809
rect 281960 161800 281962 161809
rect 281906 161735 281962 161744
rect 281814 158808 281870 158817
rect 281814 158743 281870 158752
rect 282092 158704 282144 158710
rect 282092 158646 282144 158652
rect 282104 158001 282132 158646
rect 282090 157992 282146 158001
rect 282090 157927 282146 157936
rect 281722 157312 281778 157321
rect 281722 157247 281778 157256
rect 281538 155680 281594 155689
rect 281538 155615 281594 155624
rect 282092 154488 282144 154494
rect 282092 154430 282144 154436
rect 282104 154193 282132 154430
rect 282090 154184 282146 154193
rect 282090 154119 282146 154128
rect 282196 152697 282224 164902
rect 282826 164863 282882 164872
rect 282840 164286 282868 164863
rect 282828 164280 282880 164286
rect 282828 164222 282880 164228
rect 282826 164112 282882 164121
rect 282826 164047 282882 164056
rect 282840 163130 282868 164047
rect 282828 163124 282880 163130
rect 282828 163066 282880 163072
rect 282828 161424 282880 161430
rect 282828 161366 282880 161372
rect 282840 161129 282868 161366
rect 282826 161120 282882 161129
rect 282826 161055 282882 161064
rect 282828 160472 282880 160478
rect 282828 160414 282880 160420
rect 282840 160313 282868 160414
rect 282826 160304 282882 160313
rect 282826 160239 282882 160248
rect 282828 160064 282880 160070
rect 282828 160006 282880 160012
rect 282840 159497 282868 160006
rect 282826 159488 282882 159497
rect 282826 159423 282882 159432
rect 282276 155916 282328 155922
rect 282276 155858 282328 155864
rect 282288 155009 282316 155858
rect 282274 155000 282330 155009
rect 282274 154935 282330 154944
rect 282828 154556 282880 154562
rect 282828 154498 282880 154504
rect 282840 153513 282868 154498
rect 282826 153504 282882 153513
rect 282826 153439 282882 153448
rect 282182 152688 282238 152697
rect 282182 152623 282238 152632
rect 281908 151768 281960 151774
rect 281908 151710 281960 151716
rect 281920 151201 281948 151710
rect 281906 151192 281962 151201
rect 281906 151127 281962 151136
rect 282276 151088 282328 151094
rect 282276 151030 282328 151036
rect 282184 148980 282236 148986
rect 282184 148922 282236 148928
rect 282196 148073 282224 148922
rect 282182 148064 282238 148073
rect 282182 147999 282238 148008
rect 281724 147620 281776 147626
rect 281724 147562 281776 147568
rect 281736 147393 281764 147562
rect 281722 147384 281778 147393
rect 281722 147319 281778 147328
rect 280896 144220 280948 144226
rect 280896 144162 280948 144168
rect 280802 143576 280858 143585
rect 280802 143511 280858 143520
rect 280908 128353 280936 144162
rect 282288 142154 282316 151030
rect 282736 150408 282788 150414
rect 282736 150350 282788 150356
rect 282826 150376 282882 150385
rect 282748 149705 282776 150350
rect 282826 150311 282828 150320
rect 282880 150311 282882 150320
rect 282828 150282 282880 150288
rect 282734 149696 282790 149705
rect 282734 149631 282790 149640
rect 282828 149048 282880 149054
rect 282828 148990 282880 148996
rect 282840 148889 282868 148990
rect 282826 148880 282882 148889
rect 282826 148815 282882 148824
rect 282828 147552 282880 147558
rect 282828 147494 282880 147500
rect 282840 146577 282868 147494
rect 282826 146568 282882 146577
rect 282826 146503 282882 146512
rect 282828 146260 282880 146266
rect 282828 146202 282880 146208
rect 282840 145897 282868 146202
rect 282826 145888 282882 145897
rect 282826 145823 282882 145832
rect 282828 144900 282880 144906
rect 282828 144842 282880 144848
rect 282840 144265 282868 144842
rect 282826 144256 282882 144265
rect 282826 144191 282882 144200
rect 283024 142154 283052 178706
rect 283116 142769 283144 181494
rect 283208 157418 283236 238818
rect 283576 178770 283604 246298
rect 284312 193089 284340 377590
rect 285586 359544 285642 359553
rect 285586 359479 285642 359488
rect 285600 349897 285628 359479
rect 285586 349888 285642 349897
rect 285586 349823 285642 349832
rect 284942 321600 284998 321609
rect 284942 321535 284998 321544
rect 284956 249150 284984 321535
rect 285692 309913 285720 377590
rect 287992 374649 288020 377604
rect 289648 375329 289676 377604
rect 291212 377590 291318 377618
rect 292592 377590 292974 377618
rect 293972 377590 294630 377618
rect 295352 377590 296286 377618
rect 289634 375320 289690 375329
rect 289634 375255 289690 375264
rect 287978 374640 288034 374649
rect 287978 374575 288034 374584
rect 290464 374060 290516 374066
rect 290464 374002 290516 374008
rect 286232 344344 286284 344350
rect 286230 344312 286232 344321
rect 286284 344312 286286 344321
rect 286230 344247 286286 344256
rect 287702 341592 287758 341601
rect 287702 341527 287758 341536
rect 287058 314936 287114 314945
rect 287058 314871 287114 314880
rect 285678 309904 285734 309913
rect 285678 309839 285734 309848
rect 286416 280832 286468 280838
rect 286416 280774 286468 280780
rect 286324 279472 286376 279478
rect 286324 279414 286376 279420
rect 285036 277432 285088 277438
rect 285036 277374 285088 277380
rect 284944 249144 284996 249150
rect 284944 249086 284996 249092
rect 284944 236088 284996 236094
rect 284944 236030 284996 236036
rect 284392 232552 284444 232558
rect 284392 232494 284444 232500
rect 284298 193080 284354 193089
rect 284298 193015 284354 193024
rect 283564 178764 283616 178770
rect 283564 178706 283616 178712
rect 284300 178016 284352 178022
rect 284298 177984 284300 177993
rect 284352 177984 284354 177993
rect 284298 177919 284354 177928
rect 283196 157412 283248 157418
rect 283196 157354 283248 157360
rect 283102 142760 283158 142769
rect 283102 142695 283158 142704
rect 282196 142126 282316 142154
rect 282932 142126 283052 142154
rect 281908 141772 281960 141778
rect 281908 141714 281960 141720
rect 281920 141273 281948 141714
rect 281906 141264 281962 141273
rect 281906 141199 281962 141208
rect 281632 137964 281684 137970
rect 281632 137906 281684 137912
rect 281644 137465 281672 137906
rect 281630 137456 281686 137465
rect 281630 137391 281686 137400
rect 281724 132388 281776 132394
rect 281724 132330 281776 132336
rect 281736 132161 281764 132330
rect 281722 132152 281778 132161
rect 281722 132087 281778 132096
rect 282092 129736 282144 129742
rect 282092 129678 282144 129684
rect 282104 129033 282132 129678
rect 282090 129024 282146 129033
rect 282090 128959 282146 128968
rect 280894 128344 280950 128353
rect 280894 128279 280950 128288
rect 282196 127537 282224 142126
rect 282828 142112 282880 142118
rect 282826 142080 282828 142089
rect 282880 142080 282882 142089
rect 282826 142015 282882 142024
rect 282736 140752 282788 140758
rect 282736 140694 282788 140700
rect 282748 139777 282776 140694
rect 282826 140448 282882 140457
rect 282826 140383 282882 140392
rect 282734 139768 282790 139777
rect 282734 139703 282790 139712
rect 282840 139602 282868 140383
rect 282828 139596 282880 139602
rect 282828 139538 282880 139544
rect 282828 139392 282880 139398
rect 282828 139334 282880 139340
rect 282840 138961 282868 139334
rect 282826 138952 282882 138961
rect 282826 138887 282882 138896
rect 282826 138272 282882 138281
rect 282932 138258 282960 142126
rect 282882 138230 282960 138258
rect 282826 138207 282882 138216
rect 282276 136060 282328 136066
rect 282276 136002 282328 136008
rect 282288 135969 282316 136002
rect 282274 135960 282330 135969
rect 282274 135895 282330 135904
rect 282828 133884 282880 133890
rect 282828 133826 282880 133832
rect 282840 132841 282868 133826
rect 282826 132832 282882 132841
rect 282826 132767 282882 132776
rect 282644 132456 282696 132462
rect 282644 132398 282696 132404
rect 282656 131345 282684 132398
rect 282642 131336 282698 131345
rect 282642 131271 282698 131280
rect 282276 131096 282328 131102
rect 282276 131038 282328 131044
rect 282288 130665 282316 131038
rect 282828 131028 282880 131034
rect 282828 130970 282880 130976
rect 282274 130656 282330 130665
rect 282274 130591 282330 130600
rect 282734 130384 282790 130393
rect 282734 130319 282790 130328
rect 282182 127528 282238 127537
rect 282182 127463 282238 127472
rect 282276 126948 282328 126954
rect 282276 126890 282328 126896
rect 281722 126848 281778 126857
rect 281722 126783 281778 126792
rect 280434 121408 280490 121417
rect 280434 121343 280490 121352
rect 280448 92478 280476 121343
rect 281540 111444 281592 111450
rect 281540 111386 281592 111392
rect 281552 110809 281580 111386
rect 281538 110800 281594 110809
rect 281538 110735 281594 110744
rect 281540 104848 281592 104854
rect 281540 104790 281592 104796
rect 281552 104009 281580 104790
rect 281538 104000 281594 104009
rect 281538 103935 281594 103944
rect 281630 103184 281686 103193
rect 281630 103119 281686 103128
rect 280526 100872 280582 100881
rect 280526 100807 280582 100816
rect 280436 92472 280488 92478
rect 280436 92414 280488 92420
rect 280344 91044 280396 91050
rect 280344 90986 280396 90992
rect 280540 88262 280568 100807
rect 280528 88256 280580 88262
rect 280528 88198 280580 88204
rect 281644 86902 281672 103119
rect 281736 90982 281764 126783
rect 282000 126268 282052 126274
rect 282000 126210 282052 126216
rect 282012 123729 282040 126210
rect 282288 126041 282316 126890
rect 282274 126032 282330 126041
rect 282274 125967 282330 125976
rect 282368 125588 282420 125594
rect 282368 125530 282420 125536
rect 282274 124808 282330 124817
rect 282274 124743 282330 124752
rect 281998 123720 282054 123729
rect 281998 123655 282054 123664
rect 282184 117972 282236 117978
rect 282184 117914 282236 117920
rect 282196 115433 282224 117914
rect 282288 116929 282316 124743
rect 282380 124545 282408 125530
rect 282748 125225 282776 130319
rect 282840 129849 282868 130970
rect 282826 129840 282882 129849
rect 282826 129775 282882 129784
rect 282828 127628 282880 127634
rect 282828 127570 282880 127576
rect 282734 125216 282790 125225
rect 282734 125151 282790 125160
rect 282366 124536 282422 124545
rect 282366 124471 282422 124480
rect 282736 123480 282788 123486
rect 282736 123422 282788 123428
rect 282748 119241 282776 123422
rect 282840 123049 282868 127570
rect 282826 123040 282882 123049
rect 282826 122975 282882 122984
rect 282828 122800 282880 122806
rect 282828 122742 282880 122748
rect 282840 122233 282868 122742
rect 282826 122224 282882 122233
rect 282826 122159 282882 122168
rect 282828 121440 282880 121446
rect 282828 121382 282880 121388
rect 282840 120737 282868 121382
rect 282826 120728 282882 120737
rect 282826 120663 282882 120672
rect 282828 120080 282880 120086
rect 282828 120022 282880 120028
rect 282840 119921 282868 120022
rect 282826 119912 282882 119921
rect 282826 119847 282882 119856
rect 282734 119232 282790 119241
rect 282734 119167 282790 119176
rect 282552 118448 282604 118454
rect 282552 118390 282604 118396
rect 282564 117609 282592 118390
rect 282550 117600 282606 117609
rect 282550 117535 282606 117544
rect 282274 116920 282330 116929
rect 282274 116855 282330 116864
rect 282276 116612 282328 116618
rect 282276 116554 282328 116560
rect 282182 115424 282238 115433
rect 282182 115359 282238 115368
rect 281814 113112 281870 113121
rect 281814 113047 281816 113056
rect 281868 113047 281870 113056
rect 281816 113018 281868 113024
rect 282288 108497 282316 116554
rect 282828 116136 282880 116142
rect 282826 116104 282828 116113
rect 282880 116104 282882 116113
rect 282826 116039 282882 116048
rect 282460 115932 282512 115938
rect 282460 115874 282512 115880
rect 282472 114617 282500 115874
rect 282458 114608 282514 114617
rect 282458 114543 282514 114552
rect 282828 114504 282880 114510
rect 282828 114446 282880 114452
rect 282840 113801 282868 114446
rect 282826 113792 282882 113801
rect 282826 113727 282882 113736
rect 282828 113144 282880 113150
rect 282828 113086 282880 113092
rect 282840 112305 282868 113086
rect 282826 112296 282882 112305
rect 282826 112231 282882 112240
rect 282826 111616 282882 111625
rect 282826 111551 282828 111560
rect 282880 111551 282882 111560
rect 282828 111522 282880 111528
rect 282828 110424 282880 110430
rect 282828 110366 282880 110372
rect 282840 109313 282868 110366
rect 282826 109304 282882 109313
rect 282826 109239 282882 109248
rect 282368 108996 282420 109002
rect 282368 108938 282420 108944
rect 282274 108488 282330 108497
rect 282274 108423 282330 108432
rect 282380 107817 282408 108938
rect 282366 107808 282422 107817
rect 282366 107743 282422 107752
rect 282828 107636 282880 107642
rect 282828 107578 282880 107584
rect 282840 107001 282868 107578
rect 282826 106992 282882 107001
rect 282826 106927 282882 106936
rect 284404 104854 284432 232494
rect 284956 224913 284984 236030
rect 285048 232558 285076 277374
rect 285128 249892 285180 249898
rect 285128 249834 285180 249840
rect 285140 238066 285168 249834
rect 285128 238060 285180 238066
rect 285128 238002 285180 238008
rect 285036 232552 285088 232558
rect 285036 232494 285088 232500
rect 285770 228304 285826 228313
rect 285770 228239 285826 228248
rect 284942 224904 284998 224913
rect 284942 224839 284998 224848
rect 284956 219434 284984 224839
rect 284496 219406 284984 219434
rect 284496 113082 284524 219406
rect 285680 217388 285732 217394
rect 285680 217330 285732 217336
rect 284944 203584 284996 203590
rect 284944 203526 284996 203532
rect 284576 187196 284628 187202
rect 284576 187138 284628 187144
rect 284484 113076 284536 113082
rect 284484 113018 284536 113024
rect 284588 111450 284616 187138
rect 284666 177440 284722 177449
rect 284956 177410 284984 203526
rect 284666 177375 284722 177384
rect 284944 177404 284996 177410
rect 284680 169726 284708 177375
rect 284944 177346 284996 177352
rect 284668 169720 284720 169726
rect 284668 169662 284720 169668
rect 285692 136066 285720 217330
rect 285680 136060 285732 136066
rect 285680 136002 285732 136008
rect 285680 127696 285732 127702
rect 285680 127638 285732 127644
rect 284576 111444 284628 111450
rect 284576 111386 284628 111392
rect 284392 104848 284444 104854
rect 284392 104790 284444 104796
rect 282000 100020 282052 100026
rect 282000 99962 282052 99968
rect 282012 97889 282040 99962
rect 281998 97880 282054 97889
rect 281998 97815 282054 97824
rect 281724 90976 281776 90982
rect 281724 90918 281776 90924
rect 281632 86896 281684 86902
rect 281632 86838 281684 86844
rect 279054 84144 279110 84153
rect 279054 84079 279110 84088
rect 278042 82104 278098 82113
rect 278042 82039 278098 82048
rect 277400 28280 277452 28286
rect 277400 28222 277452 28228
rect 277412 16574 277440 28222
rect 277412 16546 277992 16574
rect 276110 3496 276166 3505
rect 277964 3482 277992 16546
rect 278056 6186 278084 82039
rect 280802 77888 280858 77897
rect 280802 77823 280858 77832
rect 279424 33788 279476 33794
rect 279424 33730 279476 33736
rect 278044 6180 278096 6186
rect 278044 6122 278096 6128
rect 279436 4146 279464 33730
rect 280712 12504 280764 12510
rect 280712 12446 280764 12452
rect 279424 4140 279476 4146
rect 279424 4082 279476 4088
rect 279436 4026 279464 4082
rect 279436 3998 279556 4026
rect 276110 3431 276112 3440
rect 276164 3431 276166 3440
rect 277124 3460 277176 3466
rect 276112 3402 276164 3408
rect 277964 3454 278360 3482
rect 277124 3402 277176 3408
rect 277136 480 277164 3402
rect 278332 480 278360 3454
rect 279528 480 279556 3998
rect 280724 480 280752 12446
rect 280816 3913 280844 77823
rect 283562 64288 283618 64297
rect 283562 64223 283618 64232
rect 282182 55856 282238 55865
rect 282182 55791 282238 55800
rect 280894 26888 280950 26897
rect 280894 26823 280950 26832
rect 280908 13802 280936 26823
rect 280896 13796 280948 13802
rect 280896 13738 280948 13744
rect 280908 12510 280936 13738
rect 280896 12504 280948 12510
rect 280896 12446 280948 12452
rect 280802 3904 280858 3913
rect 280802 3839 280858 3848
rect 282196 3466 282224 55791
rect 283576 42770 283604 64223
rect 284944 64184 284996 64190
rect 284944 64126 284996 64132
rect 283564 42764 283616 42770
rect 283564 42706 283616 42712
rect 282276 29640 282328 29646
rect 282276 29582 282328 29588
rect 282288 4049 282316 29582
rect 283576 5574 283604 42706
rect 284956 24857 284984 64126
rect 284942 24848 284998 24857
rect 284942 24783 284998 24792
rect 284956 23497 284984 24783
rect 284298 23488 284354 23497
rect 284298 23423 284354 23432
rect 284942 23488 284998 23497
rect 284942 23423 284998 23432
rect 282828 5568 282880 5574
rect 282828 5510 282880 5516
rect 283564 5568 283616 5574
rect 283564 5510 283616 5516
rect 282274 4040 282330 4049
rect 282274 3975 282330 3984
rect 282184 3460 282236 3466
rect 282184 3402 282236 3408
rect 282288 1034 282316 3975
rect 282840 3482 282868 5510
rect 282840 3454 283144 3482
rect 281920 1006 282316 1034
rect 281920 480 281948 1006
rect 283116 480 283144 3454
rect 284312 480 284340 23423
rect 285692 16574 285720 127638
rect 285784 118454 285812 228239
rect 285864 180192 285916 180198
rect 285864 180134 285916 180140
rect 285876 141778 285904 180134
rect 286336 161838 286364 279414
rect 286428 236094 286456 280774
rect 286416 236088 286468 236094
rect 286416 236030 286468 236036
rect 286324 161832 286376 161838
rect 286324 161774 286376 161780
rect 285864 141772 285916 141778
rect 285864 141714 285916 141720
rect 285772 118448 285824 118454
rect 285772 118390 285824 118396
rect 287072 111586 287100 314871
rect 287716 311166 287744 341527
rect 287704 311160 287756 311166
rect 287704 311102 287756 311108
rect 288440 302252 288492 302258
rect 288440 302194 288492 302200
rect 288348 240848 288400 240854
rect 288348 240790 288400 240796
rect 288360 240174 288388 240790
rect 287244 240168 287296 240174
rect 287244 240110 287296 240116
rect 288348 240168 288400 240174
rect 288348 240110 288400 240116
rect 287256 219434 287284 240110
rect 287164 219406 287284 219434
rect 287164 116142 287192 219406
rect 287244 199504 287296 199510
rect 287244 199446 287296 199452
rect 287256 164286 287284 199446
rect 287334 177576 287390 177585
rect 287334 177511 287390 177520
rect 287244 164280 287296 164286
rect 287244 164222 287296 164228
rect 287348 160478 287376 177511
rect 287336 160472 287388 160478
rect 287336 160414 287388 160420
rect 288452 139602 288480 302194
rect 288532 258732 288584 258738
rect 288532 258674 288584 258680
rect 288544 258126 288572 258674
rect 288532 258120 288584 258126
rect 288532 258062 288584 258068
rect 288544 148986 288572 258062
rect 289910 251968 289966 251977
rect 289910 251903 289966 251912
rect 288624 198076 288676 198082
rect 288624 198018 288676 198024
rect 288532 148980 288584 148986
rect 288532 148922 288584 148928
rect 288440 139596 288492 139602
rect 288440 139538 288492 139544
rect 288636 129742 288664 198018
rect 288716 177948 288768 177954
rect 288716 177890 288768 177896
rect 288728 163130 288756 177890
rect 289820 177404 289872 177410
rect 289820 177346 289872 177352
rect 289832 171834 289860 177346
rect 289820 171828 289872 171834
rect 289820 171770 289872 171776
rect 288716 163124 288768 163130
rect 288716 163066 288768 163072
rect 289924 151094 289952 251903
rect 290096 227044 290148 227050
rect 290096 226986 290148 226992
rect 290004 210520 290056 210526
rect 290004 210462 290056 210468
rect 289912 151088 289964 151094
rect 289912 151030 289964 151036
rect 288624 129736 288676 129742
rect 288624 129678 288676 129684
rect 290016 121446 290044 210462
rect 290004 121440 290056 121446
rect 290004 121382 290056 121388
rect 287152 116136 287204 116142
rect 287152 116078 287204 116084
rect 290108 114510 290136 226986
rect 290476 225690 290504 374002
rect 291212 264314 291240 377590
rect 292592 327826 292620 377590
rect 292580 327820 292632 327826
rect 292580 327762 292632 327768
rect 293224 312588 293276 312594
rect 293224 312530 293276 312536
rect 293236 269006 293264 312530
rect 293972 301578 294000 377590
rect 294604 304972 294656 304978
rect 294604 304914 294656 304920
rect 293960 301572 294012 301578
rect 293960 301514 294012 301520
rect 294616 279478 294644 304914
rect 294604 279472 294656 279478
rect 294604 279414 294656 279420
rect 293960 276684 294012 276690
rect 293960 276626 294012 276632
rect 291844 269000 291896 269006
rect 291844 268942 291896 268948
rect 293224 269000 293276 269006
rect 293224 268942 293276 268948
rect 291200 264308 291252 264314
rect 291200 264250 291252 264256
rect 291106 251968 291162 251977
rect 291106 251903 291108 251912
rect 291160 251903 291162 251912
rect 291108 251874 291160 251880
rect 291200 246424 291252 246430
rect 291200 246366 291252 246372
rect 290464 225684 290516 225690
rect 290464 225626 290516 225632
rect 290096 114504 290148 114510
rect 290096 114446 290148 114452
rect 287060 111580 287112 111586
rect 287060 111522 287112 111528
rect 291212 107642 291240 246366
rect 291856 231810 291884 268942
rect 292580 265668 292632 265674
rect 292580 265610 292632 265616
rect 291292 231804 291344 231810
rect 291292 231746 291344 231752
rect 291844 231804 291896 231810
rect 291844 231746 291896 231752
rect 291304 123486 291332 231746
rect 291384 180124 291436 180130
rect 291384 180066 291436 180072
rect 291396 147558 291424 180066
rect 291474 178664 291530 178673
rect 291474 178599 291530 178608
rect 291488 167006 291516 178599
rect 291476 167000 291528 167006
rect 291476 166942 291528 166948
rect 291384 147552 291436 147558
rect 291384 147494 291436 147500
rect 291292 123480 291344 123486
rect 291292 123422 291344 123428
rect 292592 120086 292620 265610
rect 292764 258800 292816 258806
rect 292764 258742 292816 258748
rect 292670 196752 292726 196761
rect 292670 196687 292726 196696
rect 292580 120080 292632 120086
rect 292580 120022 292632 120028
rect 291200 107636 291252 107642
rect 291200 107578 291252 107584
rect 292578 100872 292634 100881
rect 292578 100807 292634 100816
rect 291198 97880 291254 97889
rect 291198 97815 291254 97824
rect 289818 93120 289874 93129
rect 289818 93055 289874 93064
rect 286322 91760 286378 91769
rect 286322 91695 286378 91704
rect 285692 16546 286272 16574
rect 285404 6180 285456 6186
rect 285404 6122 285456 6128
rect 285416 480 285444 6122
rect 286244 3482 286272 16546
rect 286336 4146 286364 91695
rect 288348 13116 288400 13122
rect 288348 13058 288400 13064
rect 288360 12209 288388 13058
rect 288346 12200 288402 12209
rect 288346 12135 288402 12144
rect 286324 4140 286376 4146
rect 286324 4082 286376 4088
rect 288360 3505 288388 12135
rect 288990 8256 289046 8265
rect 288990 8191 289046 8200
rect 289004 7614 289032 8191
rect 288992 7608 289044 7614
rect 288992 7550 289044 7556
rect 287794 3496 287850 3505
rect 286244 3454 286640 3482
rect 286612 480 286640 3454
rect 287794 3431 287850 3440
rect 288346 3496 288402 3505
rect 288346 3431 288402 3440
rect 287808 480 287836 3431
rect 289004 480 289032 7550
rect 289832 490 289860 93055
rect 291212 16574 291240 97815
rect 292486 66192 292542 66201
rect 292486 66127 292542 66136
rect 292500 65550 292528 66127
rect 292488 65544 292540 65550
rect 292488 65486 292540 65492
rect 291212 16546 291424 16574
rect 290016 598 290228 626
rect 290016 490 290044 598
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289832 462 290044 490
rect 290200 480 290228 598
rect 291396 480 291424 16546
rect 292500 3534 292528 65486
rect 292592 16574 292620 100807
rect 292684 63510 292712 196687
rect 292776 158710 292804 258742
rect 293222 184240 293278 184249
rect 293222 184175 293278 184184
rect 292764 158704 292816 158710
rect 292764 158646 292816 158652
rect 293236 101425 293264 184175
rect 293972 160070 294000 276626
rect 294604 272536 294656 272542
rect 294604 272478 294656 272484
rect 294052 181484 294104 181490
rect 294052 181426 294104 181432
rect 293960 160064 294012 160070
rect 293960 160006 294012 160012
rect 294064 144906 294092 181426
rect 294052 144900 294104 144906
rect 294052 144842 294104 144848
rect 293222 101416 293278 101425
rect 293222 101351 293278 101360
rect 293236 100881 293264 101351
rect 293222 100872 293278 100881
rect 293222 100807 293278 100816
rect 294616 82822 294644 272478
rect 294696 235272 294748 235278
rect 294696 235214 294748 235220
rect 294708 106282 294736 235214
rect 295352 229809 295380 377590
rect 297928 374066 297956 377604
rect 298744 374672 298796 374678
rect 298744 374614 298796 374620
rect 297916 374060 297968 374066
rect 297916 374002 297968 374008
rect 297364 365016 297416 365022
rect 297364 364958 297416 364964
rect 295432 292596 295484 292602
rect 295432 292538 295484 292544
rect 295338 229800 295394 229809
rect 295338 229735 295340 229744
rect 295392 229735 295394 229744
rect 295340 229706 295392 229712
rect 295338 185600 295394 185609
rect 295338 185535 295394 185544
rect 295352 163538 295380 185535
rect 295340 163532 295392 163538
rect 295340 163474 295392 163480
rect 295338 149152 295394 149161
rect 295338 149087 295394 149096
rect 294696 106276 294748 106282
rect 294696 106218 294748 106224
rect 294604 82816 294656 82822
rect 294604 82758 294656 82764
rect 292672 63504 292724 63510
rect 292672 63446 292724 63452
rect 292684 62830 292712 63446
rect 292672 62824 292724 62830
rect 292672 62766 292724 62772
rect 294616 28286 294644 82758
rect 294604 28280 294656 28286
rect 294604 28222 294656 28228
rect 295352 16574 295380 149087
rect 295444 110430 295472 292538
rect 295892 290488 295944 290494
rect 295892 290430 295944 290436
rect 295904 290057 295932 290430
rect 295522 290048 295578 290057
rect 295522 289983 295578 289992
rect 295890 290048 295946 290057
rect 295890 289983 295946 289992
rect 295536 142118 295564 289983
rect 297376 225622 297404 364958
rect 298100 298784 298152 298790
rect 298100 298726 298152 298732
rect 297454 289912 297510 289921
rect 297454 289847 297510 289856
rect 297468 283529 297496 289847
rect 297454 283520 297510 283529
rect 297454 283455 297510 283464
rect 298006 246392 298062 246401
rect 298006 246327 298062 246336
rect 298020 245721 298048 246327
rect 298006 245712 298062 245721
rect 298006 245647 298062 245656
rect 296812 225616 296864 225622
rect 296812 225558 296864 225564
rect 297364 225616 297416 225622
rect 297364 225558 297416 225564
rect 295982 224360 296038 224369
rect 295982 224295 296038 224304
rect 295996 144974 296024 224295
rect 296718 223000 296774 223009
rect 296718 222935 296774 222944
rect 295984 144968 296036 144974
rect 295984 144910 296036 144916
rect 295524 142112 295576 142118
rect 295524 142054 295576 142060
rect 295996 127702 296024 144910
rect 295984 127696 296036 127702
rect 295984 127638 296036 127644
rect 296732 117978 296760 222935
rect 296824 144226 296852 225558
rect 297914 223000 297970 223009
rect 297914 222935 297970 222944
rect 297928 222902 297956 222935
rect 297916 222896 297968 222902
rect 297916 222838 297968 222844
rect 296904 188352 296956 188358
rect 296904 188294 296956 188300
rect 296812 144220 296864 144226
rect 296812 144162 296864 144168
rect 296916 139398 296944 188294
rect 296904 139392 296956 139398
rect 296904 139334 296956 139340
rect 296720 117972 296772 117978
rect 296720 117914 296772 117920
rect 295432 110424 295484 110430
rect 295432 110366 295484 110372
rect 298020 96529 298048 245647
rect 298112 125594 298140 298726
rect 298756 240854 298784 374614
rect 299478 325000 299534 325009
rect 299478 324935 299534 324944
rect 298834 251832 298890 251841
rect 298834 251767 298890 251776
rect 298744 240848 298796 240854
rect 298744 240790 298796 240796
rect 298466 225584 298522 225593
rect 298466 225519 298522 225528
rect 298480 225010 298508 225519
rect 298468 225004 298520 225010
rect 298468 224946 298520 224952
rect 298742 218784 298798 218793
rect 298742 218719 298798 218728
rect 298192 178764 298244 178770
rect 298192 178706 298244 178712
rect 298204 126954 298232 178706
rect 298756 177342 298784 218719
rect 298744 177336 298796 177342
rect 298744 177278 298796 177284
rect 298848 146946 298876 251767
rect 298836 146940 298888 146946
rect 298836 146882 298888 146888
rect 298192 126948 298244 126954
rect 298192 126890 298244 126896
rect 298100 125588 298152 125594
rect 298100 125530 298152 125536
rect 298100 106956 298152 106962
rect 298100 106898 298152 106904
rect 298006 96520 298062 96529
rect 298006 96455 298062 96464
rect 297364 49020 297416 49026
rect 297364 48962 297416 48968
rect 297376 17950 297404 48962
rect 296720 17944 296772 17950
rect 296720 17886 296772 17892
rect 297364 17944 297416 17950
rect 297364 17886 297416 17892
rect 292592 16546 293264 16574
rect 295352 16546 295656 16574
rect 292578 7576 292634 7585
rect 292578 7511 292634 7520
rect 292592 3777 292620 7511
rect 292578 3768 292634 3777
rect 292578 3703 292634 3712
rect 292488 3528 292540 3534
rect 292488 3470 292540 3476
rect 292592 480 292620 3703
rect 293236 490 293264 16546
rect 294880 3528 294932 3534
rect 294880 3470 294932 3476
rect 293512 598 293724 626
rect 293512 490 293540 598
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 462 293540 490
rect 293696 480 293724 598
rect 294892 480 294920 3470
rect 295628 490 295656 16546
rect 296732 3534 296760 17886
rect 296720 3528 296772 3534
rect 296720 3470 296772 3476
rect 297272 3528 297324 3534
rect 297272 3470 297324 3476
rect 295904 598 296116 626
rect 295904 490 295932 598
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 462 295932 490
rect 296088 480 296116 598
rect 297284 480 297312 3470
rect 298112 490 298140 106898
rect 299492 46238 299520 324935
rect 299584 213926 299612 377604
rect 300872 377590 301254 377618
rect 302252 377590 302910 377618
rect 303632 377590 304566 377618
rect 305012 377590 306222 377618
rect 307878 377590 308444 377618
rect 300124 261588 300176 261594
rect 300124 261530 300176 261536
rect 299572 213920 299624 213926
rect 299572 213862 299624 213868
rect 299572 178696 299624 178702
rect 299572 178638 299624 178644
rect 299584 147626 299612 178638
rect 300136 173194 300164 261530
rect 300872 255338 300900 377590
rect 300860 255332 300912 255338
rect 300860 255274 300912 255280
rect 300216 213920 300268 213926
rect 300216 213862 300268 213868
rect 300124 173188 300176 173194
rect 300124 173130 300176 173136
rect 300228 164898 300256 213862
rect 300308 196648 300360 196654
rect 300308 196590 300360 196596
rect 300320 188358 300348 196590
rect 300308 188352 300360 188358
rect 300308 188294 300360 188300
rect 300216 164892 300268 164898
rect 300216 164834 300268 164840
rect 300872 151774 300900 255274
rect 300952 253224 301004 253230
rect 300952 253166 301004 253172
rect 300860 151768 300912 151774
rect 300860 151710 300912 151716
rect 299572 147620 299624 147626
rect 299572 147562 299624 147568
rect 300860 143540 300912 143546
rect 300860 143482 300912 143488
rect 300872 142186 300900 143482
rect 300860 142180 300912 142186
rect 300860 142122 300912 142128
rect 299662 86320 299718 86329
rect 299662 86255 299664 86264
rect 299716 86255 299718 86264
rect 299664 86226 299716 86232
rect 300768 46912 300820 46918
rect 300768 46854 300820 46860
rect 300780 46238 300808 46854
rect 299480 46232 299532 46238
rect 299480 46174 299532 46180
rect 300768 46232 300820 46238
rect 300768 46174 300820 46180
rect 300872 16574 300900 142122
rect 300964 137970 300992 253166
rect 302252 251938 302280 377590
rect 302884 369912 302936 369918
rect 302884 369854 302936 369860
rect 302332 313948 302384 313954
rect 302332 313890 302384 313896
rect 302344 313342 302372 313890
rect 302332 313336 302384 313342
rect 302332 313278 302384 313284
rect 302240 251932 302292 251938
rect 302240 251874 302292 251880
rect 301502 212120 301558 212129
rect 301502 212055 301558 212064
rect 301042 188456 301098 188465
rect 301042 188391 301098 188400
rect 300952 137964 301004 137970
rect 300952 137906 301004 137912
rect 301056 125497 301084 188391
rect 301516 143546 301544 212055
rect 302240 195288 302292 195294
rect 302240 195230 302292 195236
rect 302252 154494 302280 195230
rect 302240 154488 302292 154494
rect 302240 154430 302292 154436
rect 302344 146266 302372 313278
rect 302424 184952 302476 184958
rect 302424 184894 302476 184900
rect 302436 150346 302464 184894
rect 302424 150340 302476 150346
rect 302424 150282 302476 150288
rect 302332 146260 302384 146266
rect 302332 146202 302384 146208
rect 301504 143540 301556 143546
rect 301504 143482 301556 143488
rect 301042 125488 301098 125497
rect 301042 125423 301098 125432
rect 301318 125488 301374 125497
rect 301318 125423 301374 125432
rect 301332 124817 301360 125423
rect 301318 124808 301374 124817
rect 301318 124743 301374 124752
rect 300872 16546 301544 16574
rect 300766 11792 300822 11801
rect 300766 11727 300822 11736
rect 300674 7576 300730 7585
rect 300674 7511 300730 7520
rect 300688 4049 300716 7511
rect 299662 4040 299718 4049
rect 299662 3975 299718 3984
rect 300674 4040 300730 4049
rect 300674 3975 300730 3984
rect 298296 598 298508 626
rect 298296 490 298324 598
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 462 298324 490
rect 298480 480 298508 598
rect 299676 480 299704 3975
rect 300780 480 300808 11727
rect 301516 490 301544 16546
rect 302896 4078 302924 369854
rect 303632 293865 303660 377590
rect 305012 342961 305040 377590
rect 308416 374066 308444 377590
rect 309152 377590 309534 377618
rect 310532 377590 311190 377618
rect 308404 374060 308456 374066
rect 308404 374002 308456 374008
rect 307022 366344 307078 366353
rect 307022 366279 307078 366288
rect 304998 342952 305054 342961
rect 304998 342887 305054 342896
rect 305012 342281 305040 342887
rect 304998 342272 305054 342281
rect 304998 342207 305054 342216
rect 305642 342272 305698 342281
rect 305642 342207 305698 342216
rect 303618 293856 303674 293865
rect 303618 293791 303674 293800
rect 303632 292641 303660 293791
rect 303618 292632 303674 292641
rect 303618 292567 303674 292576
rect 304262 292632 304318 292641
rect 304262 292567 304318 292576
rect 303620 287700 303672 287706
rect 303620 287642 303672 287648
rect 303632 287094 303660 287642
rect 303620 287088 303672 287094
rect 303620 287030 303672 287036
rect 303632 132394 303660 287030
rect 304276 279478 304304 292567
rect 304998 291272 305054 291281
rect 304998 291207 305054 291216
rect 304264 279472 304316 279478
rect 304264 279414 304316 279420
rect 303712 260160 303764 260166
rect 303712 260102 303764 260108
rect 303724 259486 303752 260102
rect 303712 259480 303764 259486
rect 303712 259422 303764 259428
rect 303620 132388 303672 132394
rect 303620 132330 303672 132336
rect 303724 113150 303752 259422
rect 303896 195356 303948 195362
rect 303896 195298 303948 195304
rect 303804 182844 303856 182850
rect 303804 182786 303856 182792
rect 303816 131034 303844 182786
rect 303908 162858 303936 195298
rect 303896 162852 303948 162858
rect 303896 162794 303948 162800
rect 303804 131028 303856 131034
rect 303804 130970 303856 130976
rect 305012 122806 305040 291207
rect 305184 271176 305236 271182
rect 305184 271118 305236 271124
rect 305092 239488 305144 239494
rect 305092 239430 305144 239436
rect 305104 238785 305132 239430
rect 305090 238776 305146 238785
rect 305090 238711 305146 238720
rect 305000 122800 305052 122806
rect 305000 122742 305052 122748
rect 303712 113144 303764 113150
rect 303712 113086 303764 113092
rect 305104 109002 305132 238711
rect 305196 190454 305224 271118
rect 305656 225622 305684 342207
rect 306380 271924 306432 271930
rect 306380 271866 306432 271872
rect 305644 225616 305696 225622
rect 305644 225558 305696 225564
rect 305196 190426 305316 190454
rect 305184 175976 305236 175982
rect 305184 175918 305236 175924
rect 305196 175302 305224 175918
rect 305184 175296 305236 175302
rect 305184 175238 305236 175244
rect 305288 175234 305316 190426
rect 305644 175296 305696 175302
rect 305644 175238 305696 175244
rect 305276 175228 305328 175234
rect 305276 175170 305328 175176
rect 305092 108996 305144 109002
rect 305092 108938 305144 108944
rect 305656 86970 305684 175238
rect 306392 126274 306420 271866
rect 306472 200796 306524 200802
rect 306472 200738 306524 200744
rect 306484 154562 306512 200738
rect 306472 154556 306524 154562
rect 306472 154498 306524 154504
rect 306380 126268 306432 126274
rect 306380 126210 306432 126216
rect 305644 86964 305696 86970
rect 305644 86906 305696 86912
rect 304264 80708 304316 80714
rect 304264 80650 304316 80656
rect 302976 50380 303028 50386
rect 302976 50322 303028 50328
rect 302988 30977 303016 50322
rect 304276 31074 304304 80650
rect 304264 31068 304316 31074
rect 304264 31010 304316 31016
rect 302974 30968 303030 30977
rect 302974 30903 303030 30912
rect 302988 16574 303016 30903
rect 303620 28280 303672 28286
rect 303620 28222 303672 28228
rect 303632 16574 303660 28222
rect 302988 16546 303200 16574
rect 303632 16546 303936 16574
rect 302884 4072 302936 4078
rect 302884 4014 302936 4020
rect 301792 598 302004 626
rect 301792 490 301820 598
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 462 301820 490
rect 301976 480 302004 598
rect 303172 480 303200 16546
rect 303908 490 303936 16546
rect 307036 5506 307064 366279
rect 308416 363633 308444 374002
rect 308402 363624 308458 363633
rect 308402 363559 308458 363568
rect 309152 361554 309180 377590
rect 309876 374060 309928 374066
rect 309876 374002 309928 374008
rect 309784 369164 309836 369170
rect 309784 369106 309836 369112
rect 309140 361548 309192 361554
rect 309140 361490 309192 361496
rect 309796 341465 309824 369106
rect 309782 341456 309838 341465
rect 309782 341391 309838 341400
rect 309796 340921 309824 341391
rect 309782 340912 309838 340921
rect 309782 340847 309838 340856
rect 308404 318844 308456 318850
rect 308404 318786 308456 318792
rect 308416 280809 308444 318786
rect 309138 305008 309194 305017
rect 309138 304943 309194 304952
rect 308402 280800 308458 280809
rect 308402 280735 308458 280744
rect 307116 274712 307168 274718
rect 307116 274654 307168 274660
rect 307128 159390 307156 274654
rect 307668 272536 307720 272542
rect 307668 272478 307720 272484
rect 307680 271930 307708 272478
rect 307668 271924 307720 271930
rect 307668 271866 307720 271872
rect 307760 250572 307812 250578
rect 307760 250514 307812 250520
rect 307772 250073 307800 250514
rect 307758 250064 307814 250073
rect 307758 249999 307814 250008
rect 307116 159384 307168 159390
rect 307116 159326 307168 159332
rect 307116 140072 307168 140078
rect 307116 140014 307168 140020
rect 306748 5500 306800 5506
rect 306748 5442 306800 5448
rect 307024 5500 307076 5506
rect 307024 5442 307076 5448
rect 305552 4140 305604 4146
rect 305552 4082 305604 4088
rect 304184 598 304396 626
rect 304184 490 304212 598
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 462 304212 490
rect 304368 480 304396 598
rect 305564 480 305592 4082
rect 306760 480 306788 5442
rect 307128 4146 307156 140014
rect 307772 116618 307800 249999
rect 307852 249144 307904 249150
rect 307852 249086 307904 249092
rect 307864 150414 307892 249086
rect 308404 207664 308456 207670
rect 308404 207606 308456 207612
rect 308416 167686 308444 207606
rect 308404 167680 308456 167686
rect 308404 167622 308456 167628
rect 307852 150408 307904 150414
rect 307852 150350 307904 150356
rect 307760 116612 307812 116618
rect 307760 116554 307812 116560
rect 309152 115938 309180 304943
rect 309784 279540 309836 279546
rect 309784 279482 309836 279488
rect 309232 256012 309284 256018
rect 309232 255954 309284 255960
rect 309140 115932 309192 115938
rect 309140 115874 309192 115880
rect 309244 100026 309272 255954
rect 309796 153882 309824 279482
rect 309888 251938 309916 374002
rect 310428 305652 310480 305658
rect 310428 305594 310480 305600
rect 310440 305017 310468 305594
rect 310426 305008 310482 305017
rect 310426 304943 310482 304952
rect 309876 251932 309928 251938
rect 309876 251874 309928 251880
rect 309874 199336 309930 199345
rect 309874 199271 309930 199280
rect 309784 153876 309836 153882
rect 309784 153818 309836 153824
rect 309782 119368 309838 119377
rect 309782 119303 309838 119312
rect 309232 100020 309284 100026
rect 309232 99962 309284 99968
rect 309138 84824 309194 84833
rect 309138 84759 309194 84768
rect 308402 54496 308458 54505
rect 308402 54431 308458 54440
rect 308416 6866 308444 54431
rect 308404 6860 308456 6866
rect 308404 6802 308456 6808
rect 307116 4140 307168 4146
rect 307116 4082 307168 4088
rect 308416 4049 308444 6802
rect 308402 4040 308458 4049
rect 308402 3975 308458 3984
rect 309046 4040 309102 4049
rect 309046 3975 309102 3984
rect 307944 3528 307996 3534
rect 307944 3470 307996 3476
rect 307956 480 307984 3470
rect 309060 480 309088 3975
rect 309152 3534 309180 84759
rect 309796 6866 309824 119303
rect 309888 113150 309916 199271
rect 309876 113144 309928 113150
rect 309876 113086 309928 113092
rect 310532 60625 310560 377590
rect 312832 375358 312860 377604
rect 313292 377590 314502 377618
rect 311900 375352 311952 375358
rect 311900 375294 311952 375300
rect 312820 375352 312872 375358
rect 312820 375294 312872 375300
rect 311912 369170 311940 375294
rect 311900 369164 311952 369170
rect 311900 369106 311952 369112
rect 311898 340912 311954 340921
rect 311898 340847 311954 340856
rect 310612 242208 310664 242214
rect 310612 242150 310664 242156
rect 310624 241534 310652 242150
rect 310612 241528 310664 241534
rect 310612 241470 310664 241476
rect 310624 149054 310652 241470
rect 310704 188352 310756 188358
rect 310704 188294 310756 188300
rect 310716 164966 310744 188294
rect 310704 164960 310756 164966
rect 310704 164902 310756 164908
rect 310612 149048 310664 149054
rect 310612 148990 310664 148996
rect 310518 60616 310574 60625
rect 310518 60551 310574 60560
rect 311162 60616 311218 60625
rect 311162 60551 311218 60560
rect 309876 32428 309928 32434
rect 309876 32370 309928 32376
rect 309784 6860 309836 6866
rect 309784 6802 309836 6808
rect 309888 4078 309916 32370
rect 311176 15162 311204 60551
rect 311912 59362 311940 340847
rect 313292 334626 313320 377590
rect 316144 374678 316172 377604
rect 317984 375358 318012 377604
rect 319640 376689 319668 377604
rect 320284 377590 321310 377618
rect 319626 376680 319682 376689
rect 319626 376615 319682 376624
rect 317972 375352 318024 375358
rect 317972 375294 318024 375300
rect 316132 374672 316184 374678
rect 316132 374614 316184 374620
rect 319640 373994 319668 376615
rect 320180 375352 320232 375358
rect 320180 375294 320232 375300
rect 319456 373966 319668 373994
rect 318064 369164 318116 369170
rect 318064 369106 318116 369112
rect 316684 366376 316736 366382
rect 316684 366318 316736 366324
rect 313280 334620 313332 334626
rect 313280 334562 313332 334568
rect 313924 309800 313976 309806
rect 313924 309742 313976 309748
rect 311992 268388 312044 268394
rect 311992 268330 312044 268336
rect 312004 267782 312032 268330
rect 311992 267776 312044 267782
rect 311992 267718 312044 267724
rect 312004 155922 312032 267718
rect 313280 244996 313332 245002
rect 313280 244938 313332 244944
rect 311992 155916 312044 155922
rect 311992 155858 312044 155864
rect 313292 130393 313320 244938
rect 313372 236700 313424 236706
rect 313372 236642 313424 236648
rect 313384 236026 313412 236642
rect 313372 236020 313424 236026
rect 313372 235962 313424 235968
rect 313384 133890 313412 235962
rect 313372 133884 313424 133890
rect 313372 133826 313424 133832
rect 313278 130384 313334 130393
rect 313278 130319 313334 130328
rect 311900 59356 311952 59362
rect 311900 59298 311952 59304
rect 311912 58682 311940 59298
rect 311900 58676 311952 58682
rect 311900 58618 311952 58624
rect 313936 34513 313964 309742
rect 314660 253292 314712 253298
rect 314660 253234 314712 253240
rect 314672 252618 314700 253234
rect 314660 252612 314712 252618
rect 314660 252554 314712 252560
rect 314672 127634 314700 252554
rect 316040 249824 316092 249830
rect 316040 249766 316092 249772
rect 315302 193896 315358 193905
rect 315302 193831 315358 193840
rect 314660 127628 314712 127634
rect 314660 127570 314712 127576
rect 314660 37936 314712 37942
rect 314660 37878 314712 37884
rect 313922 34504 313978 34513
rect 313922 34439 313978 34448
rect 314566 34504 314622 34513
rect 314566 34439 314622 34448
rect 311164 15156 311216 15162
rect 311164 15098 311216 15104
rect 311440 10396 311492 10402
rect 311440 10338 311492 10344
rect 309876 4072 309928 4078
rect 309876 4014 309928 4020
rect 309140 3528 309192 3534
rect 309140 3470 309192 3476
rect 309888 490 309916 4014
rect 310072 598 310284 626
rect 310072 490 310100 598
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309888 462 310100 490
rect 310256 480 310284 598
rect 311452 480 311480 10338
rect 314580 3534 314608 34439
rect 313832 3528 313884 3534
rect 313832 3470 313884 3476
rect 314568 3528 314620 3534
rect 314568 3470 314620 3476
rect 312636 3460 312688 3466
rect 312636 3402 312688 3408
rect 312648 480 312676 3402
rect 313844 480 313872 3470
rect 314672 490 314700 37878
rect 315316 4146 315344 193831
rect 316052 131102 316080 249766
rect 316696 230353 316724 366318
rect 317328 363656 317380 363662
rect 317328 363598 317380 363604
rect 317340 260846 317368 363598
rect 317604 322244 317656 322250
rect 317604 322186 317656 322192
rect 317328 260840 317380 260846
rect 317328 260782 317380 260788
rect 317328 250504 317380 250510
rect 317328 250446 317380 250452
rect 317340 249830 317368 250446
rect 317328 249824 317380 249830
rect 317328 249766 317380 249772
rect 317512 239420 317564 239426
rect 317512 239362 317564 239368
rect 317524 238814 317552 239362
rect 317512 238808 317564 238814
rect 317512 238750 317564 238756
rect 316130 230344 316186 230353
rect 316130 230279 316186 230288
rect 316682 230344 316738 230353
rect 316682 230279 316738 230288
rect 316144 175982 316172 230279
rect 316774 200832 316830 200841
rect 316774 200767 316830 200776
rect 316682 189816 316738 189825
rect 316682 189751 316738 189760
rect 316132 175976 316184 175982
rect 316132 175918 316184 175924
rect 316040 131096 316092 131102
rect 316040 131038 316092 131044
rect 316040 34536 316092 34542
rect 316040 34478 316092 34484
rect 315304 4140 315356 4146
rect 315304 4082 315356 4088
rect 316052 3534 316080 34478
rect 316696 14521 316724 189751
rect 316788 35902 316816 200767
rect 317524 161430 317552 238750
rect 317512 161424 317564 161430
rect 317512 161366 317564 161372
rect 317616 151814 317644 322186
rect 318076 280838 318104 369106
rect 319456 358086 319484 373966
rect 319444 358080 319496 358086
rect 319444 358022 319496 358028
rect 318064 280832 318116 280838
rect 318064 280774 318116 280780
rect 318800 280220 318852 280226
rect 318800 280162 318852 280168
rect 318064 260840 318116 260846
rect 318064 260782 318116 260788
rect 318076 156670 318104 260782
rect 318064 156664 318116 156670
rect 318064 156606 318116 156612
rect 317616 151786 317736 151814
rect 317420 140888 317472 140894
rect 317420 140830 317472 140836
rect 316776 35896 316828 35902
rect 316776 35838 316828 35844
rect 316788 34542 316816 35838
rect 316776 34536 316828 34542
rect 316776 34478 316828 34484
rect 317432 16574 317460 140830
rect 317708 140078 317736 151786
rect 318812 140758 318840 280162
rect 319442 243536 319498 243545
rect 319442 243471 319498 243480
rect 319456 152522 319484 243471
rect 320192 221921 320220 375294
rect 320284 349081 320312 377590
rect 322204 360936 322256 360942
rect 322204 360878 322256 360884
rect 320270 349072 320326 349081
rect 320270 349007 320326 349016
rect 320822 349072 320878 349081
rect 320822 349007 320878 349016
rect 320836 347857 320864 349007
rect 320822 347848 320878 347857
rect 320822 347783 320878 347792
rect 320178 221912 320234 221921
rect 320178 221847 320234 221856
rect 320638 221912 320694 221921
rect 320638 221847 320694 221856
rect 320652 221474 320680 221847
rect 320640 221468 320692 221474
rect 320640 221410 320692 221416
rect 319444 152516 319496 152522
rect 319444 152458 319496 152464
rect 319444 141432 319496 141438
rect 319444 141374 319496 141380
rect 318800 140752 318852 140758
rect 318800 140694 318852 140700
rect 317696 140072 317748 140078
rect 317696 140014 317748 140020
rect 318708 140072 318760 140078
rect 318708 140014 318760 140020
rect 318720 139466 318748 140014
rect 318708 139460 318760 139466
rect 318708 139402 318760 139408
rect 319456 16574 319484 141374
rect 320836 37262 320864 347783
rect 322216 347070 322244 360878
rect 322204 347064 322256 347070
rect 322204 347006 322256 347012
rect 322204 329112 322256 329118
rect 322204 329054 322256 329060
rect 322216 302938 322244 329054
rect 322204 302932 322256 302938
rect 322204 302874 322256 302880
rect 322202 298208 322258 298217
rect 322202 298143 322258 298152
rect 322216 273970 322244 298143
rect 322296 289876 322348 289882
rect 322296 289818 322348 289824
rect 322204 273964 322256 273970
rect 322204 273906 322256 273912
rect 322204 254652 322256 254658
rect 322204 254594 322256 254600
rect 320914 205048 320970 205057
rect 320914 204983 320970 204992
rect 320928 117298 320956 204983
rect 320916 117292 320968 117298
rect 320916 117234 320968 117240
rect 322216 93838 322244 254594
rect 322308 239465 322336 289818
rect 322952 239494 322980 377604
rect 324332 377590 324622 377618
rect 326278 377590 326384 377618
rect 324332 345681 324360 377590
rect 325608 374060 325660 374066
rect 325608 374002 325660 374008
rect 324318 345672 324374 345681
rect 324318 345607 324374 345616
rect 324962 308408 325018 308417
rect 324962 308343 325018 308352
rect 323674 277536 323730 277545
rect 323674 277471 323730 277480
rect 322940 239488 322992 239494
rect 322294 239456 322350 239465
rect 322940 239430 322992 239436
rect 322294 239391 322350 239400
rect 322294 237416 322350 237425
rect 322294 237351 322350 237360
rect 322308 158030 322336 237351
rect 323582 224224 323638 224233
rect 323582 224159 323638 224168
rect 322296 158024 322348 158030
rect 322296 157966 322348 157972
rect 322296 138100 322348 138106
rect 322296 138042 322348 138048
rect 322204 93832 322256 93838
rect 322204 93774 322256 93780
rect 321560 50380 321612 50386
rect 321560 50322 321612 50328
rect 320824 37256 320876 37262
rect 320824 37198 320876 37204
rect 320836 36922 320864 37198
rect 320180 36916 320232 36922
rect 320180 36858 320232 36864
rect 320824 36916 320876 36922
rect 320824 36858 320876 36864
rect 320192 16574 320220 36858
rect 321572 16574 321600 50322
rect 317432 16546 318104 16574
rect 319456 16546 319760 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 316682 14512 316738 14521
rect 316682 14447 316738 14456
rect 316040 3528 316092 3534
rect 316040 3470 316092 3476
rect 314856 598 315068 626
rect 314856 490 314884 598
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 462 314884 490
rect 315040 480 315068 598
rect 316236 598 316448 626
rect 316236 480 316264 598
rect 316420 490 316448 598
rect 316696 490 316724 14447
rect 317328 3528 317380 3534
rect 317328 3470 317380 3476
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 316420 462 316724 490
rect 317340 480 317368 3470
rect 318076 490 318104 16546
rect 319732 4146 319760 16546
rect 319720 4140 319772 4146
rect 319720 4082 319772 4088
rect 318352 598 318564 626
rect 318352 490 318380 598
rect 317298 -960 317410 480
rect 318076 462 318380 490
rect 318536 480 318564 598
rect 319732 480 319760 4082
rect 320468 490 320496 16546
rect 320744 598 320956 626
rect 320744 490 320772 598
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 322124 480 322152 16546
rect 322308 3777 322336 138042
rect 323596 19378 323624 224159
rect 323688 200802 323716 277471
rect 324320 234592 324372 234598
rect 324318 234560 324320 234569
rect 324372 234560 324374 234569
rect 324318 234495 324374 234504
rect 323676 200796 323728 200802
rect 323676 200738 323728 200744
rect 324976 108361 325004 308343
rect 325620 234598 325648 374002
rect 326356 337385 326384 377590
rect 327920 374066 327948 377604
rect 328472 377590 329590 377618
rect 327908 374060 327960 374066
rect 327908 374002 327960 374008
rect 328472 351937 328500 377590
rect 331232 365022 331260 377604
rect 332612 377590 332902 377618
rect 333992 377590 334558 377618
rect 335372 377590 336214 377618
rect 336752 377590 337870 377618
rect 331864 366444 331916 366450
rect 331864 366386 331916 366392
rect 331220 365016 331272 365022
rect 331220 364958 331272 364964
rect 331876 354657 331904 366386
rect 331862 354648 331918 354657
rect 331862 354583 331918 354592
rect 328458 351928 328514 351937
rect 328458 351863 328514 351872
rect 329102 351928 329158 351937
rect 329102 351863 329158 351872
rect 326342 337376 326398 337385
rect 326342 337311 326398 337320
rect 327722 337376 327778 337385
rect 327722 337311 327778 337320
rect 326988 322244 327040 322250
rect 326988 322186 327040 322192
rect 327000 321638 327028 322186
rect 325700 321632 325752 321638
rect 325700 321574 325752 321580
rect 326988 321632 327040 321638
rect 326988 321574 327040 321580
rect 325608 234592 325660 234598
rect 325608 234534 325660 234540
rect 325056 219496 325108 219502
rect 325056 219438 325108 219444
rect 324962 108352 325018 108361
rect 324962 108287 325018 108296
rect 325068 102814 325096 219438
rect 325712 132462 325740 321574
rect 327736 301578 327764 337311
rect 327816 319456 327868 319462
rect 327816 319398 327868 319404
rect 327724 301572 327776 301578
rect 327724 301514 327776 301520
rect 327724 234592 327776 234598
rect 327724 234534 327776 234540
rect 327736 137970 327764 234534
rect 327828 228410 327856 319398
rect 327816 228404 327868 228410
rect 327816 228346 327868 228352
rect 327724 137964 327776 137970
rect 327724 137906 327776 137912
rect 327078 135960 327134 135969
rect 327078 135895 327134 135904
rect 328366 135960 328422 135969
rect 328366 135895 328368 135904
rect 325700 132456 325752 132462
rect 325700 132398 325752 132404
rect 325056 102808 325108 102814
rect 325056 102750 325108 102756
rect 326342 89040 326398 89049
rect 326342 88975 326398 88984
rect 324964 83496 325016 83502
rect 324964 83438 325016 83444
rect 323676 66904 323728 66910
rect 323676 66846 323728 66852
rect 323584 19372 323636 19378
rect 323584 19314 323636 19320
rect 323596 6914 323624 19314
rect 323320 6886 323624 6914
rect 322294 3768 322350 3777
rect 322294 3703 322350 3712
rect 323320 480 323348 6886
rect 323688 3466 323716 66846
rect 324976 26217 325004 83438
rect 325054 37904 325110 37913
rect 325054 37839 325110 37848
rect 324410 26208 324466 26217
rect 324410 26143 324466 26152
rect 324962 26208 325018 26217
rect 324962 26143 325018 26152
rect 324424 3534 324452 26143
rect 325068 6866 325096 37839
rect 325056 6860 325108 6866
rect 325056 6802 325108 6808
rect 325068 5574 325096 6802
rect 324504 5568 324556 5574
rect 324504 5510 324556 5516
rect 325056 5568 325108 5574
rect 325056 5510 325108 5516
rect 324412 3528 324464 3534
rect 324412 3470 324464 3476
rect 323676 3460 323728 3466
rect 323676 3402 323728 3408
rect 324516 3346 324544 5510
rect 326356 4146 326384 88975
rect 327092 28286 327120 135895
rect 328420 135895 328422 135904
rect 328368 135866 328420 135872
rect 329116 101454 329144 351863
rect 330484 301572 330536 301578
rect 330484 301514 330536 301520
rect 329104 101448 329156 101454
rect 329104 101390 329156 101396
rect 329102 68232 329158 68241
rect 329102 68167 329158 68176
rect 327080 28280 327132 28286
rect 327080 28222 327132 28228
rect 327080 24200 327132 24206
rect 327080 24142 327132 24148
rect 327092 19378 327120 24142
rect 327080 19372 327132 19378
rect 327080 19314 327132 19320
rect 328000 8968 328052 8974
rect 328000 8910 328052 8916
rect 326344 4140 326396 4146
rect 326344 4082 326396 4088
rect 326804 4140 326856 4146
rect 326804 4082 326856 4088
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 324424 3318 324544 3346
rect 324424 480 324452 3318
rect 325620 480 325648 3470
rect 326816 480 326844 4082
rect 328012 480 328040 8910
rect 329116 4146 329144 68167
rect 330496 67726 330524 301514
rect 331876 80034 331904 354583
rect 332612 288454 332640 377590
rect 332600 288448 332652 288454
rect 332598 288416 332600 288425
rect 332652 288416 332654 288425
rect 332598 288351 332654 288360
rect 332598 284336 332654 284345
rect 332598 284271 332600 284280
rect 332652 284271 332654 284280
rect 333888 284300 333940 284306
rect 332600 284242 332652 284248
rect 333888 284242 333940 284248
rect 333900 175982 333928 284242
rect 333992 236706 334020 377590
rect 335372 332586 335400 377590
rect 336752 366382 336780 377590
rect 339512 375329 339540 377604
rect 340892 377590 341182 377618
rect 342272 377590 342838 377618
rect 344020 377590 344494 377618
rect 345032 377590 346150 377618
rect 339498 375320 339554 375329
rect 339498 375255 339554 375264
rect 338764 374740 338816 374746
rect 338764 374682 338816 374688
rect 336740 366376 336792 366382
rect 336740 366318 336792 366324
rect 337382 358048 337438 358057
rect 337382 357983 337438 357992
rect 336002 354784 336058 354793
rect 336002 354719 336058 354728
rect 335360 332580 335412 332586
rect 335360 332522 335412 332528
rect 334806 283520 334862 283529
rect 334806 283455 334862 283464
rect 333980 236700 334032 236706
rect 333980 236642 334032 236648
rect 334624 225616 334676 225622
rect 334624 225558 334676 225564
rect 333888 175976 333940 175982
rect 333888 175918 333940 175924
rect 331220 80028 331272 80034
rect 331220 79970 331272 79976
rect 331864 80028 331916 80034
rect 331864 79970 331916 79976
rect 330484 67720 330536 67726
rect 330484 67662 330536 67668
rect 329196 7676 329248 7682
rect 329196 7618 329248 7624
rect 329104 4140 329156 4146
rect 329104 4082 329156 4088
rect 329208 480 329236 7618
rect 330496 6914 330524 67662
rect 330404 6886 330524 6914
rect 330404 480 330432 6886
rect 331232 490 331260 79970
rect 332600 76560 332652 76566
rect 332600 76502 332652 76508
rect 332612 3534 332640 76502
rect 334636 67658 334664 225558
rect 334714 184376 334770 184385
rect 334714 184311 334770 184320
rect 334624 67652 334676 67658
rect 334624 67594 334676 67600
rect 334636 9654 334664 67594
rect 334728 20670 334756 184311
rect 334820 184210 334848 283455
rect 334808 184204 334860 184210
rect 334808 184146 334860 184152
rect 336016 129062 336044 354719
rect 336096 267028 336148 267034
rect 336096 266970 336148 266976
rect 336004 129056 336056 129062
rect 336004 128998 336056 129004
rect 336108 99414 336136 266970
rect 336096 99408 336148 99414
rect 336096 99350 336148 99356
rect 337396 74534 337424 357983
rect 338776 312594 338804 374682
rect 340892 366382 340920 377590
rect 342168 374672 342220 374678
rect 342168 374614 342220 374620
rect 340880 366376 340932 366382
rect 340880 366318 340932 366324
rect 340236 365016 340288 365022
rect 340236 364958 340288 364964
rect 338856 347064 338908 347070
rect 338856 347006 338908 347012
rect 338764 312588 338816 312594
rect 338764 312530 338816 312536
rect 338762 285696 338818 285705
rect 338762 285631 338818 285640
rect 338776 144226 338804 285631
rect 338868 276010 338896 347006
rect 340142 329896 340198 329905
rect 340142 329831 340198 329840
rect 338856 276004 338908 276010
rect 338856 275946 338908 275952
rect 338854 215928 338910 215937
rect 338854 215863 338910 215872
rect 338764 144220 338816 144226
rect 338764 144162 338816 144168
rect 338868 120086 338896 215863
rect 338856 120080 338908 120086
rect 338856 120022 338908 120028
rect 338120 117564 338172 117570
rect 338120 117506 338172 117512
rect 337396 74506 337516 74534
rect 335360 73840 335412 73846
rect 335360 73782 335412 73788
rect 335372 67726 335400 73782
rect 336740 69692 336792 69698
rect 336740 69634 336792 69640
rect 335360 67720 335412 67726
rect 335360 67662 335412 67668
rect 336752 67658 336780 69634
rect 336740 67652 336792 67658
rect 336740 67594 336792 67600
rect 337488 67590 337516 74506
rect 337476 67584 337528 67590
rect 337476 67526 337528 67532
rect 337488 66910 337516 67526
rect 337476 66904 337528 66910
rect 337476 66846 337528 66852
rect 335360 54528 335412 54534
rect 335360 54470 335412 54476
rect 334716 20664 334768 20670
rect 334716 20606 334768 20612
rect 335268 20664 335320 20670
rect 335268 20606 335320 20612
rect 334624 9648 334676 9654
rect 334624 9590 334676 9596
rect 332692 9036 332744 9042
rect 332692 8978 332744 8984
rect 332600 3528 332652 3534
rect 332600 3470 332652 3476
rect 331416 598 331628 626
rect 331416 490 331444 598
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 462 331444 490
rect 331600 480 331628 598
rect 332704 480 332732 8978
rect 335280 6914 335308 20606
rect 335372 16574 335400 54470
rect 338132 16574 338160 117506
rect 340156 53310 340184 329831
rect 340248 322250 340276 364958
rect 341522 362264 341578 362273
rect 341522 362199 341578 362208
rect 340236 322244 340288 322250
rect 340236 322186 340288 322192
rect 340880 317552 340932 317558
rect 340880 317494 340932 317500
rect 340892 317393 340920 317494
rect 340878 317384 340934 317393
rect 340878 317319 340934 317328
rect 340234 126304 340290 126313
rect 340234 126239 340290 126248
rect 340248 117570 340276 126239
rect 340236 117564 340288 117570
rect 340236 117506 340288 117512
rect 340788 53780 340840 53786
rect 340788 53722 340840 53728
rect 340800 53310 340828 53722
rect 340144 53304 340196 53310
rect 340144 53246 340196 53252
rect 340788 53304 340840 53310
rect 340788 53246 340840 53252
rect 335372 16546 336320 16574
rect 338132 16546 338712 16574
rect 335096 6886 335308 6914
rect 333888 3528 333940 3534
rect 333888 3470 333940 3476
rect 333900 480 333928 3470
rect 335096 480 335124 6886
rect 336292 480 336320 16546
rect 337476 9648 337528 9654
rect 337476 9590 337528 9596
rect 337488 480 337516 9590
rect 338684 480 338712 16546
rect 340800 3534 340828 53246
rect 341536 15910 341564 362199
rect 342180 317558 342208 374614
rect 342168 317552 342220 317558
rect 342168 317494 342220 317500
rect 342272 239426 342300 377590
rect 344020 376961 344048 377590
rect 344006 376952 344062 376961
rect 344006 376887 344062 376896
rect 342902 375320 342958 375329
rect 342902 375255 342958 375264
rect 342916 374785 342944 375255
rect 342902 374776 342958 374785
rect 342902 374711 342958 374720
rect 342260 239420 342312 239426
rect 342260 239362 342312 239368
rect 342916 237289 342944 374711
rect 344020 373994 344048 376887
rect 343652 373966 344048 373994
rect 343652 343602 343680 373966
rect 345032 360874 345060 377590
rect 345756 376100 345808 376106
rect 345756 376042 345808 376048
rect 345020 360868 345072 360874
rect 345020 360810 345072 360816
rect 343640 343596 343692 343602
rect 343640 343538 343692 343544
rect 344284 326392 344336 326398
rect 344284 326334 344336 326340
rect 342994 239456 343050 239465
rect 342994 239391 343050 239400
rect 342902 237280 342958 237289
rect 342902 237215 342958 237224
rect 342916 236706 342944 237215
rect 342904 236700 342956 236706
rect 342904 236642 342956 236648
rect 341614 234696 341670 234705
rect 341614 234631 341670 234640
rect 341628 163538 341656 234631
rect 342904 221536 342956 221542
rect 342904 221478 342956 221484
rect 341616 163532 341668 163538
rect 341616 163474 341668 163480
rect 342916 133890 342944 221478
rect 343008 170406 343036 239391
rect 342996 170400 343048 170406
rect 342996 170342 343048 170348
rect 342994 140040 343050 140049
rect 342994 139975 343050 139984
rect 342904 133884 342956 133890
rect 342904 133826 342956 133832
rect 343008 57322 343036 139975
rect 343548 82136 343600 82142
rect 343548 82078 343600 82084
rect 342996 57316 343048 57322
rect 342996 57258 343048 57264
rect 341524 15904 341576 15910
rect 341524 15846 341576 15852
rect 342352 15904 342404 15910
rect 342352 15846 342404 15852
rect 342364 3534 342392 15846
rect 343560 6914 343588 82078
rect 344296 72486 344324 326334
rect 345664 251932 345716 251938
rect 345664 251874 345716 251880
rect 344284 72480 344336 72486
rect 344284 72422 344336 72428
rect 344296 16574 344324 72422
rect 345676 16574 345704 251874
rect 345768 242214 345796 376042
rect 347792 374746 347820 377604
rect 349172 377590 349462 377618
rect 348422 376544 348478 376553
rect 348422 376479 348478 376488
rect 347780 374740 347832 374746
rect 347780 374682 347832 374688
rect 347044 370592 347096 370598
rect 347044 370534 347096 370540
rect 347056 317490 347084 370534
rect 348436 334694 348464 376479
rect 349172 340202 349200 377590
rect 351104 374649 351132 377604
rect 352562 377496 352618 377505
rect 352562 377431 352618 377440
rect 351184 375352 351236 375358
rect 351184 375294 351236 375300
rect 351090 374640 351146 374649
rect 351090 374575 351146 374584
rect 349804 373380 349856 373386
rect 349804 373322 349856 373328
rect 349160 340196 349212 340202
rect 349160 340138 349212 340144
rect 348424 334688 348476 334694
rect 348424 334630 348476 334636
rect 347044 317484 347096 317490
rect 347044 317426 347096 317432
rect 345756 242208 345808 242214
rect 345756 242150 345808 242156
rect 345754 211984 345810 211993
rect 345754 211919 345810 211928
rect 345768 130422 345796 211919
rect 345756 130416 345808 130422
rect 345756 130358 345808 130364
rect 347056 104854 347084 317426
rect 348424 257440 348476 257446
rect 348424 257382 348476 257388
rect 347044 104848 347096 104854
rect 347044 104790 347096 104796
rect 346400 57248 346452 57254
rect 346400 57190 346452 57196
rect 346412 16574 346440 57190
rect 348436 16574 348464 257382
rect 349816 222902 349844 373322
rect 351196 356697 351224 375294
rect 351182 356688 351238 356697
rect 351182 356623 351238 356632
rect 350446 346488 350502 346497
rect 350446 346423 350502 346432
rect 350460 346390 350488 346423
rect 352576 346390 352604 377431
rect 352760 374678 352788 377604
rect 354128 377460 354180 377466
rect 354128 377402 354180 377408
rect 353942 376000 353998 376009
rect 353942 375935 353998 375944
rect 352748 374672 352800 374678
rect 352748 374614 352800 374620
rect 352656 373312 352708 373318
rect 352656 373254 352708 373260
rect 350448 346384 350500 346390
rect 350448 346326 350500 346332
rect 352564 346384 352616 346390
rect 352564 346326 352616 346332
rect 349804 222896 349856 222902
rect 349804 222838 349856 222844
rect 349802 142216 349858 142225
rect 349802 142151 349858 142160
rect 344296 16546 344600 16574
rect 345676 16546 345796 16574
rect 346412 16546 346992 16574
rect 343376 6886 343588 6914
rect 339868 3528 339920 3534
rect 339868 3470 339920 3476
rect 340788 3528 340840 3534
rect 340788 3470 340840 3476
rect 340972 3528 341024 3534
rect 340972 3470 341024 3476
rect 342352 3528 342404 3534
rect 342352 3470 342404 3476
rect 339880 480 339908 3470
rect 340984 480 341012 3470
rect 342166 3360 342222 3369
rect 342166 3295 342222 3304
rect 342180 480 342208 3295
rect 343376 480 343404 6886
rect 344572 480 344600 16546
rect 345768 4078 345796 16546
rect 345756 4072 345808 4078
rect 345756 4014 345808 4020
rect 345768 480 345796 4014
rect 346964 480 346992 16546
rect 348068 16546 348464 16574
rect 348068 12442 348096 16546
rect 348056 12436 348108 12442
rect 348056 12378 348108 12384
rect 348068 480 348096 12378
rect 349816 12374 349844 142151
rect 349804 12368 349856 12374
rect 349804 12310 349856 12316
rect 350460 9654 350488 346326
rect 352562 306504 352618 306513
rect 352562 306439 352618 306448
rect 351182 195256 351238 195265
rect 351182 195191 351238 195200
rect 349988 9648 350040 9654
rect 349988 9590 350040 9596
rect 350448 9648 350500 9654
rect 350448 9590 350500 9596
rect 350000 9042 350028 9590
rect 349988 9036 350040 9042
rect 349988 8978 350040 8984
rect 351196 3670 351224 195191
rect 352576 114510 352604 306439
rect 352668 245002 352696 373254
rect 353956 354686 353984 375935
rect 354034 374096 354090 374105
rect 354034 374031 354090 374040
rect 353944 354680 353996 354686
rect 353944 354622 353996 354628
rect 353944 301504 353996 301510
rect 353944 301446 353996 301452
rect 352656 244996 352708 245002
rect 352656 244938 352708 244944
rect 352654 232520 352710 232529
rect 352654 232455 352710 232464
rect 352668 118658 352696 232455
rect 352746 124128 352802 124137
rect 352746 124063 352802 124072
rect 352656 118652 352708 118658
rect 352656 118594 352708 118600
rect 352564 114504 352616 114510
rect 352564 114446 352616 114452
rect 352562 90400 352618 90409
rect 352562 90335 352618 90344
rect 351642 3904 351698 3913
rect 351642 3839 351698 3848
rect 351656 3670 351684 3839
rect 351184 3664 351236 3670
rect 351184 3606 351236 3612
rect 351644 3664 351696 3670
rect 351644 3606 351696 3612
rect 350446 3496 350502 3505
rect 349252 3460 349304 3466
rect 350446 3431 350502 3440
rect 349252 3402 349304 3408
rect 349264 480 349292 3402
rect 350460 480 350488 3431
rect 351656 480 351684 3606
rect 352576 3505 352604 90335
rect 352760 64190 352788 124063
rect 353956 95198 353984 301446
rect 354048 246401 354076 374031
rect 354140 357406 354168 377402
rect 354416 375358 354444 377604
rect 354678 375728 354734 375737
rect 354678 375663 354734 375672
rect 354404 375352 354456 375358
rect 354404 375294 354456 375300
rect 354692 367713 354720 375663
rect 354678 367704 354734 367713
rect 354678 367639 354734 367648
rect 354128 357400 354180 357406
rect 354128 357342 354180 357348
rect 355324 302932 355376 302938
rect 355324 302874 355376 302880
rect 354128 274032 354180 274038
rect 354128 273974 354180 273980
rect 354034 246392 354090 246401
rect 354034 246327 354090 246336
rect 354140 171834 354168 273974
rect 354128 171828 354180 171834
rect 354128 171770 354180 171776
rect 355336 129810 355364 302874
rect 356072 250578 356100 377604
rect 356164 377505 356192 451246
rect 356242 423736 356298 423745
rect 356242 423671 356298 423680
rect 356150 377496 356206 377505
rect 356150 377431 356206 377440
rect 356256 366450 356284 423671
rect 356334 394496 356390 394505
rect 356334 394431 356390 394440
rect 356348 393378 356376 394431
rect 356336 393372 356388 393378
rect 356336 393314 356388 393320
rect 356348 371890 356376 393314
rect 356426 387152 356482 387161
rect 356426 387087 356482 387096
rect 356440 373425 356468 387087
rect 356426 373416 356482 373425
rect 356426 373351 356482 373360
rect 357452 371929 357480 458351
rect 358726 455968 358782 455977
rect 358726 455903 358782 455912
rect 358740 455462 358768 455903
rect 358728 455456 358780 455462
rect 358728 455398 358780 455404
rect 358726 453520 358782 453529
rect 358726 453455 358782 453464
rect 358740 452674 358768 453455
rect 358728 452668 358780 452674
rect 358728 452610 358780 452616
rect 358726 451072 358782 451081
rect 358726 451007 358782 451016
rect 358740 449954 358768 451007
rect 358728 449948 358780 449954
rect 358728 449890 358780 449896
rect 358726 448624 358782 448633
rect 358726 448559 358728 448568
rect 358780 448559 358782 448568
rect 358728 448530 358780 448536
rect 358726 446176 358782 446185
rect 358726 446111 358782 446120
rect 358740 445806 358768 446111
rect 358728 445800 358780 445806
rect 358728 445742 358780 445748
rect 358726 443728 358782 443737
rect 358726 443663 358782 443672
rect 358740 443018 358768 443663
rect 358728 443012 358780 443018
rect 358728 442954 358780 442960
rect 358726 438968 358782 438977
rect 358726 438903 358728 438912
rect 358780 438903 358782 438912
rect 358728 438874 358780 438880
rect 358726 436384 358782 436393
rect 358726 436319 358782 436328
rect 358740 436150 358768 436319
rect 358728 436144 358780 436150
rect 358728 436086 358780 436092
rect 358726 433936 358782 433945
rect 358726 433871 358782 433880
rect 358740 433362 358768 433871
rect 358728 433356 358780 433362
rect 358728 433298 358780 433304
rect 358726 429040 358782 429049
rect 358726 428975 358782 428984
rect 358740 427854 358768 428975
rect 358728 427848 358780 427854
rect 358728 427790 358780 427796
rect 358726 426592 358782 426601
rect 358726 426527 358782 426536
rect 358740 426494 358768 426527
rect 358728 426488 358780 426494
rect 358728 426430 358780 426436
rect 357530 421696 357586 421705
rect 357530 421631 357586 421640
rect 357438 371920 357494 371929
rect 356336 371884 356388 371890
rect 357438 371855 357494 371864
rect 356336 371826 356388 371832
rect 356794 370560 356850 370569
rect 356794 370495 356850 370504
rect 356244 366444 356296 366450
rect 356244 366386 356296 366392
rect 356704 355360 356756 355366
rect 356704 355302 356756 355308
rect 356716 320210 356744 355302
rect 356808 347070 356836 370495
rect 357544 358057 357572 421631
rect 358726 419248 358782 419257
rect 358726 419183 358782 419192
rect 358740 418198 358768 419183
rect 358728 418192 358780 418198
rect 358728 418134 358780 418140
rect 358728 416832 358780 416838
rect 358726 416800 358728 416809
rect 358780 416800 358782 416809
rect 358726 416735 358782 416744
rect 358726 414352 358782 414361
rect 358726 414287 358782 414296
rect 358740 414050 358768 414287
rect 358728 414044 358780 414050
rect 358728 413986 358780 413992
rect 358726 411904 358782 411913
rect 358726 411839 358782 411848
rect 358740 411330 358768 411839
rect 358728 411324 358780 411330
rect 358728 411266 358780 411272
rect 358726 407008 358782 407017
rect 358726 406943 358782 406952
rect 358740 405754 358768 406943
rect 358728 405748 358780 405754
rect 358728 405690 358780 405696
rect 358726 404288 358782 404297
rect 358726 404223 358782 404232
rect 358740 403034 358768 404223
rect 358728 403028 358780 403034
rect 358728 402970 358780 402976
rect 358726 401840 358782 401849
rect 358726 401775 358782 401784
rect 358740 401674 358768 401775
rect 358728 401668 358780 401674
rect 358728 401610 358780 401616
rect 358634 399392 358690 399401
rect 358634 399327 358690 399336
rect 358648 398886 358676 399327
rect 358636 398880 358688 398886
rect 358636 398822 358688 398828
rect 357622 392048 357678 392057
rect 357622 391983 357678 391992
rect 357636 370530 357664 391983
rect 357714 389600 357770 389609
rect 357714 389535 357770 389544
rect 357728 376106 357756 389535
rect 357898 384704 357954 384713
rect 357898 384639 357954 384648
rect 357912 383722 357940 384639
rect 357900 383716 357952 383722
rect 357900 383658 357952 383664
rect 357898 379808 357954 379817
rect 357898 379743 357954 379752
rect 357912 379574 357940 379743
rect 357900 379568 357952 379574
rect 357900 379510 357952 379516
rect 357716 376100 357768 376106
rect 357716 376042 357768 376048
rect 358082 371376 358138 371385
rect 358082 371311 358138 371320
rect 357624 370524 357676 370530
rect 357624 370466 357676 370472
rect 357530 358048 357586 358057
rect 357530 357983 357586 357992
rect 358096 349858 358124 371311
rect 358176 358080 358228 358086
rect 358176 358022 358228 358028
rect 358084 349852 358136 349858
rect 358084 349794 358136 349800
rect 356796 347064 356848 347070
rect 356796 347006 356848 347012
rect 356704 320204 356756 320210
rect 356704 320146 356756 320152
rect 356716 286142 356744 320146
rect 358084 304292 358136 304298
rect 358084 304234 358136 304240
rect 356704 286136 356756 286142
rect 356704 286078 356756 286084
rect 356796 262268 356848 262274
rect 356796 262210 356848 262216
rect 356060 250572 356112 250578
rect 356060 250514 356112 250520
rect 356704 210452 356756 210458
rect 356704 210394 356756 210400
rect 355324 129804 355376 129810
rect 355324 129746 355376 129752
rect 354034 124128 354090 124137
rect 354034 124063 354090 124072
rect 354048 123486 354076 124063
rect 354036 123480 354088 123486
rect 354036 123422 354088 123428
rect 354036 109064 354088 109070
rect 354036 109006 354088 109012
rect 353944 95192 353996 95198
rect 353944 95134 353996 95140
rect 352748 64184 352800 64190
rect 352748 64126 352800 64132
rect 354048 7614 354076 109006
rect 356716 97986 356744 210394
rect 356808 160750 356836 262210
rect 356796 160744 356848 160750
rect 356796 160686 356848 160692
rect 358096 155242 358124 304234
rect 358188 284306 358216 358022
rect 358832 313954 358860 538290
rect 358912 535560 358964 535566
rect 358912 535502 358964 535508
rect 358924 348430 358952 535502
rect 359016 532030 359044 560254
rect 360292 545148 360344 545154
rect 360292 545090 360344 545096
rect 360200 541680 360252 541686
rect 360200 541622 360252 541628
rect 359004 532024 359056 532030
rect 359004 531966 359056 531972
rect 360212 496806 360240 541622
rect 360200 496800 360252 496806
rect 360200 496742 360252 496748
rect 360200 473340 360252 473346
rect 360200 473282 360252 473288
rect 359094 441280 359150 441289
rect 359094 441215 359150 441224
rect 359002 431488 359058 431497
rect 359002 431423 359058 431432
rect 358912 348424 358964 348430
rect 358912 348366 358964 348372
rect 358820 313948 358872 313954
rect 358820 313890 358872 313896
rect 358176 284300 358228 284306
rect 358176 284242 358228 284248
rect 358176 266348 358228 266354
rect 358176 266290 358228 266296
rect 358084 155236 358136 155242
rect 358084 155178 358136 155184
rect 358082 137728 358138 137737
rect 358082 137663 358138 137672
rect 356704 97980 356756 97986
rect 356704 97922 356756 97928
rect 354036 7608 354088 7614
rect 354036 7550 354088 7556
rect 352562 3496 352618 3505
rect 352562 3431 352618 3440
rect 358096 3369 358124 137663
rect 358188 115938 358216 266290
rect 359016 253298 359044 431423
rect 359108 369170 359136 441215
rect 359096 369164 359148 369170
rect 359096 369106 359148 369112
rect 359462 289096 359518 289105
rect 359462 289031 359518 289040
rect 359004 253292 359056 253298
rect 359004 253234 359056 253240
rect 358820 129804 358872 129810
rect 358820 129746 358872 129752
rect 358176 115932 358228 115938
rect 358176 115874 358228 115880
rect 358832 8974 358860 129746
rect 359476 103494 359504 289031
rect 360212 276690 360240 473282
rect 360304 377466 360332 545090
rect 360856 543833 360884 702578
rect 376116 700324 376168 700330
rect 376116 700266 376168 700272
rect 367100 545216 367152 545222
rect 367100 545158 367152 545164
rect 360842 543824 360898 543833
rect 360842 543759 360898 543768
rect 363052 543788 363104 543794
rect 363052 543730 363104 543736
rect 361580 539708 361632 539714
rect 361580 539650 361632 539656
rect 360384 462392 360436 462398
rect 360384 462334 360436 462340
rect 360292 377460 360344 377466
rect 360292 377402 360344 377408
rect 360396 363662 360424 462334
rect 360476 379568 360528 379574
rect 360476 379510 360528 379516
rect 360488 373386 360516 379510
rect 360476 373380 360528 373386
rect 360476 373322 360528 373328
rect 360384 363656 360436 363662
rect 360384 363598 360436 363604
rect 360200 276684 360252 276690
rect 360200 276626 360252 276632
rect 360934 143576 360990 143585
rect 360934 143511 360990 143520
rect 359464 103488 359516 103494
rect 359464 103430 359516 103436
rect 360844 101448 360896 101454
rect 360844 101390 360896 101396
rect 360856 89690 360884 101390
rect 360844 89684 360896 89690
rect 360844 89626 360896 89632
rect 358820 8968 358872 8974
rect 358820 8910 358872 8916
rect 360856 3466 360884 89626
rect 360948 80714 360976 143511
rect 361592 120057 361620 539650
rect 362958 538520 363014 538529
rect 362958 538455 363014 538464
rect 361672 443012 361724 443018
rect 361672 442954 361724 442960
rect 361684 258806 361712 442954
rect 361764 418192 361816 418198
rect 361764 418134 361816 418140
rect 361776 360942 361804 418134
rect 361856 398880 361908 398886
rect 361856 398822 361908 398828
rect 361868 376009 361896 398822
rect 361854 376000 361910 376009
rect 361854 375935 361910 375944
rect 361764 360936 361816 360942
rect 361764 360878 361816 360884
rect 362972 327758 363000 538455
rect 363064 352578 363092 543730
rect 364432 536920 364484 536926
rect 364432 536862 364484 536868
rect 363604 516180 363656 516186
rect 363604 516122 363656 516128
rect 363616 497486 363644 516122
rect 364340 502444 364392 502450
rect 364340 502386 364392 502392
rect 363604 497480 363656 497486
rect 363604 497422 363656 497428
rect 363144 436144 363196 436150
rect 363144 436086 363196 436092
rect 363052 352572 363104 352578
rect 363052 352514 363104 352520
rect 362960 327752 363012 327758
rect 362960 327694 363012 327700
rect 361672 258800 361724 258806
rect 361672 258742 361724 258748
rect 363156 256018 363184 436086
rect 363236 427848 363288 427854
rect 363236 427790 363288 427796
rect 363248 305658 363276 427790
rect 363236 305652 363288 305658
rect 363236 305594 363288 305600
rect 364352 287706 364380 502386
rect 364444 370569 364472 536862
rect 365720 477556 365772 477562
rect 365720 477498 365772 477504
rect 364524 405748 364576 405754
rect 364524 405690 364576 405696
rect 364430 370560 364486 370569
rect 364430 370495 364486 370504
rect 364536 351898 364564 405690
rect 364524 351892 364576 351898
rect 364524 351834 364576 351840
rect 365732 291825 365760 477498
rect 365812 433356 365864 433362
rect 365812 433298 365864 433304
rect 365824 370598 365852 433298
rect 365904 403028 365956 403034
rect 365904 402970 365956 402976
rect 365916 373318 365944 402970
rect 365904 373312 365956 373318
rect 365904 373254 365956 373260
rect 365812 370592 365864 370598
rect 365812 370534 365864 370540
rect 367112 304978 367140 545158
rect 367376 541000 367428 541006
rect 367376 540942 367428 540948
rect 367284 528624 367336 528630
rect 367284 528566 367336 528572
rect 367192 481704 367244 481710
rect 367192 481646 367244 481652
rect 367100 304972 367152 304978
rect 367100 304914 367152 304920
rect 365718 291816 365774 291825
rect 365718 291751 365774 291760
rect 364340 287700 364392 287706
rect 364340 287642 364392 287648
rect 363604 286136 363656 286142
rect 363604 286078 363656 286084
rect 363144 256012 363196 256018
rect 363144 255954 363196 255960
rect 363616 135250 363644 286078
rect 366362 282160 366418 282169
rect 366362 282095 366418 282104
rect 363696 236700 363748 236706
rect 363696 236642 363748 236648
rect 363604 135244 363656 135250
rect 363604 135186 363656 135192
rect 361578 120048 361634 120057
rect 361578 119983 361634 119992
rect 361592 119377 361620 119983
rect 361578 119368 361634 119377
rect 361578 119303 361634 119312
rect 363708 101590 363736 236642
rect 363696 101584 363748 101590
rect 363696 101526 363748 101532
rect 366376 88262 366404 282095
rect 367204 268394 367232 481646
rect 367296 337414 367324 528566
rect 367388 365022 367416 540942
rect 369860 538280 369912 538286
rect 369860 538222 369912 538228
rect 368572 474768 368624 474774
rect 368572 474710 368624 474716
rect 368480 416832 368532 416838
rect 368480 416774 368532 416780
rect 367376 365016 367428 365022
rect 367376 364958 367428 364964
rect 367284 337408 367336 337414
rect 367284 337350 367336 337356
rect 367744 269816 367796 269822
rect 367744 269758 367796 269764
rect 367192 268388 367244 268394
rect 367192 268330 367244 268336
rect 367756 149734 367784 269758
rect 368492 250510 368520 416774
rect 368584 359514 368612 474710
rect 368572 359508 368624 359514
rect 368572 359450 368624 359456
rect 369872 298790 369900 538222
rect 371240 524476 371292 524482
rect 371240 524418 371292 524424
rect 369952 445800 370004 445806
rect 369952 445742 370004 445748
rect 369860 298784 369912 298790
rect 369860 298726 369912 298732
rect 369964 258738 369992 445742
rect 370044 414044 370096 414050
rect 370044 413986 370096 413992
rect 370056 372570 370084 413986
rect 370044 372564 370096 372570
rect 370044 372506 370096 372512
rect 371252 290494 371280 524418
rect 374092 472048 374144 472054
rect 374092 471990 374144 471996
rect 371424 470620 371476 470626
rect 371424 470562 371476 470568
rect 371332 448588 371384 448594
rect 371332 448530 371384 448536
rect 371344 362409 371372 448530
rect 371330 362400 371386 362409
rect 371330 362335 371386 362344
rect 371330 323640 371386 323649
rect 371330 323575 371386 323584
rect 371240 290488 371292 290494
rect 371240 290430 371292 290436
rect 370502 280800 370558 280809
rect 370502 280735 370558 280744
rect 369952 258732 370004 258738
rect 369952 258674 370004 258680
rect 368480 250504 368532 250510
rect 368480 250446 368532 250452
rect 369122 200696 369178 200705
rect 369122 200631 369178 200640
rect 367744 149728 367796 149734
rect 367744 149670 367796 149676
rect 369136 132462 369164 200631
rect 369124 132456 369176 132462
rect 369124 132398 369176 132404
rect 367836 129124 367888 129130
rect 367836 129066 367888 129072
rect 367744 121508 367796 121514
rect 367744 121450 367796 121456
rect 366916 102808 366968 102814
rect 366916 102750 366968 102756
rect 366928 95130 366956 102750
rect 366916 95124 366968 95130
rect 366916 95066 366968 95072
rect 366364 88256 366416 88262
rect 366364 88198 366416 88204
rect 360936 80708 360988 80714
rect 360936 80650 360988 80656
rect 367756 13802 367784 121450
rect 367848 106962 367876 129066
rect 367836 106956 367888 106962
rect 367836 106898 367888 106904
rect 370516 103193 370544 280735
rect 371344 132494 371372 323575
rect 371436 319462 371464 470562
rect 372988 460216 373040 460222
rect 372988 460158 373040 460164
rect 373000 459610 373028 460158
rect 372712 459604 372764 459610
rect 372712 459546 372764 459552
rect 372988 459604 373040 459610
rect 372988 459546 373040 459552
rect 371516 449200 371568 449206
rect 371516 449142 371568 449148
rect 371528 448594 371556 449142
rect 371516 448588 371568 448594
rect 371516 448530 371568 448536
rect 372620 426488 372672 426494
rect 372620 426430 372672 426436
rect 371424 319456 371476 319462
rect 371424 319398 371476 319404
rect 372632 253230 372660 426430
rect 372724 329089 372752 459546
rect 374000 449948 374052 449954
rect 374000 449890 374052 449896
rect 372710 329080 372766 329089
rect 372710 329015 372766 329024
rect 374012 260166 374040 449890
rect 374104 358086 374132 471990
rect 376024 438932 376076 438938
rect 376024 438874 376076 438880
rect 374642 373416 374698 373425
rect 374642 373351 374698 373360
rect 374092 358080 374144 358086
rect 374092 358022 374144 358028
rect 374000 260160 374052 260166
rect 374000 260102 374052 260108
rect 372620 253224 372672 253230
rect 372620 253166 372672 253172
rect 373262 231160 373318 231169
rect 373262 231095 373318 231104
rect 371884 206304 371936 206310
rect 371884 206246 371936 206252
rect 371896 166297 371924 206246
rect 371976 177336 372028 177342
rect 371976 177278 372028 177284
rect 371882 166288 371938 166297
rect 371882 166223 371938 166232
rect 371252 132466 371372 132494
rect 371252 126954 371280 132466
rect 371884 127016 371936 127022
rect 371884 126958 371936 126964
rect 371240 126948 371292 126954
rect 371240 126890 371292 126896
rect 371252 126313 371280 126890
rect 371238 126304 371294 126313
rect 371238 126239 371294 126248
rect 370596 106344 370648 106350
rect 370596 106286 370648 106292
rect 370502 103184 370558 103193
rect 370502 103119 370558 103128
rect 370608 16590 370636 106286
rect 371896 26246 371924 126958
rect 371988 99482 372016 177278
rect 371976 99476 372028 99482
rect 371976 99418 372028 99424
rect 373276 92478 373304 231095
rect 374656 105602 374684 373351
rect 374734 190496 374790 190505
rect 374734 190431 374790 190440
rect 374748 151162 374776 190431
rect 374736 151156 374788 151162
rect 374736 151098 374788 151104
rect 374736 117360 374788 117366
rect 374736 117302 374788 117308
rect 374644 105596 374696 105602
rect 374644 105538 374696 105544
rect 373264 92472 373316 92478
rect 373264 92414 373316 92420
rect 371884 26240 371936 26246
rect 371884 26182 371936 26188
rect 374748 24138 374776 117302
rect 376036 99385 376064 438874
rect 376128 376038 376156 700266
rect 379428 539640 379480 539646
rect 379428 539582 379480 539588
rect 379440 538218 379468 539582
rect 379428 538212 379480 538218
rect 379428 538154 379480 538160
rect 378140 536852 378192 536858
rect 378140 536794 378192 536800
rect 376760 455456 376812 455462
rect 376760 455398 376812 455404
rect 376116 376032 376168 376038
rect 376116 375974 376168 375980
rect 376128 287706 376156 375974
rect 376772 369073 376800 455398
rect 377404 452668 377456 452674
rect 377404 452610 377456 452616
rect 376758 369064 376814 369073
rect 376758 368999 376814 369008
rect 376116 287700 376168 287706
rect 376116 287642 376168 287648
rect 376116 133952 376168 133958
rect 376116 133894 376168 133900
rect 376022 99376 376078 99385
rect 376022 99311 376078 99320
rect 374736 24132 374788 24138
rect 374736 24074 374788 24080
rect 370596 16584 370648 16590
rect 370596 16526 370648 16532
rect 367744 13796 367796 13802
rect 367744 13738 367796 13744
rect 376128 12345 376156 133894
rect 377416 124234 377444 452610
rect 377496 264240 377548 264246
rect 377496 264182 377548 264188
rect 377404 124228 377456 124234
rect 377404 124170 377456 124176
rect 377404 106412 377456 106418
rect 377404 106354 377456 106360
rect 376114 12336 376170 12345
rect 376114 12271 376170 12280
rect 377416 9625 377444 106354
rect 377508 99346 377536 264182
rect 378152 193225 378180 536794
rect 380900 487212 380952 487218
rect 380900 487154 380952 487160
rect 379520 465112 379572 465118
rect 379520 465054 379572 465060
rect 378232 411324 378284 411330
rect 378232 411266 378284 411272
rect 378244 278050 378272 411266
rect 379532 338774 379560 465054
rect 379520 338768 379572 338774
rect 379520 338710 379572 338716
rect 380164 282940 380216 282946
rect 380164 282882 380216 282888
rect 378232 278044 378284 278050
rect 378232 277986 378284 277992
rect 378784 232552 378836 232558
rect 378784 232494 378836 232500
rect 378138 193216 378194 193225
rect 378138 193151 378194 193160
rect 378796 111790 378824 232494
rect 378874 193216 378930 193225
rect 378874 193151 378930 193160
rect 378888 132433 378916 193151
rect 378874 132424 378930 132433
rect 378874 132359 378930 132368
rect 378876 129056 378928 129062
rect 378876 128998 378928 129004
rect 378784 111784 378836 111790
rect 378784 111726 378836 111732
rect 378784 108316 378836 108322
rect 378784 108258 378836 108264
rect 377496 99340 377548 99346
rect 377496 99282 377548 99288
rect 378796 10402 378824 108258
rect 378888 93809 378916 128998
rect 380176 104145 380204 282882
rect 380912 271182 380940 487154
rect 381556 374785 381584 702646
rect 388442 541104 388498 541113
rect 388442 541039 388498 541048
rect 382280 506524 382332 506530
rect 382280 506466 382332 506472
rect 381542 374776 381598 374785
rect 381542 374711 381598 374720
rect 382292 355366 382320 506466
rect 385040 494760 385092 494766
rect 385040 494702 385092 494708
rect 382280 355360 382332 355366
rect 382280 355302 382332 355308
rect 381544 307828 381596 307834
rect 381544 307770 381596 307776
rect 380900 271176 380952 271182
rect 380900 271118 380952 271124
rect 380162 104136 380218 104145
rect 380162 104071 380218 104080
rect 381556 97753 381584 307770
rect 382924 278044 382976 278050
rect 382924 277986 382976 277992
rect 381728 164892 381780 164898
rect 381728 164834 381780 164840
rect 381634 102776 381690 102785
rect 381634 102711 381690 102720
rect 381542 97744 381598 97753
rect 381542 97679 381598 97688
rect 378874 93800 378930 93809
rect 378874 93735 378930 93744
rect 378784 10396 378836 10402
rect 378784 10338 378836 10344
rect 377402 9616 377458 9625
rect 377402 9551 377458 9560
rect 381648 7682 381676 102711
rect 381740 93770 381768 164834
rect 382936 96626 382964 277986
rect 385052 272542 385080 494702
rect 387062 312488 387118 312497
rect 387062 312423 387118 312432
rect 385040 272536 385092 272542
rect 385040 272478 385092 272484
rect 384304 254584 384356 254590
rect 384304 254526 384356 254532
rect 383014 138680 383070 138689
rect 383014 138615 383070 138624
rect 382924 96620 382976 96626
rect 382924 96562 382976 96568
rect 381728 93764 381780 93770
rect 381728 93706 381780 93712
rect 382924 54596 382976 54602
rect 382924 54538 382976 54544
rect 381636 7676 381688 7682
rect 381636 7618 381688 7624
rect 382936 4049 382964 54538
rect 383028 54534 383056 138615
rect 384316 114442 384344 254526
rect 385684 238060 385736 238066
rect 385684 238002 385736 238008
rect 385040 124228 385092 124234
rect 385040 124170 385092 124176
rect 384304 114436 384356 114442
rect 384304 114378 384356 114384
rect 383016 54528 383068 54534
rect 383016 54470 383068 54476
rect 385052 19990 385080 124170
rect 385696 124166 385724 238002
rect 385776 199436 385828 199442
rect 385776 199378 385828 199384
rect 385684 124160 385736 124166
rect 385684 124102 385736 124108
rect 385788 120018 385816 199378
rect 387076 121446 387104 312423
rect 388456 148345 388484 541039
rect 389178 535528 389234 535537
rect 389178 535463 389234 535472
rect 388536 217320 388588 217326
rect 388536 217262 388588 217268
rect 388442 148336 388498 148345
rect 388442 148271 388498 148280
rect 388444 136672 388496 136678
rect 388444 136614 388496 136620
rect 387064 121440 387116 121446
rect 387064 121382 387116 121388
rect 385776 120012 385828 120018
rect 385776 119954 385828 119960
rect 388456 40633 388484 136614
rect 388548 112470 388576 217262
rect 389192 140729 389220 535463
rect 398840 527196 398892 527202
rect 398840 527138 398892 527144
rect 395988 520940 396040 520946
rect 395988 520882 396040 520888
rect 396000 520334 396028 520882
rect 395988 520328 396040 520334
rect 395988 520270 396040 520276
rect 392216 493332 392268 493338
rect 392216 493274 392268 493280
rect 392228 492726 392256 493274
rect 392216 492720 392268 492726
rect 392216 492662 392268 492668
rect 392584 492720 392636 492726
rect 392584 492662 392636 492668
rect 392596 306374 392624 492662
rect 393320 393372 393372 393378
rect 393320 393314 393372 393320
rect 392596 306346 392716 306374
rect 392688 295322 392716 306346
rect 392676 295316 392728 295322
rect 392676 295258 392728 295264
rect 392688 294642 392716 295258
rect 392676 294636 392728 294642
rect 392676 294578 392728 294584
rect 392584 287700 392636 287706
rect 392584 287642 392636 287648
rect 389824 213240 389876 213246
rect 389824 213182 389876 213188
rect 389178 140720 389234 140729
rect 389178 140655 389234 140664
rect 389192 140049 389220 140655
rect 389178 140040 389234 140049
rect 389178 139975 389234 139984
rect 388536 112464 388588 112470
rect 388536 112406 388588 112412
rect 389836 109002 389864 213182
rect 392596 145586 392624 287642
rect 392674 192536 392730 192545
rect 392674 192471 392730 192480
rect 392584 145580 392636 145586
rect 392584 145522 392636 145528
rect 390558 132424 390614 132433
rect 390558 132359 390614 132368
rect 390572 131209 390600 132359
rect 390558 131200 390614 131209
rect 390558 131135 390614 131144
rect 391204 130416 391256 130422
rect 391204 130358 391256 130364
rect 389914 129976 389970 129985
rect 389914 129911 389970 129920
rect 389824 108996 389876 109002
rect 389824 108938 389876 108944
rect 388442 40624 388498 40633
rect 388442 40559 388498 40568
rect 389928 29646 389956 129911
rect 391216 104786 391244 130358
rect 392688 115870 392716 192471
rect 392768 170400 392820 170406
rect 392768 170342 392820 170348
rect 392676 115864 392728 115870
rect 392676 115806 392728 115812
rect 391204 104780 391256 104786
rect 391204 104722 391256 104728
rect 392584 100768 392636 100774
rect 392584 100710 392636 100716
rect 392596 37262 392624 100710
rect 392780 97918 392808 170342
rect 393332 129130 393360 393314
rect 395896 193860 395948 193866
rect 395896 193802 395948 193808
rect 393410 183016 393466 183025
rect 393410 182951 393466 182960
rect 393424 138825 393452 182951
rect 395436 160744 395488 160750
rect 395436 160686 395488 160692
rect 395342 142760 395398 142769
rect 395342 142695 395398 142704
rect 393410 138816 393466 138825
rect 393410 138751 393466 138760
rect 393410 131336 393466 131345
rect 393410 131271 393466 131280
rect 393320 129124 393372 129130
rect 393320 129066 393372 129072
rect 392768 97912 392820 97918
rect 392768 97854 392820 97860
rect 393424 76566 393452 131271
rect 394608 129124 394660 129130
rect 394608 129066 394660 129072
rect 394620 128761 394648 129066
rect 394606 128752 394662 128761
rect 394606 128687 394662 128696
rect 393964 128376 394016 128382
rect 393964 128318 394016 128324
rect 393412 76560 393464 76566
rect 393412 76502 393464 76508
rect 392584 37256 392636 37262
rect 392584 37198 392636 37204
rect 393976 32434 394004 128318
rect 393964 32428 394016 32434
rect 393964 32370 394016 32376
rect 389916 29640 389968 29646
rect 389916 29582 389968 29588
rect 395356 22846 395384 142695
rect 395448 136610 395476 160686
rect 395436 136604 395488 136610
rect 395436 136546 395488 136552
rect 395908 117298 395936 193802
rect 396000 146305 396028 520270
rect 396724 317552 396776 317558
rect 396724 317494 396776 317500
rect 396736 210361 396764 317494
rect 397366 266384 397422 266393
rect 397366 266319 397422 266328
rect 397380 262857 397408 266319
rect 396814 262848 396870 262857
rect 396814 262783 396870 262792
rect 397366 262848 397422 262857
rect 397366 262783 397422 262792
rect 396722 210352 396778 210361
rect 396722 210287 396778 210296
rect 395986 146296 396042 146305
rect 395986 146231 396042 146240
rect 396724 142248 396776 142254
rect 396724 142190 396776 142196
rect 395896 117292 395948 117298
rect 395896 117234 395948 117240
rect 395344 22840 395396 22846
rect 395344 22782 395396 22788
rect 385040 19984 385092 19990
rect 385040 19926 385092 19932
rect 396736 5506 396764 142190
rect 396828 126041 396856 262783
rect 397458 226944 397514 226953
rect 397458 226879 397514 226888
rect 396908 184204 396960 184210
rect 396908 184146 396960 184152
rect 396814 126032 396870 126041
rect 396814 125967 396870 125976
rect 396920 95169 396948 184146
rect 397472 111874 397500 226879
rect 398748 151088 398800 151094
rect 398748 151030 398800 151036
rect 398012 139528 398064 139534
rect 398012 139470 398064 139476
rect 397552 137964 397604 137970
rect 397552 137906 397604 137912
rect 397564 137601 397592 137906
rect 397550 137592 397606 137601
rect 397550 137527 397606 137536
rect 397550 136776 397606 136785
rect 397550 136711 397606 136720
rect 397564 136678 397592 136711
rect 397552 136672 397604 136678
rect 397552 136614 397604 136620
rect 397644 136604 397696 136610
rect 397644 136546 397696 136552
rect 397656 135561 397684 136546
rect 398024 135930 398052 139470
rect 398104 139392 398156 139398
rect 398104 139334 398156 139340
rect 398116 138106 398144 139334
rect 398104 138100 398156 138106
rect 398104 138042 398156 138048
rect 398656 138032 398708 138038
rect 398656 137974 398708 137980
rect 398012 135924 398064 135930
rect 398012 135866 398064 135872
rect 397642 135552 397698 135561
rect 397642 135487 397698 135496
rect 398668 135250 398696 137974
rect 398656 135244 398708 135250
rect 398656 135186 398708 135192
rect 398668 134881 398696 135186
rect 398654 134872 398710 134881
rect 398654 134807 398710 134816
rect 397550 134056 397606 134065
rect 397550 133991 397606 134000
rect 397564 133958 397592 133991
rect 397552 133952 397604 133958
rect 397552 133894 397604 133900
rect 397644 133884 397696 133890
rect 397644 133826 397696 133832
rect 397656 133521 397684 133826
rect 397642 133512 397698 133521
rect 397642 133447 397698 133456
rect 397552 132456 397604 132462
rect 397552 132398 397604 132404
rect 397564 132161 397592 132398
rect 397550 132152 397606 132161
rect 397550 132087 397606 132096
rect 397550 130656 397606 130665
rect 397550 130591 397606 130600
rect 397564 129810 397592 130591
rect 397552 129804 397604 129810
rect 397552 129746 397604 129752
rect 397550 129296 397606 129305
rect 397550 129231 397606 129240
rect 397564 128382 397592 129231
rect 397552 128376 397604 128382
rect 397552 128318 397604 128324
rect 397550 127936 397606 127945
rect 397550 127871 397606 127880
rect 397564 127022 397592 127871
rect 397552 127016 397604 127022
rect 397552 126958 397604 126964
rect 398104 126948 398156 126954
rect 398104 126890 398156 126896
rect 398116 126721 398144 126890
rect 398102 126712 398158 126721
rect 398102 126647 398158 126656
rect 397550 125216 397606 125225
rect 397550 125151 397606 125160
rect 397564 124234 397592 125151
rect 398760 124681 398788 151030
rect 398852 126721 398880 527138
rect 405740 497480 405792 497486
rect 405740 497422 405792 497428
rect 398932 494760 398984 494766
rect 398932 494702 398984 494708
rect 398944 493338 398972 494702
rect 398932 493332 398984 493338
rect 398932 493274 398984 493280
rect 400864 383716 400916 383722
rect 400864 383658 400916 383664
rect 400218 214704 400274 214713
rect 400218 214639 400274 214648
rect 399574 146296 399630 146305
rect 399574 146231 399630 146240
rect 399482 142352 399538 142361
rect 399482 142287 399538 142296
rect 398838 126712 398894 126721
rect 398838 126647 398894 126656
rect 398746 124672 398802 124681
rect 398746 124607 398802 124616
rect 397552 124228 397604 124234
rect 397552 124170 397604 124176
rect 397644 124160 397696 124166
rect 397644 124102 397696 124108
rect 397550 123856 397606 123865
rect 397550 123791 397606 123800
rect 397564 123486 397592 123791
rect 397552 123480 397604 123486
rect 397552 123422 397604 123428
rect 397656 123321 397684 124102
rect 397642 123312 397698 123321
rect 397642 123247 397698 123256
rect 397550 122496 397606 122505
rect 397550 122431 397606 122440
rect 397564 121514 397592 122431
rect 397552 121508 397604 121514
rect 397552 121450 397604 121456
rect 397644 121440 397696 121446
rect 397644 121382 397696 121388
rect 397656 120601 397684 121382
rect 397734 121136 397790 121145
rect 397734 121071 397790 121080
rect 397642 120592 397698 120601
rect 397642 120527 397698 120536
rect 397644 120080 397696 120086
rect 397748 120057 397776 121071
rect 397644 120022 397696 120028
rect 397734 120048 397790 120057
rect 397552 120012 397604 120018
rect 397552 119954 397604 119960
rect 397564 119241 397592 119954
rect 397656 119921 397684 120022
rect 397734 119983 397790 119992
rect 397642 119912 397698 119921
rect 397642 119847 397698 119856
rect 397550 119232 397606 119241
rect 397550 119167 397606 119176
rect 397552 118652 397604 118658
rect 397552 118594 397604 118600
rect 397564 117881 397592 118594
rect 397642 118416 397698 118425
rect 397642 118351 397698 118360
rect 397550 117872 397606 117881
rect 397550 117807 397606 117816
rect 397656 117366 397684 118351
rect 397644 117360 397696 117366
rect 397644 117302 397696 117308
rect 397552 117292 397604 117298
rect 397552 117234 397604 117240
rect 397564 117201 397592 117234
rect 397550 117192 397606 117201
rect 397550 117127 397606 117136
rect 397552 115932 397604 115938
rect 397552 115874 397604 115880
rect 397564 115841 397592 115874
rect 397644 115864 397696 115870
rect 397550 115832 397606 115841
rect 397644 115806 397696 115812
rect 397550 115767 397606 115776
rect 397656 115161 397684 115806
rect 397642 115152 397698 115161
rect 397642 115087 397698 115096
rect 397552 114504 397604 114510
rect 397550 114472 397552 114481
rect 397604 114472 397606 114481
rect 397550 114407 397606 114416
rect 397644 114436 397696 114442
rect 397644 114378 397696 114384
rect 397656 113801 397684 114378
rect 397642 113792 397698 113801
rect 397642 113727 397698 113736
rect 397552 113144 397604 113150
rect 397552 113086 397604 113092
rect 397564 112441 397592 113086
rect 398746 112976 398802 112985
rect 398746 112911 398802 112920
rect 398760 112470 398788 112911
rect 398748 112464 398800 112470
rect 397550 112432 397606 112441
rect 398748 112406 398800 112412
rect 397550 112367 397606 112376
rect 397472 111846 397684 111874
rect 397460 111784 397512 111790
rect 397458 111752 397460 111761
rect 397512 111752 397514 111761
rect 397458 111687 397514 111696
rect 397550 110256 397606 110265
rect 397550 110191 397606 110200
rect 397564 109070 397592 110191
rect 397552 109064 397604 109070
rect 397458 109032 397514 109041
rect 397552 109006 397604 109012
rect 397458 108967 397460 108976
rect 397512 108967 397514 108976
rect 397460 108938 397512 108944
rect 397656 108361 397684 111846
rect 398194 111072 398250 111081
rect 398194 111007 398250 111016
rect 397642 108352 397698 108361
rect 397642 108287 397644 108296
rect 397696 108287 397698 108296
rect 397644 108258 397696 108264
rect 397458 107536 397514 107545
rect 397458 107471 397514 107480
rect 397472 106418 397500 107471
rect 397550 106856 397606 106865
rect 397550 106791 397606 106800
rect 397460 106412 397512 106418
rect 397460 106354 397512 106360
rect 397564 106350 397592 106791
rect 397552 106344 397604 106350
rect 397552 106286 397604 106292
rect 397460 106276 397512 106282
rect 397460 106218 397512 106224
rect 397472 106185 397500 106218
rect 397458 106176 397514 106185
rect 397458 106111 397514 106120
rect 397920 105596 397972 105602
rect 397920 105538 397972 105544
rect 397460 104848 397512 104854
rect 397458 104816 397460 104825
rect 397512 104816 397514 104825
rect 397458 104751 397514 104760
rect 397552 104780 397604 104786
rect 397552 104722 397604 104728
rect 397564 104281 397592 104722
rect 397550 104272 397606 104281
rect 397550 104207 397606 104216
rect 397460 103488 397512 103494
rect 397458 103456 397460 103465
rect 397512 103456 397514 103465
rect 397458 103391 397514 103400
rect 397458 100872 397514 100881
rect 397458 100807 397514 100816
rect 397472 100774 397500 100807
rect 397460 100768 397512 100774
rect 397460 100710 397512 100716
rect 397932 96393 397960 105538
rect 398208 102105 398236 111007
rect 398654 104136 398710 104145
rect 398654 104071 398710 104080
rect 398194 102096 398250 102105
rect 398194 102031 398250 102040
rect 398668 99278 398696 104071
rect 398656 99272 398708 99278
rect 398656 99214 398708 99220
rect 397918 96384 397974 96393
rect 397918 96319 397974 96328
rect 396906 95160 396962 95169
rect 396906 95095 396962 95104
rect 398760 91798 398788 112406
rect 398748 91792 398800 91798
rect 398748 91734 398800 91740
rect 399496 61470 399524 142287
rect 399588 139890 399616 146231
rect 400232 140758 400260 214639
rect 400876 192506 400904 383658
rect 403622 316160 403678 316169
rect 403622 316095 403678 316104
rect 400864 192500 400916 192506
rect 400864 192442 400916 192448
rect 400310 181384 400366 181393
rect 400310 181319 400366 181328
rect 400220 140752 400272 140758
rect 400220 140694 400272 140700
rect 399588 139862 400062 139890
rect 400324 139618 400352 181319
rect 401692 175976 401744 175982
rect 401692 175918 401744 175924
rect 400956 140752 401008 140758
rect 400956 140694 401008 140700
rect 400968 139890 400996 140694
rect 401704 139890 401732 175918
rect 403636 146266 403664 316095
rect 405002 202192 405058 202201
rect 405002 202127 405058 202136
rect 404728 146940 404780 146946
rect 404728 146882 404780 146888
rect 403624 146260 403676 146266
rect 403624 146202 403676 146208
rect 403440 144968 403492 144974
rect 403440 144910 403492 144916
rect 402612 142180 402664 142186
rect 402612 142122 402664 142128
rect 400968 139862 401350 139890
rect 401704 139862 401994 139890
rect 402624 139876 402652 142122
rect 403452 139890 403480 144910
rect 404740 139890 404768 146882
rect 405016 143546 405044 202127
rect 405004 143540 405056 143546
rect 405004 143482 405056 143488
rect 405752 142361 405780 497422
rect 412652 494766 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 700330 429884 703520
rect 462332 702710 462360 703520
rect 478524 702914 478552 703520
rect 478512 702908 478564 702914
rect 478512 702850 478564 702856
rect 494808 702846 494836 703520
rect 494796 702840 494848 702846
rect 494796 702782 494848 702788
rect 462320 702704 462372 702710
rect 462320 702646 462372 702652
rect 527192 702506 527220 703520
rect 543476 702642 543504 703520
rect 543464 702636 543516 702642
rect 543464 702578 543516 702584
rect 559668 702574 559696 703520
rect 559656 702568 559708 702574
rect 559656 702510 559708 702516
rect 527180 702500 527232 702506
rect 527180 702442 527232 702448
rect 429844 700324 429896 700330
rect 429844 700266 429896 700272
rect 582654 697232 582710 697241
rect 582654 697167 582710 697176
rect 582562 683904 582618 683913
rect 582562 683839 582618 683848
rect 582470 644056 582526 644065
rect 582470 643991 582526 644000
rect 582378 564360 582434 564369
rect 582378 564295 582434 564304
rect 582392 557534 582420 564295
rect 582484 558210 582512 643991
rect 582472 558204 582524 558210
rect 582472 558146 582524 558152
rect 582392 557506 582512 557534
rect 582484 556238 582512 557506
rect 582472 556232 582524 556238
rect 582472 556174 582524 556180
rect 580356 554804 580408 554810
rect 580356 554746 580408 554752
rect 580262 538248 580318 538257
rect 580172 538212 580224 538218
rect 580262 538183 580318 538192
rect 580172 538154 580224 538160
rect 580184 537849 580212 538154
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 425060 534812 425112 534818
rect 425060 534754 425112 534760
rect 412640 494760 412692 494766
rect 412640 494702 412692 494708
rect 410524 484424 410576 484430
rect 410524 484366 410576 484372
rect 407854 374640 407910 374649
rect 407854 374575 407910 374584
rect 407120 198008 407172 198014
rect 407120 197950 407172 197956
rect 406014 146976 406070 146985
rect 406014 146911 406070 146920
rect 405738 142352 405794 142361
rect 405738 142287 405794 142296
rect 405752 142154 405780 142287
rect 405752 142126 405872 142154
rect 403452 139862 403926 139890
rect 404740 139862 405214 139890
rect 405844 139876 405872 142126
rect 406028 139890 406056 146911
rect 406028 139862 406502 139890
rect 407132 139876 407160 197950
rect 407868 151814 407896 374575
rect 409878 247616 409934 247625
rect 409878 247551 409934 247560
rect 409892 242962 409920 247551
rect 409880 242956 409932 242962
rect 409880 242898 409932 242904
rect 408590 218648 408646 218657
rect 408590 218583 408646 218592
rect 408604 151814 408632 218583
rect 407868 151786 407988 151814
rect 408604 151786 409368 151814
rect 407304 145580 407356 145586
rect 407304 145522 407356 145528
rect 407316 139890 407344 145522
rect 407960 140049 407988 151786
rect 409052 143540 409104 143546
rect 409052 143482 409104 143488
rect 407946 140040 408002 140049
rect 407946 139975 408002 139984
rect 407316 139862 407790 139890
rect 409064 139876 409092 143482
rect 409340 139890 409368 151786
rect 409892 139890 409920 242898
rect 409972 159384 410024 159390
rect 410536 159361 410564 484366
rect 416780 401668 416832 401674
rect 416780 401610 416832 401616
rect 412546 376816 412602 376825
rect 412546 376751 412602 376760
rect 411258 203688 411314 203697
rect 411258 203623 411314 203632
rect 409972 159326 410024 159332
rect 410522 159352 410578 159361
rect 409984 151814 410012 159326
rect 410522 159287 410578 159296
rect 409984 151786 410656 151814
rect 410628 139890 410656 151786
rect 411272 139890 411300 203623
rect 412560 146266 412588 376751
rect 412640 366376 412692 366382
rect 412640 366318 412692 366324
rect 411904 146260 411956 146266
rect 411904 146202 411956 146208
rect 412548 146260 412600 146266
rect 412548 146202 412600 146208
rect 411916 139890 411944 146202
rect 412652 142769 412680 366318
rect 414664 294636 414716 294642
rect 414664 294578 414716 294584
rect 414676 146946 414704 294578
rect 415400 192500 415452 192506
rect 415400 192442 415452 192448
rect 414664 146940 414716 146946
rect 414664 146882 414716 146888
rect 414480 146260 414532 146266
rect 414480 146202 414532 146208
rect 412638 142760 412694 142769
rect 412638 142695 412694 142704
rect 414204 142248 414256 142254
rect 414204 142190 414256 142196
rect 409340 139862 409722 139890
rect 409892 139862 410366 139890
rect 410628 139862 411010 139890
rect 411272 139862 411654 139890
rect 411916 139862 412298 139890
rect 414216 139876 414244 142190
rect 414492 139890 414520 146202
rect 415412 143449 415440 192442
rect 415398 143440 415454 143449
rect 415398 143375 415454 143384
rect 416134 143440 416190 143449
rect 416134 143375 416190 143384
rect 415490 142760 415546 142769
rect 415490 142695 415546 142704
rect 414492 139862 414874 139890
rect 415504 139876 415532 142695
rect 416148 142225 416176 143375
rect 416134 142216 416190 142225
rect 416134 142151 416190 142160
rect 416148 139876 416176 142151
rect 416792 141438 416820 401610
rect 418804 360868 418856 360874
rect 418804 360810 418856 360816
rect 417424 171828 417476 171834
rect 417424 171770 417476 171776
rect 417436 144906 417464 171770
rect 417424 144900 417476 144906
rect 417424 144842 417476 144848
rect 418068 144900 418120 144906
rect 418068 144842 418120 144848
rect 416780 141432 416832 141438
rect 416780 141374 416832 141380
rect 416792 139876 416820 141374
rect 418080 139876 418108 144842
rect 399852 139596 399904 139602
rect 400324 139596 400706 139618
rect 400324 139590 400404 139596
rect 399852 139538 399904 139544
rect 400456 139590 400706 139596
rect 400404 139538 400456 139544
rect 399864 137737 399892 139538
rect 404360 139528 404412 139534
rect 418816 139482 418844 360810
rect 420920 344344 420972 344350
rect 420920 344286 420972 344292
rect 420182 214568 420238 214577
rect 420182 214503 420238 214512
rect 418894 204912 418950 204921
rect 418894 204847 418950 204856
rect 418908 143546 418936 204847
rect 419632 173188 419684 173194
rect 419632 173130 419684 173136
rect 419644 151814 419672 173130
rect 420196 151814 420224 214503
rect 419644 151786 420132 151814
rect 420196 151786 420316 151814
rect 418896 143540 418948 143546
rect 418896 143482 418948 143488
rect 420000 143540 420052 143546
rect 420000 143482 420052 143488
rect 420012 139876 420040 143482
rect 420104 142154 420132 151786
rect 420104 142126 420224 142154
rect 420196 139890 420224 142126
rect 420288 140078 420316 151786
rect 420276 140072 420328 140078
rect 420276 140014 420328 140020
rect 420932 139890 420960 344286
rect 423678 208448 423734 208457
rect 423678 208383 423734 208392
rect 422942 206272 422998 206281
rect 422942 206207 422998 206216
rect 422300 156664 422352 156670
rect 422300 156606 422352 156612
rect 422312 151814 422340 156606
rect 422312 151786 422800 151814
rect 421472 145580 421524 145586
rect 421472 145522 421524 145528
rect 421484 139890 421512 145522
rect 422576 140888 422628 140894
rect 422576 140830 422628 140836
rect 420196 139862 420670 139890
rect 420932 139862 421314 139890
rect 421484 139862 421958 139890
rect 422588 139876 422616 140830
rect 422772 139890 422800 151786
rect 422956 142866 422984 206207
rect 423036 153876 423088 153882
rect 423036 153818 423088 153824
rect 422944 142860 422996 142866
rect 422944 142802 422996 142808
rect 423048 140894 423076 153818
rect 423036 140888 423088 140894
rect 423036 140830 423088 140836
rect 423692 140826 423720 208383
rect 425072 143449 425100 534754
rect 445760 518968 445812 518974
rect 445760 518910 445812 518916
rect 434720 505164 434772 505170
rect 434720 505106 434772 505112
rect 427818 317520 427874 317529
rect 427818 317455 427874 317464
rect 426438 203552 426494 203561
rect 426438 203487 426494 203496
rect 425150 149152 425206 149161
rect 425150 149087 425206 149096
rect 425058 143440 425114 143449
rect 425058 143375 425114 143384
rect 423680 140820 423732 140826
rect 423680 140762 423732 140768
rect 424508 140820 424560 140826
rect 424508 140762 424560 140768
rect 422772 139862 423246 139890
rect 424520 139876 424548 140762
rect 425164 139876 425192 149087
rect 425794 143440 425850 143449
rect 425794 143375 425850 143384
rect 419630 139496 419686 139505
rect 404412 139476 404570 139482
rect 404360 139470 404570 139476
rect 404372 139454 404570 139470
rect 417160 139466 417450 139482
rect 417148 139460 417450 139466
rect 417200 139454 417450 139460
rect 418816 139454 419630 139482
rect 419630 139431 419686 139440
rect 425518 139496 425574 139505
rect 425808 139482 425836 143375
rect 425574 139468 425836 139482
rect 426452 139482 426480 203487
rect 427832 151814 427860 317455
rect 432602 314800 432658 314809
rect 432602 314735 432658 314744
rect 428464 284368 428516 284374
rect 428464 284310 428516 284316
rect 427832 151786 427952 151814
rect 427082 142216 427138 142225
rect 427082 142151 427138 142160
rect 427096 139876 427124 142151
rect 427924 139890 427952 151786
rect 428476 142186 428504 284310
rect 429844 249076 429896 249082
rect 429844 249018 429896 249024
rect 429198 197976 429254 197985
rect 429198 197911 429254 197920
rect 428464 142180 428516 142186
rect 428464 142122 428516 142128
rect 429212 139890 429240 197911
rect 429856 148442 429884 249018
rect 431868 214600 431920 214606
rect 431868 214542 431920 214548
rect 431224 200796 431276 200802
rect 431224 200738 431276 200744
rect 430580 158024 430632 158030
rect 430580 157966 430632 157972
rect 429936 151156 429988 151162
rect 429936 151098 429988 151104
rect 429844 148436 429896 148442
rect 429844 148378 429896 148384
rect 429948 139890 429976 151098
rect 430592 139890 430620 157966
rect 431236 141438 431264 200738
rect 431224 141432 431276 141438
rect 431224 141374 431276 141380
rect 427924 139862 428398 139890
rect 429212 139862 429686 139890
rect 429948 139862 430330 139890
rect 430592 139862 430974 139890
rect 427450 139496 427506 139505
rect 426452 139468 426848 139482
rect 425574 139454 425822 139468
rect 426466 139466 426848 139468
rect 426466 139460 426860 139466
rect 426466 139454 426808 139460
rect 425518 139431 425574 139440
rect 417148 139402 417200 139408
rect 431314 139496 431370 139505
rect 427506 139454 427754 139482
rect 427450 139431 427506 139440
rect 431880 139482 431908 214542
rect 432236 142860 432288 142866
rect 432236 142802 432288 142808
rect 432248 139876 432276 142802
rect 432616 140865 432644 314735
rect 434732 214606 434760 505106
rect 443000 299532 443052 299538
rect 443000 299474 443052 299480
rect 439412 295384 439464 295390
rect 439412 295326 439464 295332
rect 436744 273964 436796 273970
rect 436744 273906 436796 273912
rect 434812 234660 434864 234666
rect 434812 234602 434864 234608
rect 434720 214600 434772 214606
rect 434720 214542 434772 214548
rect 432696 193248 432748 193254
rect 432696 193190 432748 193196
rect 432708 147014 432736 193190
rect 434720 167680 434772 167686
rect 434720 167622 434772 167628
rect 432696 147008 432748 147014
rect 432696 146950 432748 146956
rect 433522 143576 433578 143585
rect 433522 143511 433578 143520
rect 432880 142180 432932 142186
rect 432880 142122 432932 142128
rect 432602 140856 432658 140865
rect 432602 140791 432658 140800
rect 432892 139876 432920 142122
rect 433536 139876 433564 143511
rect 434732 140758 434760 167622
rect 434720 140752 434772 140758
rect 434720 140694 434772 140700
rect 434824 139876 434852 234602
rect 436100 225004 436152 225010
rect 436100 224946 436152 224952
rect 436112 140758 436140 224946
rect 436756 151162 436784 273906
rect 439134 211848 439190 211857
rect 439134 211783 439190 211792
rect 438124 209092 438176 209098
rect 438124 209034 438176 209040
rect 436836 155236 436888 155242
rect 436836 155178 436888 155184
rect 436744 151156 436796 151162
rect 436744 151098 436796 151104
rect 436376 146940 436428 146946
rect 436376 146882 436428 146888
rect 435180 140752 435232 140758
rect 435180 140694 435232 140700
rect 436100 140752 436152 140758
rect 436100 140694 436152 140700
rect 435192 139890 435220 140694
rect 436388 139890 436416 146882
rect 436848 143546 436876 155178
rect 438136 151814 438164 209034
rect 438136 151786 438256 151814
rect 437664 148368 437716 148374
rect 437664 148310 437716 148316
rect 436836 143540 436888 143546
rect 436836 143482 436888 143488
rect 437020 140752 437072 140758
rect 437020 140694 437072 140700
rect 437032 139890 437060 140694
rect 437676 139890 437704 148310
rect 435192 139862 435482 139890
rect 436388 139862 436770 139890
rect 437032 139862 437414 139890
rect 437676 139862 438058 139890
rect 436374 139496 436430 139505
rect 431370 139454 431908 139482
rect 436126 139454 436374 139482
rect 431314 139431 431370 139440
rect 436374 139431 436430 139440
rect 426808 139402 426860 139408
rect 438228 139398 438256 151786
rect 412732 139392 412784 139398
rect 438216 139392 438268 139398
rect 412784 139340 412942 139346
rect 412732 139334 412942 139340
rect 438858 139360 438914 139369
rect 438216 139334 438268 139340
rect 412744 139318 412942 139334
rect 438702 139318 438858 139346
rect 438858 139295 438914 139304
rect 399850 137728 399906 137737
rect 399850 137663 399906 137672
rect 439148 132494 439176 211783
rect 439320 143540 439372 143546
rect 439320 143482 439372 143488
rect 439332 139876 439360 143482
rect 439148 132466 439360 132494
rect 439332 111897 439360 132466
rect 439424 131753 439452 295326
rect 441620 257372 441672 257378
rect 441620 257314 441672 257320
rect 440238 207088 440294 207097
rect 440238 207023 440294 207032
rect 440252 206990 440280 207023
rect 440240 206984 440292 206990
rect 440240 206926 440292 206932
rect 440884 206984 440936 206990
rect 440884 206926 440936 206932
rect 439596 149728 439648 149734
rect 439596 149670 439648 149676
rect 439504 139392 439556 139398
rect 439504 139334 439556 139340
rect 439516 135833 439544 139334
rect 439608 138553 439636 149670
rect 440424 148436 440476 148442
rect 440424 148378 440476 148384
rect 440332 141432 440384 141438
rect 440332 141374 440384 141380
rect 440240 140072 440292 140078
rect 440240 140014 440292 140020
rect 439594 138544 439650 138553
rect 439594 138479 439650 138488
rect 439502 135824 439558 135833
rect 439502 135759 439558 135768
rect 440252 132841 440280 140014
rect 440238 132832 440294 132841
rect 440238 132767 440294 132776
rect 439410 131744 439466 131753
rect 439410 131679 439466 131688
rect 440238 127936 440294 127945
rect 440238 127871 440294 127880
rect 439410 120864 439466 120873
rect 439410 120799 439466 120808
rect 439424 115977 439452 120799
rect 439410 115968 439466 115977
rect 439410 115903 439466 115912
rect 439318 111888 439374 111897
rect 439318 111823 439374 111832
rect 439318 104408 439374 104417
rect 439318 104343 439374 104352
rect 439332 103514 439360 104343
rect 439410 103864 439466 103873
rect 439410 103799 439466 103808
rect 439148 103486 439360 103514
rect 400048 97889 400076 100028
rect 400034 97880 400090 97889
rect 400034 97815 400090 97824
rect 399484 61464 399536 61470
rect 399484 61406 399536 61412
rect 400692 46918 400720 100028
rect 400862 96928 400918 96937
rect 400862 96863 400918 96872
rect 400680 46912 400732 46918
rect 400680 46854 400732 46860
rect 400876 44878 400904 96863
rect 401336 95266 401364 100028
rect 401324 95260 401376 95266
rect 401324 95202 401376 95208
rect 401980 67590 402008 100028
rect 402624 96937 402652 100028
rect 403268 99278 403296 100028
rect 403256 99272 403308 99278
rect 403256 99214 403308 99220
rect 403912 97918 403940 100028
rect 404556 99385 404584 100028
rect 405844 99414 405872 100028
rect 405832 99408 405884 99414
rect 404542 99376 404598 99385
rect 405832 99350 405884 99356
rect 404542 99311 404598 99320
rect 403900 97912 403952 97918
rect 403900 97854 403952 97860
rect 402610 96928 402666 96937
rect 402610 96863 402666 96872
rect 402980 95260 403032 95266
rect 402980 95202 403032 95208
rect 401968 67584 402020 67590
rect 401968 67526 402020 67532
rect 400864 44872 400916 44878
rect 400864 44814 400916 44820
rect 396724 5500 396776 5506
rect 396724 5442 396776 5448
rect 402992 4078 403020 95202
rect 404556 84194 404584 99311
rect 405844 99278 405872 99350
rect 405832 99272 405884 99278
rect 405832 99214 405884 99220
rect 406488 96393 406516 100028
rect 405738 96384 405794 96393
rect 405738 96319 405794 96328
rect 406474 96384 406530 96393
rect 406474 96319 406530 96328
rect 404372 84166 404584 84194
rect 404372 82142 404400 84166
rect 404360 82136 404412 82142
rect 404360 82078 404412 82084
rect 405752 43450 405780 96319
rect 407132 59362 407160 100028
rect 407120 59356 407172 59362
rect 407120 59298 407172 59304
rect 405740 43444 405792 43450
rect 405740 43386 405792 43392
rect 407776 15910 407804 100028
rect 408420 99482 408448 100028
rect 408408 99476 408460 99482
rect 408408 99418 408460 99424
rect 409064 96898 409092 100028
rect 409052 96892 409104 96898
rect 409052 96834 409104 96840
rect 409708 93809 409736 100028
rect 409972 96892 410024 96898
rect 409972 96834 410024 96840
rect 409694 93800 409750 93809
rect 409694 93735 409750 93744
rect 409708 92585 409736 93735
rect 408498 92576 408554 92585
rect 408498 92511 408554 92520
rect 409694 92576 409750 92585
rect 409694 92511 409750 92520
rect 408512 50386 408540 92511
rect 408500 50380 408552 50386
rect 408500 50322 408552 50328
rect 409984 18630 410012 96834
rect 410996 89729 411024 100028
rect 410982 89720 411038 89729
rect 410982 89655 411038 89664
rect 409972 18624 410024 18630
rect 409972 18566 410024 18572
rect 407764 15904 407816 15910
rect 407764 15846 407816 15852
rect 411640 6866 411668 100028
rect 412284 95130 412312 100028
rect 412928 96422 412956 100028
rect 413572 99929 413600 100028
rect 413558 99920 413614 99929
rect 413558 99855 413614 99864
rect 413284 96960 413336 96966
rect 413284 96902 413336 96908
rect 412916 96416 412968 96422
rect 412916 96358 412968 96364
rect 412272 95124 412324 95130
rect 412272 95066 412324 95072
rect 412284 93129 412312 95066
rect 412270 93120 412326 93129
rect 412270 93055 412326 93064
rect 413296 17270 413324 96902
rect 413376 96416 413428 96422
rect 413376 96358 413428 96364
rect 413388 95266 413416 96358
rect 413376 95260 413428 95266
rect 413376 95202 413428 95208
rect 413388 85542 413416 95202
rect 413376 85536 413428 85542
rect 413376 85478 413428 85484
rect 414216 72486 414244 100028
rect 414860 99929 414888 100028
rect 414846 99920 414902 99929
rect 414846 99855 414902 99864
rect 414662 97200 414718 97209
rect 414662 97135 414718 97144
rect 414204 72480 414256 72486
rect 414204 72422 414256 72428
rect 413284 17264 413336 17270
rect 413284 17206 413336 17212
rect 414676 13122 414704 97135
rect 416148 96966 416176 100028
rect 416136 96960 416188 96966
rect 416136 96902 416188 96908
rect 416792 51814 416820 100028
rect 416780 51808 416832 51814
rect 416780 51750 416832 51756
rect 417436 27606 417464 100028
rect 418080 91769 418108 100028
rect 418724 96529 418752 100028
rect 418710 96520 418766 96529
rect 418710 96455 418766 96464
rect 418066 91760 418122 91769
rect 418066 91695 418122 91704
rect 417424 27600 417476 27606
rect 417424 27542 417476 27548
rect 419368 24206 419396 100028
rect 420012 99113 420040 100028
rect 419998 99104 420054 99113
rect 419998 99039 420054 99048
rect 420012 96626 420040 99039
rect 420000 96620 420052 96626
rect 420000 96562 420052 96568
rect 421300 93906 421328 100028
rect 421944 99249 421972 100028
rect 421930 99240 421986 99249
rect 421930 99175 421986 99184
rect 421288 93900 421340 93906
rect 421288 93842 421340 93848
rect 421300 91089 421328 93842
rect 421286 91080 421342 91089
rect 421286 91015 421342 91024
rect 422588 54602 422616 100028
rect 423232 96898 423260 100028
rect 423876 97209 423904 100028
rect 423862 97200 423918 97209
rect 423862 97135 423918 97144
rect 423220 96892 423272 96898
rect 423220 96834 423272 96840
rect 424520 93770 424548 100028
rect 424508 93764 424560 93770
rect 424508 93706 424560 93712
rect 425164 88262 425192 100028
rect 425702 97064 425758 97073
rect 425702 96999 425758 97008
rect 425152 88256 425204 88262
rect 425152 88198 425204 88204
rect 425716 63510 425744 96999
rect 426452 93838 426480 100028
rect 427096 96937 427124 100028
rect 427740 97073 427768 100028
rect 427726 97064 427782 97073
rect 427726 96999 427782 97008
rect 427082 96928 427138 96937
rect 427082 96863 427138 96872
rect 427910 96928 427966 96937
rect 427910 96863 427966 96872
rect 426440 93832 426492 93838
rect 426440 93774 426492 93780
rect 425704 63504 425756 63510
rect 425704 63446 425756 63452
rect 422576 54596 422628 54602
rect 422576 54538 422628 54544
rect 419356 24200 419408 24206
rect 419356 24142 419408 24148
rect 414664 13116 414716 13122
rect 414664 13058 414716 13064
rect 411628 6860 411680 6866
rect 411628 6802 411680 6808
rect 427924 6186 427952 96863
rect 428384 65550 428412 100028
rect 429028 99346 429056 100028
rect 429016 99340 429068 99346
rect 429016 99282 429068 99288
rect 429292 96892 429344 96898
rect 429292 96834 429344 96840
rect 428372 65544 428424 65550
rect 428372 65486 428424 65492
rect 429304 20670 429332 96834
rect 429672 95198 429700 100028
rect 429660 95192 429712 95198
rect 429660 95134 429712 95140
rect 430316 89690 430344 100028
rect 431604 97753 431632 100028
rect 431590 97744 431646 97753
rect 431590 97679 431646 97688
rect 432248 92478 432276 100028
rect 432892 97986 432920 100028
rect 433536 99929 433564 100028
rect 433522 99920 433578 99929
rect 433522 99855 433578 99864
rect 434180 99210 434208 100028
rect 434824 99929 434852 100028
rect 434810 99920 434866 99929
rect 434810 99855 434866 99864
rect 434168 99204 434220 99210
rect 434168 99146 434220 99152
rect 432880 97980 432932 97986
rect 432880 97922 432932 97928
rect 434824 97889 434852 99855
rect 434810 97880 434866 97889
rect 434810 97815 434866 97824
rect 432696 97232 432748 97238
rect 432696 97174 432748 97180
rect 432604 95872 432656 95878
rect 432604 95814 432656 95820
rect 432236 92472 432288 92478
rect 432236 92414 432288 92420
rect 430304 89684 430356 89690
rect 430304 89626 430356 89632
rect 432616 82822 432644 95814
rect 432708 86970 432736 97174
rect 432696 86964 432748 86970
rect 432696 86906 432748 86912
rect 432604 82816 432656 82822
rect 432604 82758 432656 82764
rect 435468 53786 435496 100028
rect 436756 96914 436784 100028
rect 436836 99340 436888 99346
rect 436836 99282 436888 99288
rect 436112 96886 436784 96914
rect 435456 53780 435508 53786
rect 435456 53722 435508 53728
rect 436112 39370 436140 96886
rect 436848 84194 436876 99282
rect 437400 97889 437428 100028
rect 438044 97986 438072 100028
rect 438032 97980 438084 97986
rect 438032 97922 438084 97928
rect 437386 97880 437442 97889
rect 437386 97815 437442 97824
rect 438688 95169 438716 100028
rect 439148 95878 439176 103486
rect 439318 101688 439374 101697
rect 439318 101623 439374 101632
rect 439332 101590 439360 101623
rect 439320 101584 439372 101590
rect 439320 101526 439372 101532
rect 439136 95872 439188 95878
rect 439136 95814 439188 95820
rect 438674 95160 438730 95169
rect 438674 95095 438730 95104
rect 439332 84194 439360 100028
rect 436756 84166 436876 84194
rect 439240 84166 439360 84194
rect 436756 80034 436784 84166
rect 436744 80028 436796 80034
rect 436744 79970 436796 79976
rect 439240 75886 439268 84166
rect 439228 75880 439280 75886
rect 439228 75822 439280 75828
rect 436100 39364 436152 39370
rect 436100 39306 436152 39312
rect 429292 20664 429344 20670
rect 429292 20606 429344 20612
rect 439424 9654 439452 103799
rect 439502 102368 439558 102377
rect 439502 102303 439558 102312
rect 439516 99346 439544 102303
rect 439504 99340 439556 99346
rect 439504 99282 439556 99288
rect 440252 69698 440280 127871
rect 440344 121961 440372 141374
rect 440436 137465 440464 148378
rect 440422 137456 440478 137465
rect 440422 137391 440478 137400
rect 440436 136678 440464 137391
rect 440424 136672 440476 136678
rect 440424 136614 440476 136620
rect 440330 121952 440386 121961
rect 440330 121887 440386 121896
rect 440422 119096 440478 119105
rect 440422 119031 440478 119040
rect 440330 115016 440386 115025
rect 440330 114951 440386 114960
rect 440344 83502 440372 114951
rect 440436 97238 440464 119031
rect 440896 114481 440924 206926
rect 441632 124001 441660 257314
rect 441710 180024 441766 180033
rect 441710 179959 441766 179968
rect 441724 147098 441752 179959
rect 441804 152516 441856 152522
rect 441804 152458 441856 152464
rect 441816 151814 441844 152458
rect 441816 151786 442028 151814
rect 441724 147070 441936 147098
rect 441804 146872 441856 146878
rect 441804 146814 441856 146820
rect 441712 144220 441764 144226
rect 441712 144162 441764 144168
rect 441724 136241 441752 144162
rect 441710 136232 441766 136241
rect 441710 136167 441766 136176
rect 441816 132161 441844 146814
rect 441908 138961 441936 147070
rect 442000 146878 442028 151786
rect 441988 146872 442040 146878
rect 441988 146814 442040 146820
rect 441894 138952 441950 138961
rect 441894 138887 441950 138896
rect 441986 138136 442042 138145
rect 441986 138071 442042 138080
rect 442000 136610 442028 138071
rect 442906 136776 442962 136785
rect 442906 136711 442908 136720
rect 442960 136711 442962 136720
rect 442908 136682 442960 136688
rect 441988 136604 442040 136610
rect 441988 136546 442040 136552
rect 442906 134872 442962 134881
rect 442906 134807 442962 134816
rect 442920 134570 442948 134807
rect 442908 134564 442960 134570
rect 442908 134506 442960 134512
rect 442908 133884 442960 133890
rect 442908 133826 442960 133832
rect 442920 133521 442948 133826
rect 442906 133512 442962 133521
rect 442906 133447 442962 133456
rect 441802 132152 441858 132161
rect 441802 132087 441858 132096
rect 442908 130824 442960 130830
rect 442906 130792 442908 130801
rect 442960 130792 442962 130801
rect 442906 130727 442962 130736
rect 442906 129976 442962 129985
rect 442906 129911 442962 129920
rect 442920 129810 442948 129911
rect 442908 129804 442960 129810
rect 442908 129746 442960 129752
rect 442170 129296 442226 129305
rect 442170 129231 442226 129240
rect 442184 128382 442212 129231
rect 442172 128376 442224 128382
rect 442172 128318 442224 128324
rect 442906 127256 442962 127265
rect 442906 127191 442908 127200
rect 442960 127191 442962 127200
rect 442908 127162 442960 127168
rect 442908 126948 442960 126954
rect 442908 126890 442960 126896
rect 442816 126880 442868 126886
rect 442816 126822 442868 126828
rect 442828 126041 442856 126822
rect 442920 126721 442948 126890
rect 442906 126712 442962 126721
rect 442906 126647 442962 126656
rect 442814 126032 442870 126041
rect 442814 125967 442870 125976
rect 442908 125588 442960 125594
rect 442908 125530 442960 125536
rect 442920 124681 442948 125530
rect 442906 124672 442962 124681
rect 442906 124607 442962 124616
rect 442632 124160 442684 124166
rect 442632 124102 442684 124108
rect 442644 124001 442672 124102
rect 441618 123992 441674 124001
rect 441618 123927 441674 123936
rect 442630 123992 442686 124001
rect 442630 123927 442686 123936
rect 441896 122664 441948 122670
rect 441894 122632 441896 122641
rect 441948 122632 441950 122641
rect 441894 122567 441950 122576
rect 441618 120456 441674 120465
rect 441618 120391 441674 120400
rect 440882 114472 440938 114481
rect 440882 114407 440938 114416
rect 440424 97232 440476 97238
rect 440424 97174 440476 97180
rect 441632 84833 441660 120391
rect 442908 118584 442960 118590
rect 442906 118552 442908 118561
rect 442960 118552 442962 118561
rect 442906 118487 442962 118496
rect 442906 117192 442962 117201
rect 443012 117178 443040 299474
rect 444378 220144 444434 220153
rect 444378 220079 444434 220088
rect 443090 188320 443146 188329
rect 443090 188255 443146 188264
rect 443104 134570 443132 188255
rect 443182 148336 443238 148345
rect 443182 148271 443238 148280
rect 443092 134564 443144 134570
rect 443092 134506 443144 134512
rect 443090 125216 443146 125225
rect 443090 125151 443146 125160
rect 442962 117150 443040 117178
rect 442906 117127 442962 117136
rect 442906 116376 442962 116385
rect 442906 116311 442908 116320
rect 442960 116311 442962 116320
rect 442908 116282 442960 116288
rect 442908 115864 442960 115870
rect 442906 115832 442908 115841
rect 442960 115832 442962 115841
rect 442906 115767 442962 115776
rect 442906 113656 442962 113665
rect 442906 113591 442962 113600
rect 442920 113422 442948 113591
rect 442908 113416 442960 113422
rect 442908 113358 442960 113364
rect 442908 113144 442960 113150
rect 442906 113112 442908 113121
rect 442960 113112 442962 113121
rect 442906 113047 442962 113056
rect 442170 109576 442226 109585
rect 442170 109511 442226 109520
rect 442184 109070 442212 109511
rect 442172 109064 442224 109070
rect 442172 109006 442224 109012
rect 442446 109032 442502 109041
rect 442446 108967 442448 108976
rect 442500 108967 442502 108976
rect 442448 108938 442500 108944
rect 441710 108216 441766 108225
rect 441710 108151 441766 108160
rect 441618 84824 441674 84833
rect 441618 84759 441674 84768
rect 440332 83496 440384 83502
rect 440332 83438 440384 83444
rect 441724 73846 441752 108151
rect 442906 107536 442962 107545
rect 442962 107494 443040 107522
rect 442906 107471 442962 107480
rect 442724 106276 442776 106282
rect 442724 106218 442776 106224
rect 442354 106176 442410 106185
rect 442354 106111 442410 106120
rect 442368 104922 442396 106111
rect 442736 105641 442764 106218
rect 442722 105632 442778 105641
rect 442722 105567 442778 105576
rect 442356 104916 442408 104922
rect 442356 104858 442408 104864
rect 442172 101652 442224 101658
rect 442172 101594 442224 101600
rect 442184 100881 442212 101594
rect 442170 100872 442226 100881
rect 442170 100807 442226 100816
rect 442908 100700 442960 100706
rect 442908 100642 442960 100648
rect 442920 100201 442948 100642
rect 442906 100192 442962 100201
rect 442906 100127 442962 100136
rect 441712 73840 441764 73846
rect 441712 73782 441764 73788
rect 440240 69692 440292 69698
rect 440240 69634 440292 69640
rect 443012 35902 443040 107494
rect 443104 71777 443132 125151
rect 443196 103465 443224 148271
rect 443276 147008 443328 147014
rect 443276 146950 443328 146956
rect 443288 109002 443316 146950
rect 444392 130830 444420 220079
rect 444564 163532 444616 163538
rect 444564 163474 444616 163480
rect 444380 130824 444432 130830
rect 444380 130766 444432 130772
rect 444472 128376 444524 128382
rect 444472 128318 444524 128324
rect 444380 113416 444432 113422
rect 444380 113358 444432 113364
rect 443368 109064 443420 109070
rect 443368 109006 443420 109012
rect 443276 108996 443328 109002
rect 443276 108938 443328 108944
rect 443182 103456 443238 103465
rect 443182 103391 443238 103400
rect 443380 88330 443408 109006
rect 443368 88324 443420 88330
rect 443368 88266 443420 88272
rect 443090 71768 443146 71777
rect 443090 71703 443146 71712
rect 444392 49026 444420 113358
rect 444484 86290 444512 128318
rect 444576 122670 444604 163474
rect 444564 122664 444616 122670
rect 444564 122606 444616 122612
rect 445772 99346 445800 518910
rect 580276 484673 580304 538183
rect 580368 524521 580396 554746
rect 580354 524512 580410 524521
rect 580354 524447 580410 524456
rect 582380 520328 582432 520334
rect 582380 520270 582432 520276
rect 582392 511329 582420 520270
rect 582378 511320 582434 511329
rect 582378 511255 582434 511264
rect 580262 484664 580318 484673
rect 580262 484599 580318 484608
rect 582380 455456 582432 455462
rect 582380 455398 582432 455404
rect 582392 431633 582420 455398
rect 582378 431624 582434 431633
rect 582378 431559 582434 431568
rect 582378 365120 582434 365129
rect 582378 365055 582434 365064
rect 582392 336025 582420 365055
rect 582378 336016 582434 336025
rect 582378 335951 582434 335960
rect 582378 333296 582434 333305
rect 582378 333231 582434 333240
rect 447140 288448 447192 288454
rect 447140 288390 447192 288396
rect 445942 182880 445998 182889
rect 445942 182815 445998 182824
rect 445850 177304 445906 177313
rect 445850 177239 445906 177248
rect 445864 118590 445892 177239
rect 445852 118584 445904 118590
rect 445852 118526 445904 118532
rect 445852 104916 445904 104922
rect 445852 104858 445904 104864
rect 445760 99340 445812 99346
rect 445760 99282 445812 99288
rect 444472 86284 444524 86290
rect 444472 86226 444524 86232
rect 444380 49020 444432 49026
rect 444380 48962 444432 48968
rect 443000 35896 443052 35902
rect 443000 35838 443052 35844
rect 439412 9648 439464 9654
rect 439412 9590 439464 9596
rect 427912 6180 427964 6186
rect 427912 6122 427964 6128
rect 402980 4072 403032 4078
rect 382922 4040 382978 4049
rect 402980 4014 403032 4020
rect 382922 3975 382978 3984
rect 360844 3460 360896 3466
rect 360844 3402 360896 3408
rect 358082 3360 358138 3369
rect 358082 3295 358138 3304
rect 445864 2786 445892 104858
rect 445956 101658 445984 182815
rect 446034 109848 446090 109857
rect 446034 109783 446090 109792
rect 445944 101652 445996 101658
rect 445944 101594 445996 101600
rect 446048 57254 446076 109783
rect 447152 97986 447180 288390
rect 449900 279472 449952 279478
rect 449900 279414 449952 279420
rect 449162 246256 449218 246265
rect 449162 246191 449218 246200
rect 447324 191140 447376 191146
rect 447324 191082 447376 191088
rect 447230 119368 447286 119377
rect 447230 119303 447286 119312
rect 447140 97980 447192 97986
rect 447140 97922 447192 97928
rect 446036 57248 446088 57254
rect 446036 57190 446088 57196
rect 447244 21418 447272 119303
rect 447336 115870 447364 191082
rect 448612 151156 448664 151162
rect 448612 151098 448664 151104
rect 448520 127220 448572 127226
rect 448520 127162 448572 127168
rect 447324 115864 447376 115870
rect 447324 115806 447376 115812
rect 447232 21412 447284 21418
rect 447232 21354 447284 21360
rect 448532 12442 448560 127162
rect 448624 97889 448652 151098
rect 449176 102134 449204 246191
rect 449912 149054 449940 279414
rect 460940 251864 460992 251870
rect 460940 251806 460992 251812
rect 452660 240780 452712 240786
rect 452660 240722 452712 240728
rect 449990 189680 450046 189689
rect 449990 189615 450046 189624
rect 449900 149048 449952 149054
rect 449900 148990 449952 148996
rect 449912 148374 449940 148990
rect 449900 148368 449952 148374
rect 449900 148310 449952 148316
rect 449900 116340 449952 116346
rect 449900 116282 449952 116288
rect 449164 102128 449216 102134
rect 449164 102070 449216 102076
rect 449176 100706 449204 102070
rect 449164 100700 449216 100706
rect 449164 100642 449216 100648
rect 448610 97880 448666 97889
rect 448610 97815 448666 97824
rect 448520 12436 448572 12442
rect 448520 12378 448572 12384
rect 449912 10334 449940 116282
rect 450004 109857 450032 189615
rect 449990 109848 450046 109857
rect 449990 109783 450046 109792
rect 452672 106282 452700 240722
rect 454040 221468 454092 221474
rect 454040 221410 454092 221416
rect 452752 136740 452804 136746
rect 452752 136682 452804 136688
rect 452660 106276 452712 106282
rect 452660 106218 452712 106224
rect 452764 42770 452792 136682
rect 454052 126886 454080 221410
rect 456800 215960 456852 215966
rect 456800 215902 456852 215908
rect 454132 129804 454184 129810
rect 454132 129746 454184 129752
rect 454040 126880 454092 126886
rect 454040 126822 454092 126828
rect 454144 47598 454172 129746
rect 456812 113150 456840 215902
rect 456892 134564 456944 134570
rect 456892 134506 456944 134512
rect 456800 113144 456852 113150
rect 456800 113086 456852 113092
rect 454132 47592 454184 47598
rect 454132 47534 454184 47540
rect 452752 42764 452804 42770
rect 452752 42706 452804 42712
rect 456904 37942 456932 134506
rect 460952 125594 460980 251806
rect 580906 165880 580962 165889
rect 580906 165815 580962 165824
rect 580920 147014 580948 165815
rect 580908 147008 580960 147014
rect 580908 146950 580960 146956
rect 580264 140820 580316 140826
rect 580264 140762 580316 140768
rect 580170 139360 580226 139369
rect 580170 139295 580226 139304
rect 580184 138038 580212 139295
rect 580172 138032 580224 138038
rect 580172 137974 580224 137980
rect 580276 126041 580304 140762
rect 580262 126032 580318 126041
rect 580262 125967 580318 125976
rect 460940 125588 460992 125594
rect 460940 125530 460992 125536
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580184 99414 580212 99447
rect 580172 99408 580224 99414
rect 580172 99350 580224 99356
rect 456892 37936 456944 37942
rect 456892 37878 456944 37884
rect 582392 16574 582420 333231
rect 582484 133890 582512 556174
rect 582576 460222 582604 683839
rect 582564 460216 582616 460222
rect 582564 460158 582616 460164
rect 582562 458144 582618 458153
rect 582562 458079 582618 458088
rect 582576 145586 582604 458079
rect 582668 449206 582696 697167
rect 583206 670712 583262 670721
rect 583206 670647 583262 670656
rect 582746 630864 582802 630873
rect 582746 630799 582802 630808
rect 582760 554033 582788 630799
rect 582930 617536 582986 617545
rect 582930 617471 582986 617480
rect 582838 577688 582894 577697
rect 582838 577623 582894 577632
rect 582746 554024 582802 554033
rect 582746 553959 582802 553968
rect 582748 535492 582800 535498
rect 582748 535434 582800 535440
rect 582656 449200 582708 449206
rect 582656 449142 582708 449148
rect 582654 404968 582710 404977
rect 582654 404903 582710 404912
rect 582668 146985 582696 404903
rect 582760 298761 582788 535434
rect 582852 376689 582880 577623
rect 582944 543726 582972 617471
rect 583022 591016 583078 591025
rect 583022 590951 583078 590960
rect 582932 543720 582984 543726
rect 582932 543662 582984 543668
rect 582932 532024 582984 532030
rect 582932 531966 582984 531972
rect 582944 404977 582972 531966
rect 583036 496806 583064 590951
rect 583114 559056 583170 559065
rect 583114 558991 583170 559000
rect 583024 496800 583076 496806
rect 583024 496742 583076 496748
rect 583022 471472 583078 471481
rect 583022 471407 583078 471416
rect 582930 404968 582986 404977
rect 582930 404903 582986 404912
rect 582838 376680 582894 376689
rect 582838 376615 582894 376624
rect 583036 364313 583064 471407
rect 583128 458153 583156 558991
rect 583114 458144 583170 458153
rect 583114 458079 583170 458088
rect 583220 377369 583248 670647
rect 583300 465112 583352 465118
rect 583300 465054 583352 465060
rect 583312 418305 583340 465054
rect 583298 418296 583354 418305
rect 583298 418231 583354 418240
rect 583206 377360 583262 377369
rect 583206 377295 583262 377304
rect 583022 364304 583078 364313
rect 583022 364239 583078 364248
rect 582838 351928 582894 351937
rect 582838 351863 582894 351872
rect 582852 311001 582880 351863
rect 583022 325272 583078 325281
rect 583022 325207 583078 325216
rect 582838 310992 582894 311001
rect 582838 310927 582894 310936
rect 582746 298752 582802 298761
rect 582746 298687 582802 298696
rect 582930 298752 582986 298761
rect 582930 298687 582986 298696
rect 582746 272232 582802 272241
rect 582746 272167 582802 272176
rect 582760 206990 582788 272167
rect 582838 258904 582894 258913
rect 582838 258839 582894 258848
rect 582748 206984 582800 206990
rect 582748 206926 582800 206932
rect 582852 149054 582880 258839
rect 582944 193866 582972 298687
rect 583036 247625 583064 325207
rect 583298 312080 583354 312089
rect 583298 312015 583354 312024
rect 583114 310992 583170 311001
rect 583114 310927 583170 310936
rect 583128 310593 583156 310927
rect 583114 310584 583170 310593
rect 583114 310519 583170 310528
rect 583022 247616 583078 247625
rect 583022 247551 583078 247560
rect 583022 245576 583078 245585
rect 583022 245511 583078 245520
rect 583036 244934 583064 245511
rect 583024 244928 583076 244934
rect 583024 244870 583076 244876
rect 582932 193860 582984 193866
rect 582932 193802 582984 193808
rect 583036 151094 583064 244870
rect 583024 151088 583076 151094
rect 583024 151030 583076 151036
rect 582840 149048 582892 149054
rect 582840 148990 582892 148996
rect 582748 147008 582800 147014
rect 582654 146976 582710 146985
rect 582748 146950 582800 146956
rect 582654 146911 582710 146920
rect 582564 145580 582616 145586
rect 582564 145522 582616 145528
rect 582656 139460 582708 139466
rect 582656 139402 582708 139408
rect 582564 136672 582616 136678
rect 582564 136614 582616 136620
rect 582472 133884 582524 133890
rect 582472 133826 582524 133832
rect 582470 97200 582526 97209
rect 582470 97135 582526 97144
rect 582484 73001 582512 97135
rect 582470 72992 582526 73001
rect 582470 72927 582526 72936
rect 582576 19825 582604 136614
rect 582668 59673 582696 139402
rect 582760 125594 582788 146950
rect 583024 142180 583076 142186
rect 583024 142122 583076 142128
rect 582748 125588 582800 125594
rect 582748 125530 582800 125536
rect 583036 112849 583064 142122
rect 583128 126954 583156 310519
rect 583206 266384 583262 266393
rect 583312 266354 583340 312015
rect 583206 266319 583262 266328
rect 583300 266348 583352 266354
rect 583220 232393 583248 266319
rect 583300 266290 583352 266296
rect 583206 232384 583262 232393
rect 583206 232319 583262 232328
rect 583574 222864 583630 222873
rect 583574 222799 583630 222808
rect 583298 219056 583354 219065
rect 583298 218991 583354 219000
rect 583206 192536 583262 192545
rect 583206 192471 583262 192480
rect 583116 126948 583168 126954
rect 583116 126890 583168 126896
rect 583022 112840 583078 112849
rect 583022 112775 583078 112784
rect 583220 102134 583248 192471
rect 583312 144906 583340 218991
rect 583390 205728 583446 205737
rect 583390 205663 583446 205672
rect 583300 144900 583352 144906
rect 583300 144842 583352 144848
rect 583404 136610 583432 205663
rect 583482 178664 583538 178673
rect 583482 178599 583538 178608
rect 583392 136604 583444 136610
rect 583392 136546 583444 136552
rect 583496 124166 583524 178599
rect 583484 124160 583536 124166
rect 583484 124102 583536 124108
rect 583208 102128 583260 102134
rect 583208 102070 583260 102076
rect 582748 95260 582800 95266
rect 582748 95202 582800 95208
rect 582760 86193 582788 95202
rect 582840 93900 582892 93906
rect 582840 93842 582892 93848
rect 582746 86184 582802 86193
rect 582746 86119 582802 86128
rect 582654 59664 582710 59673
rect 582654 59599 582710 59608
rect 582852 33153 582880 93842
rect 583114 93120 583170 93129
rect 583114 93055 583170 93064
rect 583024 91792 583076 91798
rect 583024 91734 583076 91740
rect 583036 46345 583064 91734
rect 583022 46336 583078 46345
rect 583022 46271 583078 46280
rect 582838 33144 582894 33153
rect 582838 33079 582894 33088
rect 582562 19816 582618 19825
rect 582562 19751 582618 19760
rect 582392 16546 583064 16574
rect 449900 10328 449952 10334
rect 449900 10270 449952 10276
rect 582196 3528 582248 3534
rect 582196 3470 582248 3476
rect 583036 3482 583064 16546
rect 583128 6633 583156 93055
rect 583114 6624 583170 6633
rect 583114 6559 583170 6568
rect 583588 3534 583616 222799
rect 583758 196616 583814 196625
rect 583758 196551 583814 196560
rect 583666 152280 583722 152289
rect 583666 152215 583722 152224
rect 583680 99113 583708 152215
rect 583666 99104 583722 99113
rect 583666 99039 583722 99048
rect 583576 3528 583628 3534
rect 581000 3120 581052 3126
rect 581000 3062 581052 3068
rect 445852 2780 445904 2786
rect 445852 2722 445904 2728
rect 581012 480 581040 3062
rect 582208 480 582236 3470
rect 583036 3454 583432 3482
rect 583576 3470 583628 3476
rect 583404 480 583432 3454
rect 583772 3126 583800 196551
rect 583760 3120 583812 3126
rect 583760 3062 583812 3068
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 2778 658144 2834 658200
rect 3054 579944 3110 580000
rect 3238 566888 3294 566944
rect 2778 553852 2834 553888
rect 2778 553832 2780 553852
rect 2780 553832 2832 553852
rect 2832 553832 2834 553852
rect 3514 671200 3570 671256
rect 3514 632068 3516 632088
rect 3516 632068 3568 632088
rect 3568 632068 3570 632088
rect 3514 632032 3570 632068
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 4802 534656 4858 534712
rect 3422 527856 3478 527912
rect 2778 501744 2834 501800
rect 2778 462596 2834 462632
rect 2778 462576 2780 462596
rect 2780 462576 2832 462596
rect 2832 462576 2834 462596
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 3514 475632 3570 475688
rect 3146 449520 3202 449576
rect 22742 536016 22798 536072
rect 3422 423580 3424 423600
rect 3424 423580 3476 423600
rect 3476 423580 3478 423600
rect 3422 423544 3478 423580
rect 3422 410488 3478 410544
rect 3514 397432 3570 397488
rect 3422 389136 3478 389192
rect 4802 385600 4858 385656
rect 2962 371356 2964 371376
rect 2964 371356 3016 371376
rect 3016 371356 3018 371376
rect 2962 371320 3018 371356
rect 3422 358400 3478 358456
rect 3330 306176 3386 306232
rect 3146 267144 3202 267200
rect 3146 254088 3202 254144
rect 3330 241068 3332 241088
rect 3332 241068 3384 241088
rect 3384 241068 3386 241088
rect 3330 241032 3386 241068
rect 3330 214920 3386 214976
rect 3054 201864 3110 201920
rect 2778 188844 2780 188864
rect 2780 188844 2832 188864
rect 2832 188844 2834 188864
rect 2778 188808 2834 188844
rect 3330 162832 3386 162888
rect 3330 136720 3386 136776
rect 3146 110608 3202 110664
rect 3054 58520 3110 58576
rect 18 6704 74 6760
rect 3514 353912 3570 353968
rect 3606 345344 3662 345400
rect 7562 329840 7618 329896
rect 4066 319232 4122 319288
rect 3606 293120 3662 293176
rect 21362 335416 21418 335472
rect 11702 229064 11758 229120
rect 10966 227024 11022 227080
rect 15842 213152 15898 213208
rect 3606 149776 3662 149832
rect 3514 97552 3570 97608
rect 3514 84632 3570 84688
rect 12346 80688 12402 80744
rect 5446 79464 5502 79520
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 4066 36488 4122 36544
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 1674 4800 1730 4856
rect 10966 55800 11022 55856
rect 6826 39208 6882 39264
rect 13726 77832 13782 77888
rect 15106 76472 15162 76528
rect 18602 241440 18658 241496
rect 17866 190304 17922 190360
rect 17222 189080 17278 189136
rect 17866 189080 17922 189136
rect 39946 445712 40002 445768
rect 39302 329976 39358 330032
rect 29642 191664 29698 191720
rect 30286 191664 30342 191720
rect 29642 190440 29698 190496
rect 34426 83408 34482 83464
rect 26146 79328 26202 79384
rect 23386 64096 23442 64152
rect 19246 62736 19302 62792
rect 22006 53080 22062 53136
rect 30286 72392 30342 72448
rect 28906 35128 28962 35184
rect 31666 58520 31722 58576
rect 33046 47504 33102 47560
rect 44086 536016 44142 536072
rect 43994 382880 44050 382936
rect 35162 71848 35218 71904
rect 38566 65456 38622 65512
rect 35806 57160 35862 57216
rect 48226 539552 48282 539608
rect 48134 343576 48190 343632
rect 43442 233824 43498 233880
rect 44086 43424 44142 43480
rect 42706 11600 42762 11656
rect 49606 240080 49662 240136
rect 50894 66816 50950 66872
rect 48226 54440 48282 54496
rect 49606 39344 49662 39400
rect 52182 232600 52238 232656
rect 55126 444488 55182 444544
rect 55034 379344 55090 379400
rect 53654 241440 53710 241496
rect 56322 373224 56378 373280
rect 57886 447752 57942 447808
rect 57702 346976 57758 347032
rect 57610 335960 57666 336016
rect 56414 221992 56470 222048
rect 56506 219272 56562 219328
rect 58990 334600 59046 334656
rect 59082 332560 59138 332616
rect 54850 186224 54906 186280
rect 53746 75112 53802 75168
rect 53746 68176 53802 68232
rect 53654 50224 53710 50280
rect 52274 26152 52330 26208
rect 57794 59880 57850 59936
rect 58990 230424 59046 230480
rect 59266 371320 59322 371376
rect 59082 222128 59138 222184
rect 65982 590688 66038 590744
rect 61842 456048 61898 456104
rect 60462 338136 60518 338192
rect 61750 391312 61806 391368
rect 60646 374040 60702 374096
rect 60370 223352 60426 223408
rect 61750 338272 61806 338328
rect 65890 573416 65946 573472
rect 63222 391176 63278 391232
rect 63314 363704 63370 363760
rect 62762 338136 62818 338192
rect 62026 331880 62082 331936
rect 64694 454688 64750 454744
rect 66074 559544 66130 559600
rect 65798 393252 65800 393272
rect 65800 393252 65852 393272
rect 65852 393252 65854 393272
rect 65798 393216 65854 393252
rect 64694 388864 64750 388920
rect 66810 588376 66866 588432
rect 66258 586508 66260 586528
rect 66260 586508 66312 586528
rect 66312 586508 66314 586528
rect 66258 586472 66314 586508
rect 66902 585656 66958 585712
rect 66810 582936 66866 582992
rect 66534 581712 66590 581768
rect 66810 580216 66866 580272
rect 66810 576136 66866 576192
rect 67362 574912 67418 574968
rect 66810 572056 66866 572112
rect 67086 570696 67142 570752
rect 67454 570696 67510 570752
rect 67362 569336 67418 569392
rect 66810 567976 66866 568032
rect 66810 564984 66866 565040
rect 66810 563624 66866 563680
rect 66810 562264 66866 562320
rect 66810 560904 66866 560960
rect 66810 558184 66866 558240
rect 66810 555464 66866 555520
rect 66626 554104 66682 554160
rect 66810 550024 66866 550080
rect 66810 548664 66866 548720
rect 66810 547304 66866 547360
rect 66810 545944 66866 546000
rect 66810 544584 66866 544640
rect 66810 543224 66866 543280
rect 76746 593408 76802 593464
rect 73986 592048 74042 592104
rect 70306 590688 70362 590744
rect 71134 590688 71190 590744
rect 73066 590688 73122 590744
rect 74446 589872 74502 589928
rect 77666 589328 77722 589384
rect 82266 590960 82322 591016
rect 81898 590688 81954 590744
rect 81346 589464 81402 589520
rect 79690 588648 79746 588704
rect 86866 590824 86922 590880
rect 88062 588512 88118 588568
rect 67730 584296 67786 584352
rect 67638 566616 67694 566672
rect 67546 554104 67602 554160
rect 67454 552744 67510 552800
rect 67362 542952 67418 543008
rect 66994 541864 67050 541920
rect 66902 452512 66958 452568
rect 66074 424224 66130 424280
rect 66902 440000 66958 440056
rect 66902 437688 66958 437744
rect 66902 435240 66958 435296
rect 66810 433236 66812 433256
rect 66812 433236 66864 433256
rect 66864 433236 66866 433256
rect 66810 433200 66866 433236
rect 66534 431024 66590 431080
rect 66718 428576 66774 428632
rect 66258 426264 66314 426320
rect 66258 421912 66314 421968
rect 66902 417288 66958 417344
rect 66258 415112 66314 415168
rect 66350 408312 66406 408368
rect 66810 406136 66866 406192
rect 66626 403688 66682 403744
rect 66810 401512 66866 401568
rect 66810 399492 66866 399528
rect 66810 399472 66812 399492
rect 66812 399472 66864 399492
rect 66864 399472 66866 399492
rect 66994 396888 67050 396944
rect 67362 539416 67418 539472
rect 67546 551384 67602 551440
rect 67546 540504 67602 540560
rect 67546 539552 67602 539608
rect 89718 586200 89774 586256
rect 67822 577496 67878 577552
rect 88890 560088 88946 560144
rect 88798 540096 88854 540152
rect 67730 442176 67786 442232
rect 67454 412800 67510 412856
rect 67362 410488 67418 410544
rect 67362 396888 67418 396944
rect 67270 395936 67326 395992
rect 66166 387640 66222 387696
rect 65890 376624 65946 376680
rect 65982 351872 66038 351928
rect 63130 241984 63186 242040
rect 63222 231784 63278 231840
rect 64694 237904 64750 237960
rect 63314 208256 63370 208312
rect 65982 305224 66038 305280
rect 67362 347792 67418 347848
rect 67270 345752 67326 345808
rect 66258 326712 66314 326768
rect 67270 324536 67326 324592
rect 66534 322396 66536 322416
rect 66536 322396 66588 322416
rect 66588 322396 66590 322416
rect 66534 322360 66590 322396
rect 66810 320184 66866 320240
rect 66442 319096 66498 319152
rect 66442 318008 66498 318064
rect 66902 316920 66958 316976
rect 66810 314744 66866 314800
rect 66902 313928 66958 313984
rect 66166 312840 66222 312896
rect 66994 311752 67050 311808
rect 66810 309576 66866 309632
rect 66902 307400 66958 307456
rect 66810 306312 66866 306368
rect 66902 303048 66958 303104
rect 66810 301960 66866 302016
rect 66902 300872 66958 300928
rect 66626 298696 66682 298752
rect 66810 297608 66866 297664
rect 67086 310664 67142 310720
rect 66074 294344 66130 294400
rect 66810 293256 66866 293312
rect 66810 292168 66866 292224
rect 66350 289992 66406 290048
rect 66810 288904 66866 288960
rect 66258 286728 66314 286784
rect 66810 285640 66866 285696
rect 66810 284552 66866 284608
rect 66810 283464 66866 283520
rect 66626 279112 66682 279168
rect 66810 278024 66866 278080
rect 65890 274488 65946 274544
rect 65890 274080 65946 274136
rect 65982 259800 66038 259856
rect 65798 239944 65854 240000
rect 65982 232464 66038 232520
rect 66810 277208 66866 277264
rect 66258 276120 66314 276176
rect 66258 272856 66314 272912
rect 67178 296112 67234 296168
rect 67086 291100 67142 291136
rect 67086 291080 67088 291100
rect 67088 291080 67140 291100
rect 67140 291080 67142 291100
rect 67546 395936 67602 395992
rect 67546 394848 67602 394904
rect 69570 535472 69626 535528
rect 72606 536696 72662 536752
rect 73158 536016 73214 536072
rect 72606 454688 72662 454744
rect 70398 446392 70454 446448
rect 71778 445848 71834 445904
rect 76562 535336 76618 535392
rect 80058 535744 80114 535800
rect 81438 458904 81494 458960
rect 79414 444488 79470 444544
rect 83462 469784 83518 469840
rect 82818 456048 82874 456104
rect 82818 447752 82874 447808
rect 84198 447752 84254 447808
rect 82818 444488 82874 444544
rect 83830 444488 83886 444544
rect 86866 465704 86922 465760
rect 86958 457544 87014 457600
rect 89626 560088 89682 560144
rect 87602 444896 87658 444952
rect 90362 589872 90418 589928
rect 89810 567296 89866 567352
rect 89074 449112 89130 449168
rect 91098 587560 91154 587616
rect 91282 584840 91338 584896
rect 91834 583652 91836 583672
rect 91836 583652 91888 583672
rect 91888 583652 91890 583672
rect 91834 583616 91890 583652
rect 91282 582120 91338 582176
rect 91282 578040 91338 578096
rect 91190 576680 91246 576736
rect 91742 575320 91798 575376
rect 91742 573960 91798 574016
rect 91742 572600 91798 572656
rect 91190 571412 91192 571432
rect 91192 571412 91244 571432
rect 91244 571412 91246 571432
rect 91190 571376 91246 571412
rect 91742 568656 91798 568712
rect 91558 565836 91560 565856
rect 91560 565836 91612 565856
rect 91612 565836 91614 565856
rect 91558 565800 91614 565836
rect 91558 564460 91614 564496
rect 91558 564440 91560 564460
rect 91560 564440 91612 564460
rect 91612 564440 91614 564460
rect 91558 563100 91614 563136
rect 91558 563080 91560 563100
rect 91560 563080 91612 563100
rect 91612 563080 91614 563100
rect 91190 561448 91246 561504
rect 91098 557368 91154 557424
rect 91098 556008 91154 556064
rect 91098 552100 91100 552120
rect 91100 552100 91152 552120
rect 91152 552100 91154 552120
rect 91098 552064 91154 552100
rect 91098 550704 91154 550760
rect 91098 549344 91154 549400
rect 91098 547712 91154 547768
rect 91374 553288 91430 553344
rect 91282 547884 91284 547904
rect 91284 547884 91336 547904
rect 91336 547884 91338 547904
rect 91282 547848 91338 547884
rect 91558 545148 91614 545184
rect 91558 545128 91560 545148
rect 91560 545128 91612 545148
rect 91612 545128 91614 545148
rect 91558 542428 91614 542464
rect 91558 542408 91560 542428
rect 91560 542408 91612 542428
rect 91612 542408 91614 542428
rect 90546 468424 90602 468480
rect 90362 444624 90418 444680
rect 92294 558728 92350 558784
rect 91926 541048 91982 541104
rect 92386 538872 92442 538928
rect 93122 570016 93178 570072
rect 93766 543768 93822 543824
rect 93122 539688 93178 539744
rect 93766 538736 93822 538792
rect 93122 462848 93178 462904
rect 100758 593408 100814 593464
rect 95882 592048 95938 592104
rect 94594 541048 94650 541104
rect 94594 534656 94650 534712
rect 94594 467064 94650 467120
rect 95974 471144 96030 471200
rect 92478 446936 92534 446992
rect 93030 446936 93086 446992
rect 93030 445712 93086 445768
rect 94502 444760 94558 444816
rect 97262 590824 97318 590880
rect 100666 589464 100722 589520
rect 98642 589328 98698 589384
rect 97262 465704 97318 465760
rect 97906 457408 97962 457464
rect 96618 445848 96674 445904
rect 97630 445848 97686 445904
rect 98734 449928 98790 449984
rect 100482 445712 100538 445768
rect 104162 590960 104218 591016
rect 101402 468424 101458 468480
rect 105542 588648 105598 588704
rect 108394 469784 108450 469840
rect 105542 447072 105598 447128
rect 111062 449112 111118 449168
rect 109682 444896 109738 444952
rect 111706 444896 111762 444952
rect 118698 585656 118754 585712
rect 116122 448568 116178 448624
rect 113178 445712 113234 445768
rect 114374 445712 114430 445768
rect 117594 445712 117650 445768
rect 118514 445712 118570 445768
rect 120722 435920 120778 435976
rect 120722 417016 120778 417072
rect 120630 411032 120686 411088
rect 80058 390904 80114 390960
rect 80610 390904 80666 390960
rect 71870 390496 71926 390552
rect 68558 390224 68614 390280
rect 69938 390360 69994 390416
rect 69662 380160 69718 380216
rect 67638 337184 67694 337240
rect 71686 375400 71742 375456
rect 71042 368464 71098 368520
rect 70582 358808 70638 358864
rect 69846 331744 69902 331800
rect 71594 358808 71650 358864
rect 71778 340856 71834 340912
rect 72238 336776 72294 336832
rect 74538 388864 74594 388920
rect 73158 345616 73214 345672
rect 73066 340856 73122 340912
rect 73250 333240 73306 333296
rect 73250 332560 73306 332616
rect 79322 387640 79378 387696
rect 75826 366288 75882 366344
rect 73986 333240 74042 333296
rect 75182 333240 75238 333296
rect 70030 329296 70086 329352
rect 76562 349696 76618 349752
rect 75182 332288 75238 332344
rect 75826 332288 75882 332344
rect 75182 329432 75238 329488
rect 83922 388728 83978 388784
rect 80058 381520 80114 381576
rect 85854 391040 85910 391096
rect 105082 391040 105138 391096
rect 120906 442856 120962 442912
rect 121550 444760 121606 444816
rect 121550 444352 121606 444408
rect 121458 440000 121514 440056
rect 121458 428440 121514 428496
rect 121182 410488 121238 410544
rect 89810 390360 89866 390416
rect 91282 390360 91338 390416
rect 85578 368328 85634 368384
rect 86222 368328 86278 368384
rect 86222 367104 86278 367160
rect 85486 365744 85542 365800
rect 85394 360168 85450 360224
rect 82910 357584 82966 357640
rect 84106 357584 84162 357640
rect 79322 347112 79378 347168
rect 86222 360848 86278 360904
rect 81438 342216 81494 342272
rect 83002 333240 83058 333296
rect 84106 331880 84162 331936
rect 92754 390360 92810 390416
rect 91650 385736 91706 385792
rect 91098 384240 91154 384296
rect 90362 377984 90418 378040
rect 90914 339496 90970 339552
rect 94226 390360 94282 390416
rect 95882 390360 95938 390416
rect 97354 390360 97410 390416
rect 96250 387776 96306 387832
rect 98826 390360 98882 390416
rect 97722 386960 97778 387016
rect 94502 361664 94558 361720
rect 95054 361664 95110 361720
rect 92478 356088 92534 356144
rect 93674 356088 93730 356144
rect 93122 353368 93178 353424
rect 93214 340040 93270 340096
rect 96526 353912 96582 353968
rect 99194 356632 99250 356688
rect 97814 336096 97870 336152
rect 100666 390360 100722 390416
rect 102138 390360 102194 390416
rect 100850 389000 100906 389056
rect 101862 389000 101918 389056
rect 102322 389000 102378 389056
rect 103334 389000 103390 389056
rect 100482 387776 100538 387832
rect 100666 363024 100722 363080
rect 100666 354592 100722 354648
rect 100666 351192 100722 351248
rect 103702 388864 103758 388920
rect 115754 390632 115810 390688
rect 109682 390496 109738 390552
rect 106554 390360 106610 390416
rect 105542 386416 105598 386472
rect 104162 385600 104218 385656
rect 103426 383016 103482 383072
rect 101954 360304 102010 360360
rect 101862 349696 101918 349752
rect 102138 354728 102194 354784
rect 103426 354728 103482 354784
rect 108026 390360 108082 390416
rect 109774 389136 109830 389192
rect 112902 389000 112958 389056
rect 106186 349832 106242 349888
rect 111062 369824 111118 369880
rect 108946 363568 109002 363624
rect 113178 386280 113234 386336
rect 114374 386280 114430 386336
rect 114558 373360 114614 373416
rect 114466 367648 114522 367704
rect 107750 346296 107806 346352
rect 108302 346296 108358 346352
rect 107750 345072 107806 345128
rect 107474 343032 107530 343088
rect 106646 334056 106702 334112
rect 107842 332968 107898 333024
rect 109682 338408 109738 338464
rect 109682 333240 109738 333296
rect 110142 333240 110198 333296
rect 110418 347792 110474 347848
rect 111614 341400 111670 341456
rect 113178 360168 113234 360224
rect 114466 360168 114522 360224
rect 115938 390360 115994 390416
rect 116122 389000 116178 389056
rect 117134 389000 117190 389056
rect 117318 388864 117374 388920
rect 117870 390360 117926 390416
rect 118974 388864 119030 388920
rect 119986 385736 120042 385792
rect 116582 377848 116638 377904
rect 117134 377848 117190 377904
rect 116582 376896 116638 376952
rect 118606 365608 118662 365664
rect 118606 364384 118662 364440
rect 118514 364248 118570 364304
rect 116582 344256 116638 344312
rect 118330 343712 118386 343768
rect 115846 343612 115848 343632
rect 115848 343612 115900 343632
rect 115900 343612 115902 343632
rect 115846 343576 115902 343612
rect 115846 342896 115902 342952
rect 117226 337048 117282 337104
rect 119894 344256 119950 344312
rect 122286 444352 122342 444408
rect 122194 417968 122250 418024
rect 122838 423680 122894 423736
rect 122838 412800 122894 412856
rect 124126 444216 124182 444272
rect 124126 442040 124182 442096
rect 124126 437824 124182 437880
rect 124126 433236 124128 433256
rect 124128 433236 124180 433256
rect 124180 433236 124182 433256
rect 124126 433200 124182 433236
rect 124126 430636 124182 430672
rect 124126 430616 124128 430636
rect 124128 430616 124180 430636
rect 124180 430616 124182 430636
rect 123482 423680 123538 423736
rect 123022 419600 123078 419656
rect 122930 403688 122986 403744
rect 122930 392536 122986 392592
rect 124126 422048 124182 422104
rect 124126 415112 124182 415168
rect 124126 408468 124182 408504
rect 124126 408448 124128 408468
rect 124128 408448 124180 408468
rect 124180 408448 124182 408468
rect 123942 401512 123998 401568
rect 124126 399492 124182 399528
rect 124126 399472 124128 399492
rect 124128 399472 124180 399492
rect 124180 399472 124182 399492
rect 124126 396924 124128 396944
rect 124128 396924 124180 396944
rect 124180 396924 124182 396944
rect 124126 396888 124182 396924
rect 123758 392536 123814 392592
rect 126886 546488 126942 546544
rect 124310 406272 124366 406328
rect 124218 386280 124274 386336
rect 123482 370504 123538 370560
rect 123482 362344 123538 362400
rect 121734 349696 121790 349752
rect 121458 346976 121514 347032
rect 120722 346432 120778 346488
rect 120722 333240 120778 333296
rect 121826 332696 121882 332752
rect 124954 378664 125010 378720
rect 124862 347112 124918 347168
rect 124218 335552 124274 335608
rect 126242 348064 126298 348120
rect 124954 335416 125010 335472
rect 124862 332832 124918 332888
rect 125414 332832 125470 332888
rect 125414 329976 125470 330032
rect 129002 458224 129058 458280
rect 128174 352008 128230 352064
rect 154118 702480 154174 702536
rect 130474 536832 130530 536888
rect 130474 446936 130530 446992
rect 130382 444352 130438 444408
rect 129094 376760 129150 376816
rect 129646 376760 129702 376816
rect 129002 370504 129058 370560
rect 128358 349832 128414 349888
rect 126242 329840 126298 329896
rect 129738 369008 129794 369064
rect 132498 377848 132554 377904
rect 132406 369144 132462 369200
rect 129186 334600 129242 334656
rect 129738 331064 129794 331120
rect 134522 385600 134578 385656
rect 133142 370640 133198 370696
rect 133786 360440 133842 360496
rect 133694 347792 133750 347848
rect 135258 388728 135314 388784
rect 136638 378120 136694 378176
rect 134614 339632 134670 339688
rect 142066 542544 142122 542600
rect 141422 444624 141478 444680
rect 137926 378120 137982 378176
rect 139306 355408 139362 355464
rect 138018 351056 138074 351112
rect 136454 329840 136510 329896
rect 137282 336096 137338 336152
rect 139214 335416 139270 335472
rect 139398 339632 139454 339688
rect 140778 346568 140834 346624
rect 141422 346568 141478 346624
rect 142802 391176 142858 391232
rect 144734 363160 144790 363216
rect 141422 340992 141478 341048
rect 142066 340992 142122 341048
rect 142066 331880 142122 331936
rect 145286 330384 145342 330440
rect 145378 329840 145434 329896
rect 146206 334192 146262 334248
rect 146206 331880 146262 331936
rect 151082 362344 151138 362400
rect 150346 359488 150402 359544
rect 149058 346432 149114 346488
rect 149058 345616 149114 345672
rect 151082 356088 151138 356144
rect 151726 346432 151782 346488
rect 150530 337184 150586 337240
rect 150438 336912 150494 336968
rect 150438 335960 150494 336016
rect 150438 334464 150494 334520
rect 150438 334056 150494 334112
rect 149702 331200 149758 331256
rect 150254 331200 150310 331256
rect 151910 335688 151966 335744
rect 152462 332424 152518 332480
rect 151910 331744 151966 331800
rect 155314 448568 155370 448624
rect 155222 383016 155278 383072
rect 155222 356768 155278 356824
rect 153842 347928 153898 347984
rect 155222 345616 155278 345672
rect 153842 338544 153898 338600
rect 153198 337048 153254 337104
rect 153106 335688 153162 335744
rect 153198 334600 153254 334656
rect 153106 332832 153162 332888
rect 153106 331880 153162 331936
rect 153198 331064 153254 331120
rect 154486 338408 154542 338464
rect 154026 338000 154082 338056
rect 155222 333240 155278 333296
rect 155314 332424 155370 332480
rect 154854 331744 154910 331800
rect 153842 330520 153898 330576
rect 154118 329976 154174 330032
rect 155774 331744 155830 331800
rect 155774 331336 155830 331392
rect 169114 552064 169170 552120
rect 169114 539416 169170 539472
rect 156602 465160 156658 465216
rect 158074 386960 158130 387016
rect 156602 343848 156658 343904
rect 156878 343712 156934 343768
rect 155958 329840 156014 329896
rect 67822 323448 67878 323504
rect 157338 340992 157394 341048
rect 157982 338000 158038 338056
rect 157338 337320 157394 337376
rect 157982 333376 158038 333432
rect 156878 329704 156934 329760
rect 156878 328480 156934 328536
rect 156878 327664 156934 327720
rect 67730 308488 67786 308544
rect 67638 304136 67694 304192
rect 67546 299784 67602 299840
rect 67638 295432 67694 295488
rect 67454 291080 67510 291136
rect 67362 287836 67418 287872
rect 67362 287816 67364 287836
rect 67364 287816 67416 287836
rect 67416 287816 67418 287836
rect 67362 281288 67418 281344
rect 66994 273944 67050 274000
rect 66902 270680 66958 270736
rect 66810 268504 66866 268560
rect 66810 265240 66866 265296
rect 66902 264152 66958 264208
rect 66810 263064 66866 263120
rect 66258 261976 66314 262032
rect 66810 260924 66812 260944
rect 66812 260924 66864 260944
rect 66864 260924 66866 260944
rect 66810 260888 66866 260924
rect 66258 258068 66260 258088
rect 66260 258068 66312 258088
rect 66312 258068 66314 258088
rect 66258 258032 66314 258068
rect 66902 257624 66958 257680
rect 66810 255448 66866 255504
rect 66810 254360 66866 254416
rect 66810 253272 66866 253328
rect 67178 248920 67234 248976
rect 66810 246744 66866 246800
rect 66810 245676 66866 245712
rect 66810 245656 66812 245676
rect 66812 245656 66864 245676
rect 66864 245656 66866 245676
rect 66902 244568 66958 244624
rect 66074 226888 66130 226944
rect 66166 129240 66222 129296
rect 66166 128016 66222 128072
rect 64786 127064 64842 127120
rect 66166 127064 66222 127120
rect 64694 121488 64750 121544
rect 66166 126248 66222 126304
rect 66074 122576 66130 122632
rect 66074 121488 66130 121544
rect 66074 120808 66130 120864
rect 66166 94424 66222 94480
rect 66166 48864 66222 48920
rect 64786 44784 64842 44840
rect 67546 280220 67602 280256
rect 67546 280200 67548 280220
rect 67548 280200 67600 280220
rect 67600 280200 67602 280220
rect 67546 251096 67602 251152
rect 67270 243480 67326 243536
rect 67454 243480 67510 243536
rect 67546 243344 67602 243400
rect 67270 222808 67326 222864
rect 67730 282376 67786 282432
rect 67822 250008 67878 250064
rect 156694 242800 156750 242856
rect 80978 241984 81034 242040
rect 69754 241848 69810 241904
rect 69018 238312 69074 238368
rect 69938 241712 69994 241768
rect 69938 236544 69994 236600
rect 69662 206896 69718 206952
rect 71042 239944 71098 240000
rect 72422 240080 72478 240136
rect 71686 239400 71742 239456
rect 71042 215192 71098 215248
rect 72698 240080 72754 240136
rect 73066 224848 73122 224904
rect 74078 239672 74134 239728
rect 75550 239944 75606 240000
rect 77942 240760 77998 240816
rect 76562 220632 76618 220688
rect 77942 217368 77998 217424
rect 72422 195200 72478 195256
rect 154670 241984 154726 242040
rect 82818 237904 82874 237960
rect 82818 234504 82874 234560
rect 83554 239400 83610 239456
rect 84198 238176 84254 238232
rect 86866 215872 86922 215928
rect 85670 212472 85726 212528
rect 86866 212472 86922 212528
rect 83462 205536 83518 205592
rect 81346 200640 81402 200696
rect 87602 228248 87658 228304
rect 86866 198192 86922 198248
rect 89534 224712 89590 224768
rect 87602 196560 87658 196616
rect 89810 235864 89866 235920
rect 89810 234640 89866 234696
rect 90362 234640 90418 234696
rect 89718 209344 89774 209400
rect 91006 209344 91062 209400
rect 93858 241304 93914 241360
rect 92386 228792 92442 228848
rect 91190 227704 91246 227760
rect 92386 227704 92442 227760
rect 91098 206216 91154 206272
rect 92386 203496 92442 203552
rect 91006 202272 91062 202328
rect 90362 194112 90418 194168
rect 78678 193024 78734 193080
rect 93858 229064 93914 229120
rect 94916 241304 94972 241360
rect 94502 229064 94558 229120
rect 97446 239400 97502 239456
rect 97354 229744 97410 229800
rect 96526 225528 96582 225584
rect 95238 224984 95294 225040
rect 96526 224984 96582 225040
rect 94502 221856 94558 221912
rect 98366 239944 98422 240000
rect 102414 237224 102470 237280
rect 104714 235456 104770 235512
rect 102138 228248 102194 228304
rect 103426 228248 103482 228304
rect 100942 215056 100998 215112
rect 102046 215056 102102 215112
rect 100666 212336 100722 212392
rect 99286 208120 99342 208176
rect 103426 199416 103482 199472
rect 106278 234368 106334 234424
rect 104806 193840 104862 193896
rect 108164 241304 108220 241360
rect 109038 236680 109094 236736
rect 109682 229744 109738 229800
rect 111798 230288 111854 230344
rect 114282 232600 114338 232656
rect 113086 230288 113142 230344
rect 112994 217232 113050 217288
rect 109682 216416 109738 216472
rect 108302 213696 108358 213752
rect 114650 233144 114706 233200
rect 115938 226208 115994 226264
rect 115938 224984 115994 225040
rect 117134 224984 117190 225040
rect 115018 223488 115074 223544
rect 113086 196696 113142 196752
rect 107566 190984 107622 191040
rect 96526 189624 96582 189680
rect 95146 186904 95202 186960
rect 106186 185136 106242 185192
rect 100666 185000 100722 185056
rect 98826 182144 98882 182200
rect 93766 182008 93822 182064
rect 97262 179424 97318 179480
rect 98826 177520 98882 177576
rect 97262 176840 97318 176896
rect 102046 183640 102102 183696
rect 102046 177520 102102 177576
rect 108118 180784 108174 180840
rect 119894 231104 119950 231160
rect 117410 219136 117466 219192
rect 117318 210296 117374 210352
rect 121642 239672 121698 239728
rect 120078 202816 120134 202872
rect 122286 239536 122342 239592
rect 122102 236816 122158 236872
rect 122102 220768 122158 220824
rect 123482 209616 123538 209672
rect 122838 209480 122894 209536
rect 128266 215056 128322 215112
rect 129738 224576 129794 224632
rect 131026 224576 131082 224632
rect 129646 213560 129702 213616
rect 121366 199960 121422 200016
rect 119986 198056 120042 198112
rect 117226 195880 117282 195936
rect 117134 184184 117190 184240
rect 110694 179560 110750 179616
rect 106186 177520 106242 177576
rect 108118 177520 108174 177576
rect 110326 177520 110382 177576
rect 110694 177112 110750 177168
rect 114374 177520 114430 177576
rect 118606 177384 118662 177440
rect 122746 177520 122802 177576
rect 124034 177520 124090 177576
rect 125506 177520 125562 177576
rect 126886 177520 126942 177576
rect 133694 210976 133750 211032
rect 133142 205400 133198 205456
rect 135350 235728 135406 235784
rect 135258 230152 135314 230208
rect 136546 230152 136602 230208
rect 136822 237088 136878 237144
rect 137282 236680 137338 236736
rect 137282 235592 137338 235648
rect 138018 232600 138074 232656
rect 138018 230424 138074 230480
rect 138892 241440 138948 241496
rect 138662 220496 138718 220552
rect 136546 200776 136602 200832
rect 141422 215872 141478 215928
rect 141422 202136 141478 202192
rect 143446 241032 143502 241088
rect 142158 229064 142214 229120
rect 144182 228656 144238 228712
rect 144734 228248 144790 228304
rect 144090 227568 144146 227624
rect 143446 226208 143502 226264
rect 142802 216552 142858 216608
rect 145010 228520 145066 228576
rect 147770 225528 147826 225584
rect 147586 205264 147642 205320
rect 144918 204176 144974 204232
rect 142066 193160 142122 193216
rect 131026 183096 131082 183152
rect 149058 236544 149114 236600
rect 150806 240216 150862 240272
rect 149334 236000 149390 236056
rect 149334 232600 149390 232656
rect 149150 225936 149206 225992
rect 153106 241304 153162 241360
rect 153014 241168 153070 241224
rect 153382 240216 153438 240272
rect 152278 239944 152334 240000
rect 153106 239944 153162 240000
rect 153014 237360 153070 237416
rect 152738 231920 152794 231976
rect 153014 227568 153070 227624
rect 150346 217504 150402 217560
rect 150346 213696 150402 213752
rect 151082 213696 151138 213752
rect 153382 238584 153438 238640
rect 153290 237224 153346 237280
rect 153106 199280 153162 199336
rect 155682 240760 155738 240816
rect 154670 236952 154726 237008
rect 155682 235592 155738 235648
rect 155774 232464 155830 232520
rect 155774 231240 155830 231296
rect 154486 189760 154542 189816
rect 151082 187040 151138 187096
rect 156372 241440 156428 241496
rect 155958 237260 155960 237280
rect 155960 237260 156012 237280
rect 156012 237260 156014 237280
rect 155958 237224 156014 237260
rect 156510 220632 156566 220688
rect 158166 332696 158222 332752
rect 158074 300056 158130 300112
rect 157982 254496 158038 254552
rect 157338 240080 157394 240136
rect 158074 242120 158130 242176
rect 159362 341536 159418 341592
rect 158718 326440 158774 326496
rect 158902 324400 158958 324456
rect 158718 324264 158774 324320
rect 158810 323176 158866 323232
rect 158718 322088 158774 322144
rect 158718 321000 158774 321056
rect 158902 320728 158958 320784
rect 158718 319096 158774 319152
rect 158626 277752 158682 277808
rect 158626 261432 158682 261488
rect 158166 239944 158222 240000
rect 158626 234640 158682 234696
rect 157338 228792 157394 228848
rect 156602 202816 156658 202872
rect 158810 318824 158866 318880
rect 158810 315560 158866 315616
rect 158810 313384 158866 313440
rect 158902 311208 158958 311264
rect 158810 310120 158866 310176
rect 158810 307944 158866 308000
rect 158810 306856 158866 306912
rect 158810 305768 158866 305824
rect 158810 304680 158866 304736
rect 158810 303628 158812 303648
rect 158812 303628 158864 303648
rect 158864 303628 158866 303648
rect 158810 303592 158866 303628
rect 158810 301416 158866 301472
rect 158994 300348 159050 300384
rect 158994 300328 158996 300348
rect 158996 300328 159048 300348
rect 159048 300328 159050 300348
rect 158810 298152 158866 298208
rect 158810 297064 158866 297120
rect 158810 295996 158866 296032
rect 158810 295976 158812 295996
rect 158812 295976 158864 295996
rect 158864 295976 158866 295996
rect 158810 294888 158866 294944
rect 158902 293800 158958 293856
rect 158810 292984 158866 293040
rect 158810 291896 158866 291952
rect 158810 290808 158866 290864
rect 158902 289720 158958 289776
rect 158810 288632 158866 288688
rect 158810 287544 158866 287600
rect 158810 285368 158866 285424
rect 158810 284824 158866 284880
rect 158810 282104 158866 282160
rect 158810 281016 158866 281072
rect 160742 355272 160798 355328
rect 160098 336912 160154 336968
rect 160098 334736 160154 334792
rect 159638 334192 159694 334248
rect 159546 327528 159602 327584
rect 159730 328616 159786 328672
rect 159638 324944 159694 325000
rect 159730 323584 159786 323640
rect 160006 316684 160008 316704
rect 160008 316684 160060 316704
rect 160060 316684 160062 316704
rect 160006 316648 160062 316684
rect 159822 278840 159878 278896
rect 158810 276664 158866 276720
rect 158810 275576 158866 275632
rect 159546 274896 159602 274952
rect 158810 274488 158866 274544
rect 158810 273400 158866 273456
rect 158810 271224 158866 271280
rect 158810 269068 158866 269104
rect 158810 269048 158812 269068
rect 158812 269048 158864 269068
rect 158864 269048 158866 269068
rect 159362 267960 159418 268016
rect 158810 265784 158866 265840
rect 158810 264696 158866 264752
rect 158810 262520 158866 262576
rect 158902 260344 158958 260400
rect 158810 258168 158866 258224
rect 159270 257100 159326 257136
rect 159270 257080 159272 257100
rect 159272 257080 159324 257100
rect 159324 257080 159326 257100
rect 158810 256264 158866 256320
rect 158902 255176 158958 255232
rect 158810 254088 158866 254144
rect 158810 253000 158866 253056
rect 158902 251912 158958 251968
rect 158810 250824 158866 250880
rect 158810 249736 158866 249792
rect 158902 249192 158958 249248
rect 160834 334464 160890 334520
rect 160742 309848 160798 309904
rect 160098 284280 160154 284336
rect 159454 248648 159510 248704
rect 158810 246472 158866 246528
rect 158810 245384 158866 245440
rect 158810 244316 158866 244352
rect 158810 244296 158812 244316
rect 158812 244296 158864 244316
rect 158864 244296 158866 244316
rect 158810 243208 158866 243264
rect 159362 234640 159418 234696
rect 158718 233824 158774 233880
rect 158074 216280 158130 216336
rect 158718 210432 158774 210488
rect 160006 247560 160062 247616
rect 160834 294480 160890 294536
rect 160926 292440 160982 292496
rect 161478 363568 161534 363624
rect 161386 313928 161442 313984
rect 159546 235456 159602 235512
rect 160098 230444 160154 230480
rect 160098 230424 160100 230444
rect 160100 230424 160152 230444
rect 160152 230424 160154 230444
rect 159454 224848 159510 224904
rect 161018 238584 161074 238640
rect 161570 343712 161626 343768
rect 162122 329704 162178 329760
rect 161570 317736 161626 317792
rect 163502 369008 163558 369064
rect 162950 328208 163006 328264
rect 162766 289040 162822 289096
rect 162122 233280 162178 233336
rect 161386 230560 161442 230616
rect 161294 230424 161350 230480
rect 160834 193976 160890 194032
rect 162306 245656 162362 245712
rect 162214 231104 162270 231160
rect 163594 331744 163650 331800
rect 163594 301552 163650 301608
rect 164790 331880 164846 331936
rect 164882 318688 164938 318744
rect 164882 317328 164938 317384
rect 163594 235728 163650 235784
rect 164146 235728 164202 235784
rect 163778 231648 163834 231704
rect 166262 389136 166318 389192
rect 170402 527720 170458 527776
rect 168470 445712 168526 445768
rect 169022 445712 169078 445768
rect 168470 444488 168526 444544
rect 167734 341536 167790 341592
rect 167642 338272 167698 338328
rect 166998 318688 167054 318744
rect 166262 302368 166318 302424
rect 166078 301452 166080 301472
rect 166080 301452 166132 301472
rect 166132 301452 166134 301472
rect 166078 301416 166134 301452
rect 165066 246200 165122 246256
rect 164974 240760 165030 240816
rect 163778 210976 163834 211032
rect 162122 190304 162178 190360
rect 161386 188400 161442 188456
rect 165526 242936 165582 242992
rect 165250 242120 165306 242176
rect 165250 237088 165306 237144
rect 155866 181464 155922 181520
rect 148966 179288 149022 179344
rect 130934 177520 130990 177576
rect 132406 177520 132462 177576
rect 133786 177520 133842 177576
rect 148874 177520 148930 177576
rect 100666 176704 100722 176760
rect 103334 176704 103390 176760
rect 113730 176704 113786 176760
rect 115846 176704 115902 176760
rect 119526 176704 119582 176760
rect 120814 176704 120870 176760
rect 127070 176724 127126 176760
rect 127070 176704 127072 176724
rect 127072 176704 127124 176724
rect 127124 176704 127126 176724
rect 129462 176704 129518 176760
rect 158994 176740 158996 176760
rect 158996 176740 159048 176760
rect 159048 176740 159050 176760
rect 158994 176704 159050 176740
rect 134430 175344 134486 175400
rect 135718 175344 135774 175400
rect 163594 187176 163650 187232
rect 163502 176568 163558 176624
rect 166814 224712 166870 224768
rect 166814 224168 166870 224224
rect 166906 197920 166962 197976
rect 166262 179968 166318 180024
rect 165526 174936 165582 174992
rect 165434 174528 165490 174584
rect 164974 173168 165030 173224
rect 166446 179560 166502 179616
rect 67454 125160 67510 125216
rect 67362 123528 67418 123584
rect 67638 102312 67694 102368
rect 67546 100680 67602 100736
rect 100666 94696 100722 94752
rect 120630 94696 120686 94752
rect 106922 94424 106978 94480
rect 103426 93200 103482 93256
rect 85118 92384 85174 92440
rect 75274 91160 75330 91216
rect 86866 91296 86922 91352
rect 86774 91160 86830 91216
rect 70306 76608 70362 76664
rect 68926 71032 68982 71088
rect 70214 68312 70270 68368
rect 73066 73752 73122 73808
rect 75826 69536 75882 69592
rect 77206 66952 77262 67008
rect 79966 65592 80022 65648
rect 88062 91160 88118 91216
rect 89626 91160 89682 91216
rect 90730 91160 90786 91216
rect 91926 91160 91982 91216
rect 93030 91160 93086 91216
rect 95146 91160 95202 91216
rect 96342 91160 96398 91216
rect 90730 88168 90786 88224
rect 91926 86808 91982 86864
rect 93030 85312 93086 85368
rect 96342 88032 96398 88088
rect 95146 81368 95202 81424
rect 97814 91296 97870 91352
rect 97262 81232 97318 81288
rect 95146 77968 95202 78024
rect 87602 61376 87658 61432
rect 82082 1944 82138 2000
rect 85670 3304 85726 3360
rect 93766 51720 93822 51776
rect 97906 91160 97962 91216
rect 99194 91160 99250 91216
rect 97906 75248 97962 75304
rect 97814 73072 97870 73128
rect 101954 91296 102010 91352
rect 100666 91160 100722 91216
rect 102046 91160 102102 91216
rect 103334 91160 103390 91216
rect 104162 91432 104218 91488
rect 102046 62872 102102 62928
rect 106186 91296 106242 91352
rect 104438 91160 104494 91216
rect 106094 91160 106150 91216
rect 104438 85448 104494 85504
rect 105542 82592 105598 82648
rect 110142 93200 110198 93256
rect 108118 92384 108174 92440
rect 107566 91296 107622 91352
rect 107474 91160 107530 91216
rect 106922 84088 106978 84144
rect 108670 91160 108726 91216
rect 109222 91160 109278 91216
rect 110142 91160 110198 91216
rect 160742 94424 160798 94480
rect 118238 93472 118294 93528
rect 124126 93472 124182 93528
rect 111246 92384 111302 92440
rect 115754 92384 115810 92440
rect 116766 92384 116822 92440
rect 111338 91840 111394 91896
rect 112166 91160 112222 91216
rect 111338 89664 111394 89720
rect 112166 87896 112222 87952
rect 111706 76744 111762 76800
rect 111062 74432 111118 74488
rect 115478 92112 115534 92168
rect 113086 91160 113142 91216
rect 114374 91160 114430 91216
rect 116582 91840 116638 91896
rect 115478 90344 115534 90400
rect 120722 91840 120778 91896
rect 119894 91704 119950 91760
rect 117134 91160 117190 91216
rect 118054 91160 118110 91216
rect 119986 91160 120042 91216
rect 118054 85176 118110 85232
rect 117226 83544 117282 83600
rect 120722 82728 120778 82784
rect 119986 82456 120042 82512
rect 125782 92420 125784 92440
rect 125784 92420 125836 92440
rect 125836 92420 125838 92440
rect 125782 92384 125838 92420
rect 133142 92404 133198 92440
rect 133142 92384 133144 92404
rect 133144 92384 133196 92404
rect 133196 92384 133198 92404
rect 130750 91704 130806 91760
rect 151634 91704 151690 91760
rect 124034 91432 124090 91488
rect 122286 91160 122342 91216
rect 119986 73888 120042 73944
rect 121090 3440 121146 3496
rect 126794 91296 126850 91352
rect 124126 91160 124182 91216
rect 125414 91160 125470 91216
rect 126886 91160 126942 91216
rect 129646 91160 129702 91216
rect 126886 69672 126942 69728
rect 151542 91296 151598 91352
rect 132406 91160 132462 91216
rect 135166 91160 135222 91216
rect 136546 91160 136602 91216
rect 130750 89528 130806 89584
rect 132866 86672 132922 86728
rect 132406 78512 132462 78568
rect 151726 91160 151782 91216
rect 153106 91160 153162 91216
rect 162490 93336 162546 93392
rect 162122 93200 162178 93256
rect 147034 64232 147090 64288
rect 130382 19896 130438 19952
rect 144826 40568 144882 40624
rect 141422 28192 141478 28248
rect 132958 6160 133014 6216
rect 162214 88984 162270 89040
rect 162490 85176 162546 85232
rect 162214 82456 162270 82512
rect 166354 93064 166410 93120
rect 165066 92112 165122 92168
rect 166446 85312 166502 85368
rect 168286 345616 168342 345672
rect 167642 303592 167698 303648
rect 168286 298016 168342 298072
rect 167642 280064 167698 280120
rect 167642 262792 167698 262848
rect 167090 261704 167146 261760
rect 167090 254496 167146 254552
rect 167642 251776 167698 251832
rect 168194 249056 168250 249112
rect 168194 242800 168250 242856
rect 168562 370504 168618 370560
rect 168470 298016 168526 298072
rect 169574 346568 169630 346624
rect 168378 242120 168434 242176
rect 168286 235728 168342 235784
rect 168286 235184 168342 235240
rect 169574 278160 169630 278216
rect 169022 217504 169078 217560
rect 173254 535608 173310 535664
rect 171874 449928 171930 449984
rect 170586 355408 170642 355464
rect 170402 317328 170458 317384
rect 169758 301552 169814 301608
rect 169666 269184 169722 269240
rect 170402 269184 170458 269240
rect 171046 312432 171102 312488
rect 170862 267008 170918 267064
rect 170862 266328 170918 266384
rect 170494 255448 170550 255504
rect 170402 213152 170458 213208
rect 169022 200640 169078 200696
rect 167642 185136 167698 185192
rect 167734 175480 167790 175536
rect 167826 171536 167882 171592
rect 167734 165688 167790 165744
rect 169114 183640 169170 183696
rect 170402 179424 170458 179480
rect 171046 264968 171102 265024
rect 170954 255312 171010 255368
rect 171874 349832 171930 349888
rect 173806 382336 173862 382392
rect 172518 356768 172574 356824
rect 172426 338408 172482 338464
rect 172058 326304 172114 326360
rect 171966 311072 172022 311128
rect 171966 268368 172022 268424
rect 173162 339632 173218 339688
rect 171966 224576 172022 224632
rect 171782 224304 171838 224360
rect 170954 219136 171010 219192
rect 173714 321544 173770 321600
rect 173254 313248 173310 313304
rect 177302 536968 177358 537024
rect 174542 360440 174598 360496
rect 176106 376760 176162 376816
rect 174726 360440 174782 360496
rect 174634 344392 174690 344448
rect 173806 313248 173862 313304
rect 173714 276120 173770 276176
rect 173438 240488 173494 240544
rect 173162 231648 173218 231704
rect 172426 204856 172482 204912
rect 170862 185544 170918 185600
rect 167642 111696 167698 111752
rect 167734 110064 167790 110120
rect 167550 108704 167606 108760
rect 168378 90344 168434 90400
rect 167734 89528 167790 89584
rect 167642 88032 167698 88088
rect 170402 94424 170458 94480
rect 170402 91704 170458 91760
rect 169298 82592 169354 82648
rect 166998 6160 167054 6216
rect 173162 194112 173218 194168
rect 170770 93744 170826 93800
rect 174634 316784 174690 316840
rect 176014 348064 176070 348120
rect 174910 345072 174966 345128
rect 174818 309712 174874 309768
rect 175094 293936 175150 293992
rect 174726 271088 174782 271144
rect 174634 241440 174690 241496
rect 173806 208392 173862 208448
rect 173346 180784 173402 180840
rect 173254 172352 173310 172408
rect 175094 182008 175150 182064
rect 175094 181328 175150 181384
rect 173346 92248 173402 92304
rect 174542 94016 174598 94072
rect 174726 97008 174782 97064
rect 175922 234368 175978 234424
rect 176106 323720 176162 323776
rect 176658 349832 176714 349888
rect 176658 309848 176714 309904
rect 177394 363568 177450 363624
rect 177302 307672 177358 307728
rect 178038 379344 178094 379400
rect 178406 379344 178462 379400
rect 178406 378664 178462 378720
rect 178866 375400 178922 375456
rect 178774 366424 178830 366480
rect 178682 359488 178738 359544
rect 177854 353912 177910 353968
rect 177854 353504 177910 353560
rect 178682 336912 178738 336968
rect 177486 335552 177542 335608
rect 176014 217912 176070 217968
rect 175922 173848 175978 173904
rect 176106 178064 176162 178120
rect 176014 137400 176070 137456
rect 175922 88984 175978 89040
rect 175186 10240 175242 10296
rect 177578 307672 177634 307728
rect 177578 306992 177634 307048
rect 177486 247560 177542 247616
rect 177762 202836 177818 202872
rect 177762 202816 177764 202836
rect 177764 202816 177816 202836
rect 177816 202816 177818 202836
rect 177394 198192 177450 198248
rect 178038 228404 178094 228440
rect 178038 228384 178040 228404
rect 178040 228384 178092 228404
rect 178092 228384 178094 228404
rect 177578 177248 177634 177304
rect 178866 335960 178922 336016
rect 178866 273264 178922 273320
rect 178774 250416 178830 250472
rect 178774 236000 178830 236056
rect 184846 554784 184902 554840
rect 182822 533296 182878 533352
rect 180062 350512 180118 350568
rect 179418 320048 179474 320104
rect 180430 331200 180486 331256
rect 180246 320048 180302 320104
rect 180246 318824 180302 318880
rect 179418 241304 179474 241360
rect 178958 236000 179014 236056
rect 180062 231784 180118 231840
rect 180154 185000 180210 185056
rect 178866 182144 178922 182200
rect 180246 176840 180302 176896
rect 177486 91568 177542 91624
rect 177302 3984 177358 4040
rect 170402 3440 170458 3496
rect 178682 88168 178738 88224
rect 178038 86672 178094 86728
rect 178682 86128 178738 86184
rect 181626 354592 181682 354648
rect 181442 284960 181498 285016
rect 180522 241304 180578 241360
rect 180614 231784 180670 231840
rect 184202 539824 184258 539880
rect 183098 369824 183154 369880
rect 182822 336912 182878 336968
rect 182178 312432 182234 312488
rect 181626 273400 181682 273456
rect 182178 206760 182234 206816
rect 181626 200640 181682 200696
rect 181534 103808 181590 103864
rect 181442 93064 181498 93120
rect 181626 91024 181682 91080
rect 181534 84088 181590 84144
rect 181442 64232 181498 64288
rect 182914 305632 182970 305688
rect 183190 316648 183246 316704
rect 183006 283056 183062 283112
rect 183282 282920 183338 282976
rect 183466 287136 183522 287192
rect 185674 549344 185730 549400
rect 184846 447072 184902 447128
rect 184386 370504 184442 370560
rect 184294 345888 184350 345944
rect 184294 340040 184350 340096
rect 184294 318688 184350 318744
rect 184846 318688 184902 318744
rect 184846 317464 184902 317520
rect 184846 283192 184902 283248
rect 184386 283056 184442 283112
rect 184294 273400 184350 273456
rect 184202 267008 184258 267064
rect 183374 238448 183430 238504
rect 183282 231784 183338 231840
rect 183190 170992 183246 171048
rect 182914 87896 182970 87952
rect 184294 245792 184350 245848
rect 184846 247560 184902 247616
rect 184754 239672 184810 239728
rect 184754 238312 184810 238368
rect 184294 229744 184350 229800
rect 184662 191120 184718 191176
rect 185582 375944 185638 376000
rect 187054 556144 187110 556200
rect 185674 327800 185730 327856
rect 186226 295296 186282 295352
rect 185582 282104 185638 282160
rect 184938 235184 184994 235240
rect 187146 377304 187202 377360
rect 187146 363024 187202 363080
rect 187054 289720 187110 289776
rect 187054 289040 187110 289096
rect 187054 278024 187110 278080
rect 188894 538192 188950 538248
rect 188434 367104 188490 367160
rect 188342 360304 188398 360360
rect 187238 345752 187294 345808
rect 188986 534112 189042 534168
rect 188894 351192 188950 351248
rect 188342 320864 188398 320920
rect 187146 268504 187202 268560
rect 187238 264152 187294 264208
rect 186962 263744 187018 263800
rect 186226 245792 186282 245848
rect 186318 241304 186374 241360
rect 186226 182824 186282 182880
rect 184846 151000 184902 151056
rect 184386 118768 184442 118824
rect 185582 93336 185638 93392
rect 185766 86808 185822 86864
rect 187146 235592 187202 235648
rect 188342 307128 188398 307184
rect 188342 282784 188398 282840
rect 188342 265104 188398 265160
rect 188526 285096 188582 285152
rect 188342 234504 188398 234560
rect 187422 211928 187478 211984
rect 187054 188400 187110 188456
rect 188342 188400 188398 188456
rect 189722 332968 189778 333024
rect 191194 550840 191250 550896
rect 191746 534928 191802 534984
rect 191102 367784 191158 367840
rect 189906 340856 189962 340912
rect 189814 331880 189870 331936
rect 189722 244840 189778 244896
rect 189078 242256 189134 242312
rect 191102 297472 191158 297528
rect 190274 238312 190330 238368
rect 190182 220496 190238 220552
rect 190182 219408 190238 219464
rect 188986 212336 189042 212392
rect 187054 98640 187110 98696
rect 184294 26832 184350 26888
rect 184202 7520 184258 7576
rect 182822 6840 182878 6896
rect 190458 231240 190514 231296
rect 193954 550704 194010 550760
rect 192574 537104 192630 537160
rect 192666 451832 192722 451888
rect 191194 235184 191250 235240
rect 191654 246472 191710 246528
rect 191654 245656 191710 245712
rect 192206 245656 192262 245712
rect 192206 240216 192262 240272
rect 193126 382336 193182 382392
rect 192666 376760 192722 376816
rect 193954 338680 194010 338736
rect 194046 336776 194102 336832
rect 193126 293120 193182 293176
rect 192666 233824 192722 233880
rect 192942 233824 192998 233880
rect 192482 219408 192538 219464
rect 192574 218592 192630 218648
rect 191838 202136 191894 202192
rect 191838 197240 191894 197296
rect 191102 94424 191158 94480
rect 189722 28192 189778 28248
rect 191286 90888 191342 90944
rect 192942 220224 192998 220280
rect 193218 255312 193274 255368
rect 195242 542680 195298 542736
rect 195242 380160 195298 380216
rect 195242 378664 195298 378720
rect 194506 377440 194562 377496
rect 195242 362208 195298 362264
rect 195334 338136 195390 338192
rect 195242 329024 195298 329080
rect 194506 287408 194562 287464
rect 194414 255312 194470 255368
rect 193862 241440 193918 241496
rect 193862 215872 193918 215928
rect 195150 288496 195206 288552
rect 195150 285640 195206 285696
rect 195150 265512 195206 265568
rect 195150 264968 195206 265024
rect 194782 251776 194838 251832
rect 196714 541048 196770 541104
rect 195886 376080 195942 376136
rect 195886 368328 195942 368384
rect 195518 358808 195574 358864
rect 197082 470872 197138 470928
rect 196714 384920 196770 384976
rect 205638 559000 205694 559056
rect 198554 553968 198610 554024
rect 197450 532208 197506 532264
rect 197450 529796 197452 529816
rect 197452 529796 197504 529816
rect 197504 529796 197506 529816
rect 197450 529760 197506 529796
rect 198554 529760 198610 529816
rect 197450 527312 197506 527368
rect 197542 524728 197598 524784
rect 197450 522280 197506 522336
rect 197450 517384 197506 517440
rect 197450 510176 197506 510232
rect 197450 507592 197506 507648
rect 197450 502696 197506 502752
rect 198738 538328 198794 538384
rect 197450 500384 197506 500440
rect 198646 500384 198702 500440
rect 197450 495508 197506 495544
rect 197450 495488 197452 495508
rect 197452 495488 197504 495508
rect 197504 495488 197506 495508
rect 197450 492904 197506 492960
rect 197450 490456 197506 490512
rect 197450 488008 197506 488064
rect 197450 485560 197506 485616
rect 198002 483112 198058 483168
rect 197450 480664 197506 480720
rect 197450 478216 197506 478272
rect 197450 475768 197506 475824
rect 197450 473356 197452 473376
rect 197452 473356 197504 473376
rect 197504 473356 197506 473376
rect 197450 473320 197506 473356
rect 197450 468424 197506 468480
rect 197450 465976 197506 466032
rect 197450 463256 197506 463312
rect 197450 460844 197452 460864
rect 197452 460844 197504 460864
rect 197504 460844 197506 460864
rect 197450 460808 197506 460844
rect 197450 455912 197506 455968
rect 197358 448588 197414 448624
rect 197358 448568 197360 448588
rect 197360 448568 197412 448588
rect 197412 448568 197414 448588
rect 197358 446120 197414 446176
rect 197358 443708 197360 443728
rect 197360 443708 197412 443728
rect 197412 443708 197414 443728
rect 197358 443672 197414 443708
rect 197726 441396 197728 441416
rect 197728 441396 197780 441416
rect 197780 441396 197782 441416
rect 197726 441360 197782 441396
rect 197358 436328 197414 436384
rect 197358 433880 197414 433936
rect 197358 428984 197414 429040
rect 197358 426536 197414 426592
rect 197358 424088 197414 424144
rect 197358 419192 197414 419248
rect 197358 414296 197414 414352
rect 197358 411848 197414 411904
rect 197358 409536 197414 409592
rect 197358 406952 197414 407008
rect 197358 404504 197414 404560
rect 197358 399608 197414 399664
rect 197358 394732 197414 394768
rect 197358 394712 197360 394732
rect 197360 394712 197412 394732
rect 197412 394712 197414 394732
rect 197358 389952 197414 390008
rect 197358 387368 197414 387424
rect 197358 385076 197414 385112
rect 197358 385056 197360 385076
rect 197360 385056 197412 385076
rect 197412 385056 197414 385076
rect 197358 380180 197414 380216
rect 197358 380160 197360 380180
rect 197360 380160 197412 380180
rect 197412 380160 197414 380180
rect 196714 364248 196770 364304
rect 196714 346976 196770 347032
rect 196622 319368 196678 319424
rect 196714 314064 196770 314120
rect 195334 301688 195390 301744
rect 196622 287272 196678 287328
rect 195242 231920 195298 231976
rect 195242 231512 195298 231568
rect 195242 219136 195298 219192
rect 195794 241440 195850 241496
rect 195794 224848 195850 224904
rect 195426 221856 195482 221912
rect 195426 220088 195482 220144
rect 195242 202136 195298 202192
rect 195150 199416 195206 199472
rect 193862 196696 193918 196752
rect 193126 178608 193182 178664
rect 195242 198736 195298 198792
rect 195978 235728 196034 235784
rect 196070 233280 196126 233336
rect 196070 232464 196126 232520
rect 193954 110472 194010 110528
rect 194046 89664 194102 89720
rect 196898 254360 196954 254416
rect 196806 235864 196862 235920
rect 197082 251660 197138 251696
rect 197082 251640 197084 251660
rect 197084 251640 197136 251660
rect 197136 251640 197138 251660
rect 196898 232464 196954 232520
rect 196714 214648 196770 214704
rect 205638 550840 205694 550896
rect 199750 535336 199806 535392
rect 199750 533296 199806 533352
rect 199014 505144 199070 505200
rect 198830 463256 198886 463312
rect 198094 453464 198150 453520
rect 198646 421640 198702 421696
rect 198554 392264 198610 392320
rect 198002 318824 198058 318880
rect 198094 317600 198150 317656
rect 198370 307672 198426 307728
rect 198370 306448 198426 306504
rect 197358 282376 197414 282432
rect 197358 280744 197414 280800
rect 197450 280200 197506 280256
rect 197358 279384 197414 279440
rect 197266 250008 197322 250064
rect 197450 278568 197506 278624
rect 198370 278024 198426 278080
rect 197450 276664 197506 276720
rect 197542 275848 197598 275904
rect 197450 274488 197506 274544
rect 197450 272856 197506 272912
rect 197450 271496 197506 271552
rect 197450 270136 197506 270192
rect 197542 268776 197598 268832
rect 198278 267996 198280 268016
rect 198280 267996 198332 268016
rect 198332 267996 198334 268016
rect 198278 267960 198334 267996
rect 197542 267164 197598 267200
rect 197542 267144 197544 267164
rect 197544 267144 197596 267164
rect 197596 267144 197598 267164
rect 197450 266600 197506 266656
rect 197450 264424 197506 264480
rect 197450 263628 197506 263664
rect 197450 263608 197452 263628
rect 197452 263608 197504 263628
rect 197504 263608 197506 263628
rect 198462 262248 198518 262304
rect 197450 261432 197506 261488
rect 198094 260888 198150 260944
rect 197450 260072 197506 260128
rect 197450 259256 197506 259312
rect 197450 257896 197506 257952
rect 197542 257352 197598 257408
rect 197450 256536 197506 256592
rect 197450 255212 197452 255232
rect 197452 255212 197504 255232
rect 197504 255212 197506 255232
rect 197450 255176 197506 255212
rect 197910 253544 197966 253600
rect 197450 253000 197506 253056
rect 197450 250824 197506 250880
rect 197450 249500 197452 249520
rect 197452 249500 197504 249520
rect 197504 249500 197506 249520
rect 197450 249464 197506 249500
rect 197450 248684 197452 248704
rect 197452 248684 197504 248704
rect 197504 248684 197506 248704
rect 197450 248648 197506 248684
rect 197726 247832 197782 247888
rect 197358 245112 197414 245168
rect 197358 243752 197414 243808
rect 197910 240796 197912 240816
rect 197912 240796 197964 240816
rect 197964 240796 197966 240816
rect 197910 240760 197966 240796
rect 197174 180104 197230 180160
rect 196622 178744 196678 178800
rect 198922 416744 198978 416800
rect 198830 382472 198886 382528
rect 198738 278160 198794 278216
rect 198646 252184 198702 252240
rect 198646 246472 198702 246528
rect 198554 244296 198610 244352
rect 198462 242120 198518 242176
rect 201038 546624 201094 546680
rect 203614 541048 203670 541104
rect 231858 557504 231914 557560
rect 225326 545264 225382 545320
rect 217506 538192 217562 538248
rect 222474 538464 222530 538520
rect 223210 538464 223266 538520
rect 221094 538192 221150 538248
rect 208674 535472 208730 535528
rect 200394 535336 200450 535392
rect 201038 535336 201094 535392
rect 221094 535336 221150 535392
rect 255962 589328 256018 589384
rect 240230 554784 240286 554840
rect 243542 556144 243598 556200
rect 253938 550704 253994 550760
rect 255318 545128 255374 545184
rect 261758 542680 261814 542736
rect 262218 541184 262274 541240
rect 265530 538464 265586 538520
rect 273258 546624 273314 546680
rect 270682 539552 270738 539608
rect 273994 539552 274050 539608
rect 280618 539824 280674 539880
rect 283470 542544 283526 542600
rect 290094 552064 290150 552120
rect 304998 549344 305054 549400
rect 295338 546624 295394 546680
rect 298374 544040 298430 544096
rect 306654 543904 306710 543960
rect 318246 541184 318302 541240
rect 328458 547848 328514 547904
rect 323582 541456 323638 541512
rect 322018 539688 322074 539744
rect 339958 546488 340014 546544
rect 337106 538464 337162 538520
rect 335450 537104 335506 537160
rect 333794 536968 333850 537024
rect 348238 542408 348294 542464
rect 349986 541048 350042 541104
rect 356058 542444 356060 542464
rect 356060 542444 356112 542464
rect 356112 542444 356114 542464
rect 356058 542408 356114 542444
rect 353666 536832 353722 536888
rect 308402 535744 308458 535800
rect 276018 535608 276074 535664
rect 276938 535608 276994 535664
rect 304078 535472 304134 535528
rect 356242 538328 356298 538384
rect 357622 543768 357678 543824
rect 357530 540096 357586 540152
rect 357438 522280 357494 522336
rect 356334 519832 356390 519888
rect 357622 534656 357678 534712
rect 358726 532072 358782 532128
rect 358726 529624 358782 529680
rect 358726 527196 358782 527232
rect 358726 527176 358728 527196
rect 358728 527176 358780 527196
rect 358780 527176 358782 527196
rect 358726 524728 358782 524784
rect 358726 522280 358782 522336
rect 358634 519832 358690 519888
rect 358726 517384 358782 517440
rect 357530 512624 357586 512680
rect 358082 510040 358138 510096
rect 356242 490864 356298 490920
rect 357898 482840 357954 482896
rect 357898 477944 357954 478000
rect 358726 507592 358782 507648
rect 358726 505164 358782 505200
rect 358726 505144 358728 505164
rect 358728 505144 358780 505164
rect 358780 505144 358782 505164
rect 358726 502696 358782 502752
rect 358726 497800 358782 497856
rect 358634 495488 358690 495544
rect 358726 492904 358782 492960
rect 358726 487736 358782 487792
rect 358174 485288 358230 485344
rect 358726 475496 358782 475552
rect 358726 473048 358782 473104
rect 358726 470620 358782 470656
rect 358726 470600 358728 470620
rect 358728 470600 358780 470620
rect 358780 470600 358782 470620
rect 356242 467880 356298 467936
rect 358726 465704 358782 465760
rect 358634 463256 358690 463312
rect 358726 460808 358782 460864
rect 357438 458360 357494 458416
rect 201314 377576 201370 377632
rect 200026 376488 200082 376544
rect 200210 367784 200266 367840
rect 200118 310392 200174 310448
rect 199474 272312 199530 272368
rect 201406 362208 201462 362264
rect 200394 291896 200450 291952
rect 201406 304952 201462 305008
rect 200486 290944 200542 291000
rect 201590 377440 201646 377496
rect 202234 375944 202290 376000
rect 202878 363704 202934 363760
rect 202142 291352 202198 291408
rect 200486 284008 200542 284064
rect 202142 284824 202198 284880
rect 205730 376080 205786 376136
rect 205822 366424 205878 366480
rect 208398 366288 208454 366344
rect 203614 293120 203670 293176
rect 202878 291896 202934 291952
rect 204902 295432 204958 295488
rect 203154 289720 203210 289776
rect 204258 289720 204314 289776
rect 204258 289176 204314 289232
rect 204258 284960 204314 285016
rect 206374 315288 206430 315344
rect 207754 338680 207810 338736
rect 207662 305768 207718 305824
rect 206466 298016 206522 298072
rect 207570 298016 207626 298072
rect 206650 297472 206706 297528
rect 206282 296656 206338 296712
rect 205178 285640 205234 285696
rect 204902 284824 204958 284880
rect 207570 296792 207626 296848
rect 206098 284280 206154 284336
rect 207754 291080 207810 291136
rect 209134 369144 209190 369200
rect 215206 375128 215262 375184
rect 214562 374040 214618 374096
rect 211894 351192 211950 351248
rect 209134 327800 209190 327856
rect 210974 317328 211030 317384
rect 210606 310528 210662 310584
rect 209962 289040 210018 289096
rect 211434 305632 211490 305688
rect 211434 303728 211490 303784
rect 210606 289040 210662 289096
rect 211894 338680 211950 338736
rect 213274 359488 213330 359544
rect 213182 314880 213238 314936
rect 212354 292712 212410 292768
rect 211986 289720 212042 289776
rect 211986 288496 212042 288552
rect 213366 306992 213422 307048
rect 214654 308624 214710 308680
rect 213182 289720 213238 289776
rect 218242 376760 218298 376816
rect 218242 375128 218298 375184
rect 215298 350376 215354 350432
rect 215298 349968 215354 350024
rect 215298 305768 215354 305824
rect 214746 299512 214802 299568
rect 214562 296656 214618 296712
rect 215390 293800 215446 293856
rect 215390 292712 215446 292768
rect 215298 288360 215354 288416
rect 215298 287544 215354 287600
rect 215206 287408 215262 287464
rect 216034 349968 216090 350024
rect 216034 330520 216090 330576
rect 220818 371320 220874 371376
rect 221462 371320 221518 371376
rect 218702 370776 218758 370832
rect 216034 288360 216090 288416
rect 216678 287680 216734 287736
rect 218058 289040 218114 289096
rect 217322 287272 217378 287328
rect 217230 285776 217286 285832
rect 215942 285640 215998 285696
rect 217690 287136 217746 287192
rect 221462 353912 221518 353968
rect 222842 343712 222898 343768
rect 218518 284416 218574 284472
rect 221462 320864 221518 320920
rect 220174 306992 220230 307048
rect 220174 295432 220230 295488
rect 220818 295432 220874 295488
rect 220082 290944 220138 291000
rect 220174 288496 220230 288552
rect 221186 292712 221242 292768
rect 223026 298696 223082 298752
rect 223026 289856 223082 289912
rect 222842 285776 222898 285832
rect 205362 283872 205418 283928
rect 214470 283872 214526 283928
rect 216126 283872 216182 283928
rect 220266 283872 220322 283928
rect 225694 315288 225750 315344
rect 230478 365744 230534 365800
rect 231122 365744 231178 365800
rect 229098 362480 229154 362536
rect 227718 351328 227774 351384
rect 226982 319368 227038 319424
rect 226338 297472 226394 297528
rect 226706 296928 226762 296984
rect 225694 294072 225750 294128
rect 226890 294072 226946 294128
rect 226706 291080 226762 291136
rect 223946 285640 224002 285696
rect 225602 288360 225658 288416
rect 225050 285640 225106 285696
rect 225970 285776 226026 285832
rect 227442 316648 227498 316704
rect 227442 316104 227498 316160
rect 226982 291216 227038 291272
rect 227626 291216 227682 291272
rect 227902 292440 227958 292496
rect 227902 292032 227958 292088
rect 228454 292032 228510 292088
rect 233146 362344 233202 362400
rect 232502 361664 232558 361720
rect 233146 361664 233202 361720
rect 232226 320592 232282 320648
rect 231122 306448 231178 306504
rect 230294 301688 230350 301744
rect 231122 297472 231178 297528
rect 230386 297336 230442 297392
rect 223762 283872 223818 283928
rect 232686 328616 232742 328672
rect 233882 323720 233938 323776
rect 232686 320592 232742 320648
rect 232686 320184 232742 320240
rect 232502 289040 232558 289096
rect 232778 292576 232834 292632
rect 234618 314744 234674 314800
rect 234526 298152 234582 298208
rect 233698 290400 233754 290456
rect 232778 288496 232834 288552
rect 234250 287136 234306 287192
rect 234526 290944 234582 291000
rect 235354 345888 235410 345944
rect 238022 364384 238078 364440
rect 237378 344392 237434 344448
rect 235998 322088 236054 322144
rect 235354 314744 235410 314800
rect 236642 308488 236698 308544
rect 235998 285640 236054 285696
rect 241426 375264 241482 375320
rect 241426 374040 241482 374096
rect 248050 374040 248106 374096
rect 245658 370640 245714 370696
rect 246302 360168 246358 360224
rect 244922 357584 244978 357640
rect 242162 356632 242218 356688
rect 238114 324944 238170 325000
rect 238114 286048 238170 286104
rect 237286 285912 237342 285968
rect 236642 285776 236698 285832
rect 237378 284960 237434 285016
rect 237654 285912 237710 285968
rect 237654 285504 237710 285560
rect 239034 309712 239090 309768
rect 240230 290400 240286 290456
rect 241426 288632 241482 288688
rect 242254 330384 242310 330440
rect 243082 287136 243138 287192
rect 242898 285640 242954 285696
rect 243082 286048 243138 286104
rect 243082 284144 243138 284200
rect 244278 328344 244334 328400
rect 244278 327664 244334 327720
rect 244278 315016 244334 315072
rect 244278 313928 244334 313984
rect 243542 285640 243598 285696
rect 243818 284824 243874 284880
rect 243818 284280 243874 284336
rect 242990 284008 243046 284064
rect 229466 283872 229522 283928
rect 230938 283872 230994 283928
rect 236734 283872 236790 283928
rect 200118 283464 200174 283520
rect 244002 279928 244058 279984
rect 245014 356632 245070 356688
rect 245014 344392 245070 344448
rect 245658 334736 245714 334792
rect 245014 328344 245070 328400
rect 244922 311072 244978 311128
rect 244370 278024 244426 278080
rect 244278 269592 244334 269648
rect 247038 334600 247094 334656
rect 246302 324944 246358 325000
rect 245658 294480 245714 294536
rect 244922 273400 244978 273456
rect 244462 268776 244518 268832
rect 244462 264424 244518 264480
rect 244370 261704 244426 261760
rect 244002 259256 244058 259312
rect 199474 250416 199530 250472
rect 200026 249464 200082 249520
rect 198738 237360 198794 237416
rect 198462 229744 198518 229800
rect 199934 242256 199990 242312
rect 199842 240216 199898 240272
rect 199934 240080 199990 240136
rect 199382 228792 199438 228848
rect 198370 195336 198426 195392
rect 244002 244160 244058 244216
rect 200118 240488 200174 240544
rect 200118 240080 200174 240136
rect 200578 239672 200634 239728
rect 200118 237224 200174 237280
rect 201590 238312 201646 238368
rect 201314 237088 201370 237144
rect 201314 235728 201370 235784
rect 201314 235184 201370 235240
rect 198002 186224 198058 186280
rect 197266 115096 197322 115152
rect 198002 100000 198058 100056
rect 198002 82184 198058 82240
rect 199382 113328 199438 113384
rect 198186 110472 198242 110528
rect 198186 74432 198242 74488
rect 199474 87488 199530 87544
rect 202142 238448 202198 238504
rect 202050 234368 202106 234424
rect 202510 234368 202566 234424
rect 202326 227024 202382 227080
rect 202510 227024 202566 227080
rect 202234 185544 202290 185600
rect 202142 112376 202198 112432
rect 201130 93744 201186 93800
rect 202234 88984 202290 89040
rect 202142 30232 202198 30288
rect 204074 235864 204130 235920
rect 205822 238584 205878 238640
rect 205362 237224 205418 237280
rect 204442 228792 204498 228848
rect 204442 227704 204498 227760
rect 203614 127200 203670 127256
rect 203522 123528 203578 123584
rect 203614 95784 203670 95840
rect 204994 227704 205050 227760
rect 204994 211792 205050 211848
rect 204902 95784 204958 95840
rect 203706 81368 203762 81424
rect 204994 84768 205050 84824
rect 207110 216416 207166 216472
rect 207110 215328 207166 215384
rect 207294 206216 207350 206272
rect 207938 240080 207994 240136
rect 208306 240080 208362 240136
rect 208306 238176 208362 238232
rect 208858 235728 208914 235784
rect 208858 234912 208914 234968
rect 209042 237224 209098 237280
rect 208950 227568 209006 227624
rect 208950 221856 209006 221912
rect 207938 216008 207994 216064
rect 207754 215328 207810 215384
rect 207018 187176 207074 187232
rect 206558 181600 206614 181656
rect 209226 234912 209282 234968
rect 209870 239400 209926 239456
rect 210698 240080 210754 240136
rect 209870 238312 209926 238368
rect 209962 237360 210018 237416
rect 209778 215192 209834 215248
rect 209042 206216 209098 206272
rect 209226 206216 209282 206272
rect 211250 238584 211306 238640
rect 210698 237360 210754 237416
rect 211250 237360 211306 237416
rect 210422 234504 210478 234560
rect 213090 240080 213146 240136
rect 210422 220088 210478 220144
rect 210514 215192 210570 215248
rect 209962 205400 210018 205456
rect 210422 205400 210478 205456
rect 209042 203496 209098 203552
rect 207754 177384 207810 177440
rect 206374 136720 206430 136776
rect 206466 91840 206522 91896
rect 206282 86264 206338 86320
rect 207754 85448 207810 85504
rect 209226 115096 209282 115152
rect 210514 203496 210570 203552
rect 211802 185680 211858 185736
rect 214194 240080 214250 240136
rect 213826 239536 213882 239592
rect 213826 238448 213882 238504
rect 214194 238312 214250 238368
rect 213826 217368 213882 217424
rect 213826 210976 213882 211032
rect 213182 208256 213238 208312
rect 210514 174528 210570 174584
rect 210514 131280 210570 131336
rect 209226 91024 209282 91080
rect 210606 82728 210662 82784
rect 214470 205692 214526 205728
rect 214470 205672 214472 205692
rect 214472 205672 214524 205692
rect 214524 205672 214526 205692
rect 215942 224984 215998 225040
rect 215298 216008 215354 216064
rect 215298 214512 215354 214568
rect 215298 185000 215354 185056
rect 216034 206896 216090 206952
rect 216586 237360 216642 237416
rect 216770 237360 216826 237416
rect 217506 240080 217562 240136
rect 217506 237360 217562 237416
rect 218150 234640 218206 234696
rect 218150 230288 218206 230344
rect 218150 229064 218206 229120
rect 218150 228248 218206 228304
rect 218058 221992 218114 222048
rect 218058 218592 218114 218648
rect 217138 216008 217194 216064
rect 218978 240080 219034 240136
rect 220910 240116 220912 240136
rect 220912 240116 220964 240136
rect 220964 240116 220966 240136
rect 220910 240080 220966 240116
rect 220726 239808 220782 239864
rect 219530 231648 219586 231704
rect 218978 230288 219034 230344
rect 221002 233144 221058 233200
rect 220358 231648 220414 231704
rect 220174 231240 220230 231296
rect 216770 200912 216826 200968
rect 216034 199416 216090 199472
rect 217322 185816 217378 185872
rect 213918 175616 213974 175672
rect 214102 175480 214158 175536
rect 213918 174936 213974 174992
rect 214010 174256 214066 174312
rect 213918 172896 213974 172952
rect 214562 177112 214618 177168
rect 214470 173576 214526 173632
rect 214194 172216 214250 172272
rect 214102 171536 214158 171592
rect 214010 171012 214066 171048
rect 214010 170992 214012 171012
rect 214012 170992 214064 171012
rect 214064 170992 214066 171012
rect 213918 170312 213974 170368
rect 213918 169652 213974 169688
rect 213918 169632 213920 169652
rect 213920 169632 213972 169652
rect 213972 169632 213974 169652
rect 214010 168952 214066 169008
rect 213918 168308 213920 168328
rect 213920 168308 213972 168328
rect 213972 168308 213974 168328
rect 213918 168272 213974 168308
rect 214010 167592 214066 167648
rect 213918 166932 213974 166968
rect 213918 166912 213920 166932
rect 213920 166912 213972 166932
rect 213972 166912 213974 166932
rect 214010 166368 214066 166424
rect 213918 165008 213974 165064
rect 213918 163648 213974 163704
rect 214010 162968 214066 163024
rect 213918 162288 213974 162344
rect 214010 161744 214066 161800
rect 213918 161064 213974 161120
rect 214010 160384 214066 160440
rect 213918 159704 213974 159760
rect 215482 175888 215538 175944
rect 215206 173168 215262 173224
rect 215390 173848 215446 173904
rect 215482 172352 215538 172408
rect 216770 179424 216826 179480
rect 216678 178064 216734 178120
rect 216034 177520 216090 177576
rect 216678 176568 216734 176624
rect 218794 187720 218850 187776
rect 221462 237224 221518 237280
rect 221646 233144 221702 233200
rect 223394 233180 223396 233200
rect 223396 233180 223448 233200
rect 223448 233180 223450 233200
rect 223394 233144 223450 233180
rect 221646 225664 221702 225720
rect 222382 215228 222384 215248
rect 222384 215228 222436 215248
rect 222436 215228 222438 215248
rect 222382 215192 222438 215228
rect 223394 211112 223450 211168
rect 223394 210296 223450 210352
rect 224314 240080 224370 240136
rect 224314 237360 224370 237416
rect 224774 238720 224830 238776
rect 226706 238448 226762 238504
rect 226706 237904 226762 237960
rect 226154 234640 226210 234696
rect 225786 231104 225842 231160
rect 225234 217912 225290 217968
rect 225602 217368 225658 217424
rect 224406 215872 224462 215928
rect 225234 215872 225290 215928
rect 225694 209480 225750 209536
rect 225694 200912 225750 200968
rect 225694 184456 225750 184512
rect 228362 240080 228418 240136
rect 228178 221992 228234 222048
rect 227626 219272 227682 219328
rect 227074 218048 227130 218104
rect 227626 218048 227682 218104
rect 227074 203632 227130 203688
rect 227074 180240 227130 180296
rect 226338 180104 226394 180160
rect 226246 176704 226302 176760
rect 227810 185000 227866 185056
rect 227718 176160 227774 176216
rect 229098 238040 229154 238096
rect 228454 215056 228510 215112
rect 230570 240080 230626 240136
rect 230478 238040 230534 238096
rect 229650 213832 229706 213888
rect 230570 237360 230626 237416
rect 232502 240080 232558 240136
rect 231766 237360 231822 237416
rect 231490 234504 231546 234560
rect 230478 213560 230534 213616
rect 230386 206760 230442 206816
rect 226246 175888 226302 175944
rect 229006 175888 229062 175944
rect 229190 176432 229246 176488
rect 229098 175208 229154 175264
rect 229098 174664 229154 174720
rect 215942 170856 215998 170912
rect 215206 164328 215262 164384
rect 214562 159024 214618 159080
rect 213918 158344 213974 158400
rect 214010 157664 214066 157720
rect 213918 157120 213974 157176
rect 214010 156440 214066 156496
rect 213918 155796 213920 155816
rect 213920 155796 213972 155816
rect 213972 155796 213974 155816
rect 213918 155760 213974 155796
rect 214010 155080 214066 155136
rect 214010 154400 214066 154456
rect 213918 153720 213974 153776
rect 213918 153040 213974 153096
rect 214010 152496 214066 152552
rect 214562 151816 214618 151872
rect 214010 151136 214066 151192
rect 213918 150476 213974 150512
rect 213918 150456 213920 150476
rect 213920 150456 213972 150476
rect 213972 150456 213974 150476
rect 213918 149776 213974 149832
rect 214010 149096 214066 149152
rect 213918 148416 213974 148472
rect 213918 147872 213974 147928
rect 214010 147192 214066 147248
rect 213918 146512 213974 146568
rect 213918 145152 213974 145208
rect 214194 144472 214250 144528
rect 213918 143792 213974 143848
rect 214010 143248 214066 143304
rect 213918 142568 213974 142624
rect 214010 141888 214066 141944
rect 213918 141208 213974 141264
rect 213918 140528 213974 140584
rect 230386 179324 230388 179344
rect 230388 179324 230440 179344
rect 230440 179324 230442 179344
rect 230386 179288 230442 179324
rect 229466 177248 229522 177304
rect 229374 176296 229430 176352
rect 229466 173984 229522 174040
rect 229374 173304 229430 173360
rect 229190 170856 229246 170912
rect 230018 176568 230074 176624
rect 230478 174664 230534 174720
rect 230570 173712 230626 173768
rect 229558 161880 229614 161936
rect 229098 148688 229154 148744
rect 229834 157800 229890 157856
rect 229742 147192 229798 147248
rect 213918 139168 213974 139224
rect 214102 138624 214158 138680
rect 213366 137944 213422 138000
rect 213274 103536 213330 103592
rect 189722 3304 189778 3360
rect 209042 3304 209098 3360
rect 214010 135904 214066 135960
rect 213918 135224 213974 135280
rect 213918 134544 213974 134600
rect 214562 139848 214618 139904
rect 213918 133320 213974 133376
rect 214470 132640 214526 132696
rect 213918 131960 213974 132016
rect 213918 130600 213974 130656
rect 214010 129920 214066 129976
rect 213918 129240 213974 129296
rect 213918 128016 213974 128072
rect 213918 125976 213974 126032
rect 213918 125296 213974 125352
rect 214102 128696 214158 128752
rect 214010 124072 214066 124128
rect 213918 123392 213974 123448
rect 214102 123528 214158 123584
rect 215942 136584 215998 136640
rect 214746 126656 214802 126712
rect 214010 122712 214066 122768
rect 213918 122032 213974 122088
rect 214010 121352 214066 121408
rect 213918 120672 213974 120728
rect 214010 119992 214066 120048
rect 213918 119448 213974 119504
rect 214010 118088 214066 118144
rect 213918 117428 213974 117464
rect 213918 117408 213920 117428
rect 213920 117408 213972 117428
rect 213972 117408 213974 117428
rect 214010 116728 214066 116784
rect 213918 116068 213974 116104
rect 213918 116048 213920 116068
rect 213920 116048 213972 116068
rect 213972 116048 213974 116068
rect 214010 115368 214066 115424
rect 213918 114824 213974 114880
rect 213918 114144 213974 114200
rect 214010 112784 214066 112840
rect 213918 112104 213974 112160
rect 214010 111424 214066 111480
rect 213918 110744 213974 110800
rect 214010 110200 214066 110256
rect 213918 109520 213974 109576
rect 214010 108840 214066 108896
rect 213918 108160 213974 108216
rect 214010 107480 214066 107536
rect 213918 106800 213974 106856
rect 214010 106120 214066 106176
rect 213918 105576 213974 105632
rect 213918 102196 213974 102232
rect 213918 102176 213920 102196
rect 213920 102176 213972 102196
rect 213972 102176 213974 102196
rect 214010 101496 214066 101552
rect 213918 100952 213974 101008
rect 213918 99592 213974 99648
rect 214010 98912 214066 98968
rect 213918 98232 213974 98288
rect 213918 96872 213974 96928
rect 215022 124616 215078 124672
rect 214746 104896 214802 104952
rect 214930 100272 214986 100328
rect 214838 96328 214894 96384
rect 216126 133864 216182 133920
rect 216034 95784 216090 95840
rect 215942 93880 215998 93936
rect 214930 93200 214986 93256
rect 215942 90344 215998 90400
rect 216310 100000 216366 100056
rect 216678 98640 216734 98696
rect 219162 95920 219218 95976
rect 224314 93880 224370 93936
rect 223026 82048 223082 82104
rect 228454 95240 228510 95296
rect 228362 87488 228418 87544
rect 228454 79464 228510 79520
rect 230754 170448 230810 170504
rect 231858 234096 231914 234152
rect 231950 217368 232006 217424
rect 234066 238720 234122 238776
rect 232502 214376 232558 214432
rect 231766 178200 231822 178256
rect 230846 169904 230902 169960
rect 231674 172352 231730 172408
rect 231398 171808 231454 171864
rect 231766 171400 231822 171456
rect 230938 168544 230994 168600
rect 230938 164328 230994 164384
rect 231030 163784 231086 163840
rect 231674 170312 231730 170368
rect 231490 167592 231546 167648
rect 231306 166096 231362 166152
rect 231490 165180 231492 165200
rect 231492 165180 231544 165200
rect 231544 165180 231546 165200
rect 231490 165144 231546 165180
rect 231398 165008 231454 165064
rect 231122 162832 231178 162888
rect 231030 160520 231086 160576
rect 230662 157664 230718 157720
rect 231214 156576 231270 156632
rect 230570 155216 230626 155272
rect 231214 154808 231270 154864
rect 231306 154400 231362 154456
rect 230570 153040 230626 153096
rect 230570 151952 230626 152008
rect 230478 151580 230480 151600
rect 230480 151580 230532 151600
rect 230532 151580 230534 151600
rect 230478 151544 230534 151580
rect 229834 117000 229890 117056
rect 229834 114824 229890 114880
rect 231214 153312 231270 153368
rect 230662 151000 230718 151056
rect 230570 147736 230626 147792
rect 230570 146240 230626 146296
rect 230570 140120 230626 140176
rect 231766 169532 231768 169552
rect 231768 169532 231820 169552
rect 231820 169532 231822 169552
rect 231766 169496 231822 169532
rect 231766 168952 231822 169008
rect 231766 168000 231822 168056
rect 231766 166676 231768 166696
rect 231768 166676 231820 166696
rect 231820 166676 231822 166696
rect 231766 166640 231822 166676
rect 231674 164736 231730 164792
rect 231674 161472 231730 161528
rect 231766 160656 231822 160712
rect 232134 206760 232190 206816
rect 231766 159976 231822 160032
rect 231766 158652 231768 158672
rect 231768 158652 231820 158672
rect 231820 158652 231822 158672
rect 231766 158616 231822 158652
rect 231490 158072 231546 158128
rect 231674 157936 231730 157992
rect 231674 157120 231730 157176
rect 231766 156712 231822 156768
rect 231766 155760 231822 155816
rect 231766 155216 231822 155272
rect 231766 154264 231822 154320
rect 231398 153856 231454 153912
rect 231766 153856 231822 153912
rect 231766 152904 231822 152960
rect 231674 151000 231730 151056
rect 231490 148280 231546 148336
rect 231490 144880 231546 144936
rect 233514 234640 233570 234696
rect 233514 231240 233570 231296
rect 234066 226208 234122 226264
rect 233422 220768 233478 220824
rect 234986 231648 235042 231704
rect 235354 222128 235410 222184
rect 232502 164872 232558 164928
rect 231766 146784 231822 146840
rect 231766 146104 231822 146160
rect 231766 143928 231822 143984
rect 231674 143384 231730 143440
rect 231766 142432 231822 142488
rect 231214 141616 231270 141672
rect 231306 135904 231362 135960
rect 231214 133048 231270 133104
rect 231766 138216 231822 138272
rect 231582 136856 231638 136912
rect 231766 136312 231822 136368
rect 231490 135360 231546 135416
rect 231766 135088 231822 135144
rect 231766 134408 231822 134464
rect 231490 134000 231546 134056
rect 231766 133456 231822 133512
rect 231674 132504 231730 132560
rect 231122 131144 231178 131200
rect 231398 130192 231454 130248
rect 231306 129784 231362 129840
rect 231490 129784 231546 129840
rect 231398 128832 231454 128888
rect 231306 127336 231362 127392
rect 230754 125976 230810 126032
rect 230570 123528 230626 123584
rect 230018 122032 230074 122088
rect 229926 113192 229982 113248
rect 230662 120264 230718 120320
rect 231214 123392 231270 123448
rect 230938 121624 230994 121680
rect 231122 120128 231178 120184
rect 230938 117952 230994 118008
rect 231030 117408 231086 117464
rect 230754 116048 230810 116104
rect 230662 114552 230718 114608
rect 230938 112648 230994 112704
rect 230754 110744 230810 110800
rect 231766 131552 231822 131608
rect 231766 130600 231822 130656
rect 231766 129240 231822 129296
rect 231766 128308 231822 128344
rect 231766 128288 231768 128308
rect 231768 128288 231820 128308
rect 231820 128288 231822 128308
rect 231674 127880 231730 127936
rect 231582 127608 231638 127664
rect 231766 126928 231822 126984
rect 231674 126384 231730 126440
rect 232502 125432 232558 125488
rect 231766 125296 231822 125352
rect 231766 124480 231822 124536
rect 231582 124072 231638 124128
rect 231766 123120 231822 123176
rect 231766 122168 231822 122224
rect 231766 121216 231822 121272
rect 231674 120672 231730 120728
rect 232502 120400 232558 120456
rect 231306 119312 231362 119368
rect 231766 118904 231822 118960
rect 231766 118360 231822 118416
rect 231582 117952 231638 118008
rect 231490 116456 231546 116512
rect 231490 115096 231546 115152
rect 231398 113736 231454 113792
rect 231306 107888 231362 107944
rect 231306 105576 231362 105632
rect 231214 105168 231270 105224
rect 231122 103264 231178 103320
rect 230754 102312 230810 102368
rect 230570 101768 230626 101824
rect 230938 100680 230994 100736
rect 230938 99456 230994 99512
rect 231122 98640 231178 98696
rect 230570 96600 230626 96656
rect 230478 96192 230534 96248
rect 230018 88984 230074 89040
rect 229834 57160 229890 57216
rect 231306 102720 231362 102776
rect 231306 102176 231362 102232
rect 231766 114144 231822 114200
rect 231674 113600 231730 113656
rect 231766 112240 231822 112296
rect 231582 111696 231638 111752
rect 231766 111288 231822 111344
rect 231490 111016 231546 111072
rect 231674 109792 231730 109848
rect 231766 109384 231822 109440
rect 231766 108432 231822 108488
rect 231766 107072 231822 107128
rect 231674 106528 231730 106584
rect 231582 106156 231584 106176
rect 231584 106156 231636 106176
rect 231636 106156 231638 106176
rect 231582 106120 231638 106156
rect 231674 104660 231676 104680
rect 231676 104660 231728 104680
rect 231728 104660 231730 104680
rect 231674 104624 231730 104660
rect 231766 103672 231822 103728
rect 231490 101496 231546 101552
rect 231398 101360 231454 101416
rect 231306 98504 231362 98560
rect 231582 100816 231638 100872
rect 231766 100408 231822 100464
rect 231674 99864 231730 99920
rect 231766 98912 231822 98968
rect 231674 97960 231730 98016
rect 231490 97552 231546 97608
rect 231766 97008 231822 97064
rect 231674 96636 231676 96656
rect 231676 96636 231728 96656
rect 231728 96636 231730 96656
rect 231674 96600 231730 96636
rect 231766 96464 231822 96520
rect 231214 94424 231270 94480
rect 232686 112104 232742 112160
rect 232870 120128 232926 120184
rect 236366 239944 236422 240000
rect 237470 240080 237526 240136
rect 236550 235728 236606 235784
rect 236458 235592 236514 235648
rect 235906 206896 235962 206952
rect 235354 170448 235410 170504
rect 236090 177520 236146 177576
rect 234618 166776 234674 166832
rect 234250 163376 234306 163432
rect 234158 160384 234214 160440
rect 233974 119040 234030 119096
rect 233882 105168 233938 105224
rect 232686 82184 232742 82240
rect 235262 136992 235318 137048
rect 234158 119720 234214 119776
rect 233974 76608 234030 76664
rect 236090 160928 236146 160984
rect 237378 235456 237434 235512
rect 237930 235456 237986 235512
rect 236734 156576 236790 156632
rect 236642 146920 236698 146976
rect 236642 138352 236698 138408
rect 236826 146648 236882 146704
rect 238298 236952 238354 237008
rect 238298 230288 238354 230344
rect 237562 210432 237618 210488
rect 239402 228520 239458 228576
rect 238758 220224 238814 220280
rect 240690 237224 240746 237280
rect 240046 233824 240102 233880
rect 240690 230424 240746 230480
rect 242162 240080 242218 240136
rect 241794 237360 241850 237416
rect 242806 237360 242862 237416
rect 242714 237088 242770 237144
rect 242622 236816 242678 236872
rect 241242 233824 241298 233880
rect 239402 205536 239458 205592
rect 239770 205536 239826 205592
rect 238022 204176 238078 204232
rect 237562 162424 237618 162480
rect 237470 159568 237526 159624
rect 238206 128968 238262 129024
rect 238850 180240 238906 180296
rect 238390 129784 238446 129840
rect 239402 125296 239458 125352
rect 239402 123120 239458 123176
rect 238298 110744 238354 110800
rect 239586 153176 239642 153232
rect 242806 231784 242862 231840
rect 243634 239944 243690 240000
rect 242990 209616 243046 209672
rect 240782 178064 240838 178120
rect 240322 170312 240378 170368
rect 240782 169768 240838 169824
rect 240782 168408 240838 168464
rect 240138 149096 240194 149152
rect 240782 142976 240838 143032
rect 239678 124752 239734 124808
rect 239586 117952 239642 118008
rect 239586 102856 239642 102912
rect 240874 123392 240930 123448
rect 241702 173984 241758 174040
rect 241518 150048 241574 150104
rect 241518 142860 241574 142896
rect 241518 142840 241520 142860
rect 241520 142840 241572 142860
rect 241572 142840 241574 142860
rect 242990 170448 243046 170504
rect 242898 167048 242954 167104
rect 242346 149640 242402 149696
rect 241058 109384 241114 109440
rect 241058 75248 241114 75304
rect 242254 111016 242310 111072
rect 242438 145832 242494 145888
rect 243634 167048 243690 167104
rect 243174 155216 243230 155272
rect 243542 140664 243598 140720
rect 242438 113872 242494 113928
rect 242254 107616 242310 107672
rect 244370 210432 244426 210488
rect 246302 289992 246358 290048
rect 245750 276684 245806 276720
rect 245750 276664 245752 276684
rect 245752 276664 245804 276684
rect 245804 276664 245806 276684
rect 248418 295976 248474 296032
rect 246946 283736 247002 283792
rect 246302 283192 246358 283248
rect 245934 281560 245990 281616
rect 246118 281016 246174 281072
rect 245934 279384 245990 279440
rect 245934 278840 245990 278896
rect 245934 277480 245990 277536
rect 245934 275848 245990 275904
rect 245934 275324 245990 275360
rect 245934 275304 245936 275324
rect 245936 275304 245988 275324
rect 245988 275304 245990 275324
rect 245842 274488 245898 274544
rect 245842 273164 245844 273184
rect 245844 273164 245896 273184
rect 245896 273164 245898 273184
rect 245842 273128 245898 273164
rect 245934 272312 245990 272368
rect 245934 271496 245990 271552
rect 245842 270952 245898 271008
rect 245934 270172 245936 270192
rect 245936 270172 245988 270192
rect 245988 270172 245990 270192
rect 245934 270136 245990 270172
rect 245750 266600 245806 266656
rect 245842 265784 245898 265840
rect 245842 262268 245898 262304
rect 245842 262248 245844 262268
rect 245844 262248 245896 262268
rect 245896 262248 245898 262268
rect 245658 259528 245714 259584
rect 245658 258712 245714 258768
rect 245842 258168 245898 258224
rect 245842 257352 245898 257408
rect 245842 256536 245898 256592
rect 245842 256028 245844 256048
rect 245844 256028 245896 256048
rect 245896 256028 245898 256048
rect 245842 255992 245898 256028
rect 245842 255196 245898 255232
rect 245842 255176 245844 255196
rect 245844 255176 245896 255196
rect 245896 255176 245898 255196
rect 245658 253816 245714 253872
rect 245842 252220 245844 252240
rect 245844 252220 245896 252240
rect 245896 252220 245898 252240
rect 245842 252184 245898 252220
rect 245658 250824 245714 250880
rect 245842 247288 245898 247344
rect 245658 245928 245714 245984
rect 245750 243752 245806 243808
rect 245658 241576 245714 241632
rect 245842 240760 245898 240816
rect 245750 214784 245806 214840
rect 245658 178608 245714 178664
rect 244370 169768 244426 169824
rect 244462 165008 244518 165064
rect 243818 154808 243874 154864
rect 243634 117544 243690 117600
rect 244922 150864 244978 150920
rect 244278 142432 244334 142488
rect 246302 269592 246358 269648
rect 246026 265240 246082 265296
rect 246026 260072 246082 260128
rect 246026 254360 246082 254416
rect 246026 253000 246082 253056
rect 246026 251640 246082 251696
rect 246026 249464 246082 249520
rect 246026 245112 246082 245168
rect 247222 282376 247278 282432
rect 247130 260888 247186 260944
rect 246118 242392 246174 242448
rect 245934 172760 245990 172816
rect 246302 171672 246358 171728
rect 247130 248648 247186 248704
rect 246302 157936 246358 157992
rect 245750 148144 245806 148200
rect 245658 138760 245714 138816
rect 245014 99456 245070 99512
rect 243634 50224 243690 50280
rect 177394 1944 177450 2000
rect 244094 4936 244150 4992
rect 246486 153720 246542 153776
rect 246394 132776 246450 132832
rect 246302 115504 246358 115560
rect 245198 68312 245254 68368
rect 245106 64096 245162 64152
rect 247682 285096 247738 285152
rect 247314 250280 247370 250336
rect 247314 239808 247370 239864
rect 247222 223488 247278 223544
rect 247222 159024 247278 159080
rect 247130 151000 247186 151056
rect 246578 137128 246634 137184
rect 248602 273164 248604 273184
rect 248604 273164 248656 273184
rect 248656 273164 248658 273184
rect 248602 273128 248658 273164
rect 249154 309984 249210 310040
rect 249890 232600 249946 232656
rect 248510 187720 248566 187776
rect 251914 353368 251970 353424
rect 250626 302368 250682 302424
rect 250534 285776 250590 285832
rect 251086 282784 251142 282840
rect 251086 251776 251142 251832
rect 250534 213152 250590 213208
rect 247774 143112 247830 143168
rect 247774 124616 247830 124672
rect 247038 86264 247094 86320
rect 246394 71032 246450 71088
rect 248418 123392 248474 123448
rect 247958 110336 248014 110392
rect 247958 108024 248014 108080
rect 245658 3848 245714 3904
rect 249890 185408 249946 185464
rect 251270 272992 251326 273048
rect 251270 270408 251326 270464
rect 254582 356632 254638 356688
rect 253294 355272 253350 355328
rect 253202 349832 253258 349888
rect 251822 247016 251878 247072
rect 251822 225664 251878 225720
rect 251822 207576 251878 207632
rect 251270 204992 251326 205048
rect 251178 144064 251234 144120
rect 249154 75112 249210 75168
rect 250442 98368 250498 98424
rect 250626 109248 250682 109304
rect 250810 124752 250866 124808
rect 250626 62872 250682 62928
rect 250534 58520 250590 58576
rect 247590 3304 247646 3360
rect 247774 3304 247830 3360
rect 249982 15136 250038 15192
rect 252098 168952 252154 169008
rect 255962 349832 256018 349888
rect 255410 311072 255466 311128
rect 254030 298016 254086 298072
rect 254582 298016 254638 298072
rect 254030 297336 254086 297392
rect 253846 288496 253902 288552
rect 253202 286320 253258 286376
rect 253294 284960 253350 285016
rect 252834 275712 252890 275768
rect 253110 245792 253166 245848
rect 253846 282104 253902 282160
rect 253294 269184 253350 269240
rect 253294 172760 253350 172816
rect 253202 156712 253258 156768
rect 252558 153040 252614 153096
rect 253386 148280 253442 148336
rect 252098 77968 252154 78024
rect 252006 59880 252062 59936
rect 251914 47504 251970 47560
rect 254122 287680 254178 287736
rect 254030 213832 254086 213888
rect 255410 240216 255466 240272
rect 255410 179424 255466 179480
rect 255318 171672 255374 171728
rect 253938 139712 253994 139768
rect 253386 108976 253442 109032
rect 254582 125976 254638 126032
rect 253294 65456 253350 65512
rect 254582 55800 254638 55856
rect 260838 367784 260894 367840
rect 258722 329024 258778 329080
rect 257342 313248 257398 313304
rect 256790 300056 256846 300112
rect 258170 301416 258226 301472
rect 257526 283600 257582 283656
rect 257342 277480 257398 277536
rect 257526 264832 257582 264888
rect 258078 264832 258134 264888
rect 257434 231104 257490 231160
rect 259458 322088 259514 322144
rect 258906 288632 258962 288688
rect 258814 264696 258870 264752
rect 259366 264696 259422 264752
rect 258722 243480 258778 243536
rect 259366 237904 259422 237960
rect 258814 234368 258870 234424
rect 259274 178608 259330 178664
rect 257342 174256 257398 174312
rect 258722 169768 258778 169824
rect 255962 102176 256018 102232
rect 255962 72392 256018 72448
rect 257342 127608 257398 127664
rect 256054 66816 256110 66872
rect 257342 102176 257398 102232
rect 256238 76744 256294 76800
rect 256146 48864 256202 48920
rect 258814 142568 258870 142624
rect 258722 132368 258778 132424
rect 258078 109656 258134 109712
rect 258078 109248 258134 109304
rect 257526 86128 257582 86184
rect 257434 73888 257490 73944
rect 258906 130192 258962 130248
rect 258906 107072 258962 107128
rect 259734 245792 259790 245848
rect 260746 245792 260802 245848
rect 260930 291352 260986 291408
rect 262126 312568 262182 312624
rect 264242 374040 264298 374096
rect 262310 331744 262366 331800
rect 262218 301552 262274 301608
rect 261482 266328 261538 266384
rect 261482 263472 261538 263528
rect 261574 237904 261630 237960
rect 260838 196696 260894 196752
rect 263690 351056 263746 351112
rect 262862 292712 262918 292768
rect 262770 247016 262826 247072
rect 262310 231104 262366 231160
rect 263598 282784 263654 282840
rect 261482 174392 261538 174448
rect 260102 170176 260158 170232
rect 260286 159024 260342 159080
rect 258906 65592 258962 65648
rect 252558 30232 252614 30288
rect 251914 9424 251970 9480
rect 251822 3576 251878 3632
rect 252374 3576 252430 3632
rect 262126 167184 262182 167240
rect 261482 142704 261538 142760
rect 261666 140800 261722 140856
rect 260194 69536 260250 69592
rect 261666 101496 261722 101552
rect 262862 163240 262918 163296
rect 264242 344256 264298 344312
rect 264242 318824 264298 318880
rect 263782 218592 263838 218648
rect 264978 206896 265034 206952
rect 264978 175616 265034 175672
rect 265070 175208 265126 175264
rect 264978 174800 265034 174856
rect 265254 173984 265310 174040
rect 265070 173576 265126 173632
rect 264978 172624 265034 172680
rect 264242 172352 264298 172408
rect 265254 172352 265310 172408
rect 263598 163376 263654 163432
rect 262862 122712 262918 122768
rect 262862 116864 262918 116920
rect 262862 116048 262918 116104
rect 261666 79328 261722 79384
rect 265070 172216 265126 172272
rect 264978 171400 265034 171456
rect 265162 171808 265218 171864
rect 265070 170992 265126 171048
rect 264978 170040 265034 170096
rect 265162 169768 265218 169824
rect 265070 169632 265126 169688
rect 264978 168816 265034 168872
rect 265438 168408 265494 168464
rect 265346 167864 265402 167920
rect 264978 167456 265034 167512
rect 265070 166640 265126 166696
rect 264978 166232 265034 166288
rect 265162 165824 265218 165880
rect 265070 165280 265126 165336
rect 264978 164464 265034 164520
rect 265162 164872 265218 164928
rect 265254 164056 265310 164112
rect 265070 163648 265126 163704
rect 264978 162832 265034 162888
rect 265070 162288 265126 162344
rect 265162 161472 265218 161528
rect 264978 161064 265034 161120
rect 264978 159704 265034 159760
rect 267002 305632 267058 305688
rect 265714 290400 265770 290456
rect 267186 299512 267242 299568
rect 267738 320728 267794 320784
rect 268382 284144 268438 284200
rect 267738 221992 267794 222048
rect 270406 352008 270462 352064
rect 269854 296928 269910 296984
rect 269762 235864 269818 235920
rect 267830 219136 267886 219192
rect 269026 221992 269082 222048
rect 269762 186360 269818 186416
rect 269946 237088 270002 237144
rect 270406 235864 270462 235920
rect 272706 376896 272762 376952
rect 274086 374584 274142 374640
rect 273902 374040 273958 374096
rect 271878 336640 271934 336696
rect 272522 336640 272578 336696
rect 271878 335416 271934 335472
rect 271234 317600 271290 317656
rect 270314 184456 270370 184512
rect 272430 266328 272486 266384
rect 272430 262792 272486 262848
rect 274086 339496 274142 339552
rect 273994 306584 274050 306640
rect 272614 216552 272670 216608
rect 272614 215328 272670 215384
rect 274086 215328 274142 215384
rect 275282 303728 275338 303784
rect 274086 180104 274142 180160
rect 274638 178608 274694 178664
rect 272522 177520 272578 177576
rect 275282 178064 275338 178120
rect 278042 296792 278098 296848
rect 276754 295432 276810 295488
rect 277398 267008 277454 267064
rect 276754 210976 276810 211032
rect 276662 178744 276718 178800
rect 278134 295296 278190 295352
rect 278042 186360 278098 186416
rect 278134 185680 278190 185736
rect 274638 177248 274694 177304
rect 278318 189896 278374 189952
rect 278318 178608 278374 178664
rect 281354 376760 281410 376816
rect 280158 376624 280214 376680
rect 283562 359488 283618 359544
rect 280894 338680 280950 338736
rect 279514 298696 279570 298752
rect 279422 194520 279478 194576
rect 279974 178744 280030 178800
rect 279606 178064 279662 178120
rect 279422 175752 279478 175808
rect 279330 173712 279386 173768
rect 279422 172216 279478 172272
rect 280066 170992 280122 171048
rect 279330 170448 279386 170504
rect 265622 167184 265678 167240
rect 265622 164872 265678 164928
rect 265438 160248 265494 160304
rect 265162 159024 265218 159080
rect 265162 158888 265218 158944
rect 265070 158480 265126 158536
rect 264978 157664 265034 157720
rect 265070 157120 265126 157176
rect 264978 156712 265034 156768
rect 265162 156576 265218 156632
rect 265162 156304 265218 156360
rect 265070 155896 265126 155952
rect 264978 155488 265034 155544
rect 264978 154128 265034 154184
rect 264426 153448 264482 153504
rect 264242 135088 264298 135144
rect 264334 118088 264390 118144
rect 264242 111968 264298 112024
rect 262954 66952 263010 67008
rect 259550 19352 259606 19408
rect 260102 19352 260158 19408
rect 262218 19216 262274 19272
rect 262954 19216 263010 19272
rect 261758 10276 261760 10296
rect 261760 10276 261812 10296
rect 261812 10276 261814 10296
rect 261758 10240 261814 10276
rect 260102 3440 260158 3496
rect 260654 3440 260710 3496
rect 265162 153720 265218 153776
rect 265070 152904 265126 152960
rect 264978 152496 265034 152552
rect 265346 151544 265402 151600
rect 265070 150728 265126 150784
rect 264978 149912 265034 149968
rect 267278 159296 267334 159352
rect 265714 154536 265770 154592
rect 265806 151952 265862 152008
rect 265622 148960 265678 149016
rect 265162 148552 265218 148608
rect 265070 148280 265126 148336
rect 265070 148144 265126 148200
rect 264978 147756 265034 147792
rect 264978 147736 264980 147756
rect 264980 147736 265032 147756
rect 265032 147736 265034 147756
rect 265070 147328 265126 147384
rect 264978 146376 265034 146432
rect 265162 145968 265218 146024
rect 264978 145696 265034 145752
rect 265070 145560 265126 145616
rect 264978 145152 265034 145208
rect 264978 144744 265034 144800
rect 264610 143792 264666 143848
rect 264426 108568 264482 108624
rect 265254 144336 265310 144392
rect 265070 143384 265126 143440
rect 264978 142160 265034 142216
rect 265254 141208 265310 141264
rect 264978 139984 265034 140040
rect 265070 139168 265126 139224
rect 264978 138216 265034 138272
rect 264978 137808 265034 137864
rect 265070 136584 265126 136640
rect 264978 135632 265034 135688
rect 265070 135224 265126 135280
rect 265162 134816 265218 134872
rect 265070 134408 265126 134464
rect 264978 134000 265034 134056
rect 264978 133592 265034 133648
rect 264978 131824 265034 131880
rect 265714 142976 265770 143032
rect 265622 134136 265678 134192
rect 264978 131008 265034 131064
rect 265070 129240 265126 129296
rect 264978 128832 265034 128888
rect 264978 127880 265034 127936
rect 265070 127472 265126 127528
rect 264978 125840 265034 125896
rect 264978 124480 265034 124536
rect 265070 124072 265126 124128
rect 264978 122884 264980 122904
rect 264980 122884 265032 122904
rect 265032 122884 265034 122904
rect 264978 122848 265034 122884
rect 264978 121896 265034 121952
rect 264978 120672 265034 120728
rect 265070 120264 265126 120320
rect 264978 119312 265034 119368
rect 265070 118904 265126 118960
rect 264978 118496 265034 118552
rect 265162 116728 265218 116784
rect 264978 115948 264980 115968
rect 264980 115948 265032 115968
rect 265032 115948 265034 115968
rect 264978 115912 265034 115948
rect 265070 115096 265126 115152
rect 264978 114572 265034 114608
rect 264978 114552 264980 114572
rect 264980 114552 265032 114572
rect 265032 114552 265034 114572
rect 264978 114144 265034 114200
rect 264610 113736 264666 113792
rect 265162 113872 265218 113928
rect 264978 112512 265034 112568
rect 265070 111560 265126 111616
rect 264978 111152 265034 111208
rect 265070 110336 265126 110392
rect 264978 108976 265034 109032
rect 265254 106936 265310 106992
rect 264978 105984 265034 106040
rect 265162 105576 265218 105632
rect 265070 104760 265126 104816
rect 264978 104352 265034 104408
rect 264518 103808 264574 103864
rect 264978 103400 265034 103456
rect 265070 102584 265126 102640
rect 264978 101224 265034 101280
rect 264978 100000 265034 100056
rect 265162 100836 265218 100872
rect 265162 100816 265164 100836
rect 265164 100816 265216 100836
rect 265216 100816 265218 100836
rect 265070 98912 265126 98968
rect 264978 98640 265034 98696
rect 264978 97824 265034 97880
rect 264518 97416 264574 97472
rect 264518 80688 264574 80744
rect 265806 139576 265862 139632
rect 265714 98232 265770 98288
rect 265622 61376 265678 61432
rect 267094 131416 267150 131472
rect 265898 126248 265954 126304
rect 267002 121488 267058 121544
rect 265806 91704 265862 91760
rect 267186 125296 267242 125352
rect 279330 136856 279386 136912
rect 282182 326304 282238 326360
rect 282918 310392 282974 310448
rect 283562 310392 283618 310448
rect 280434 193976 280490 194032
rect 280158 118360 280214 118416
rect 267278 106392 267334 106448
rect 267186 83544 267242 83600
rect 279330 105712 279386 105768
rect 280434 174664 280490 174720
rect 280342 151816 280398 151872
rect 280342 145016 280398 145072
rect 280250 105440 280306 105496
rect 279422 104896 279478 104952
rect 267830 96600 267886 96656
rect 267738 95784 267794 95840
rect 267278 73752 267334 73808
rect 267094 68176 267150 68232
rect 273350 94424 273406 94480
rect 269118 29552 269174 29608
rect 268382 6840 268438 6896
rect 273166 66816 273222 66872
rect 276018 91840 276074 91896
rect 273902 37984 273958 38040
rect 273350 35128 273406 35184
rect 273902 12280 273958 12336
rect 274546 12280 274602 12336
rect 279422 99592 279478 99648
rect 279330 96600 279386 96656
rect 280158 98504 280214 98560
rect 280066 95784 280122 95840
rect 279330 94968 279386 95024
rect 280158 95104 280214 95160
rect 280066 93744 280122 93800
rect 281538 175480 281594 175536
rect 281538 168680 281594 168736
rect 281630 165552 281686 165608
rect 281630 162560 281686 162616
rect 282182 246200 282238 246256
rect 282182 237904 282238 237960
rect 281814 173984 281870 174040
rect 281906 169360 281962 169416
rect 281906 166368 281962 166424
rect 281906 161780 281908 161800
rect 281908 161780 281960 161800
rect 281960 161780 281962 161800
rect 281906 161744 281962 161780
rect 281814 158752 281870 158808
rect 282090 157936 282146 157992
rect 281722 157256 281778 157312
rect 281538 155624 281594 155680
rect 282090 154128 282146 154184
rect 282826 164872 282882 164928
rect 282826 164056 282882 164112
rect 282826 161064 282882 161120
rect 282826 160248 282882 160304
rect 282826 159432 282882 159488
rect 282274 154944 282330 155000
rect 282826 153448 282882 153504
rect 282182 152632 282238 152688
rect 281906 151136 281962 151192
rect 282182 148008 282238 148064
rect 281722 147328 281778 147384
rect 280802 143520 280858 143576
rect 282826 150340 282882 150376
rect 282826 150320 282828 150340
rect 282828 150320 282880 150340
rect 282880 150320 282882 150340
rect 282734 149640 282790 149696
rect 282826 148824 282882 148880
rect 282826 146512 282882 146568
rect 282826 145832 282882 145888
rect 282826 144200 282882 144256
rect 285586 359488 285642 359544
rect 285586 349832 285642 349888
rect 284942 321544 284998 321600
rect 289634 375264 289690 375320
rect 287978 374584 288034 374640
rect 286230 344292 286232 344312
rect 286232 344292 286284 344312
rect 286284 344292 286286 344312
rect 286230 344256 286286 344292
rect 287702 341536 287758 341592
rect 287058 314880 287114 314936
rect 285678 309848 285734 309904
rect 284298 193024 284354 193080
rect 284298 177964 284300 177984
rect 284300 177964 284352 177984
rect 284352 177964 284354 177984
rect 284298 177928 284354 177964
rect 283102 142704 283158 142760
rect 281906 141208 281962 141264
rect 281630 137400 281686 137456
rect 281722 132096 281778 132152
rect 282090 128968 282146 129024
rect 280894 128288 280950 128344
rect 282826 142060 282828 142080
rect 282828 142060 282880 142080
rect 282880 142060 282882 142080
rect 282826 142024 282882 142060
rect 282826 140392 282882 140448
rect 282734 139712 282790 139768
rect 282826 138896 282882 138952
rect 282826 138216 282882 138272
rect 282274 135904 282330 135960
rect 282826 132776 282882 132832
rect 282642 131280 282698 131336
rect 282274 130600 282330 130656
rect 282734 130328 282790 130384
rect 282182 127472 282238 127528
rect 281722 126792 281778 126848
rect 280434 121352 280490 121408
rect 281538 110744 281594 110800
rect 281538 103944 281594 104000
rect 281630 103128 281686 103184
rect 280526 100816 280582 100872
rect 282274 125976 282330 126032
rect 282274 124752 282330 124808
rect 281998 123664 282054 123720
rect 282826 129784 282882 129840
rect 282734 125160 282790 125216
rect 282366 124480 282422 124536
rect 282826 122984 282882 123040
rect 282826 122168 282882 122224
rect 282826 120672 282882 120728
rect 282826 119856 282882 119912
rect 282734 119176 282790 119232
rect 282550 117544 282606 117600
rect 282274 116864 282330 116920
rect 282182 115368 282238 115424
rect 281814 113076 281870 113112
rect 281814 113056 281816 113076
rect 281816 113056 281868 113076
rect 281868 113056 281870 113076
rect 282826 116084 282828 116104
rect 282828 116084 282880 116104
rect 282880 116084 282882 116104
rect 282826 116048 282882 116084
rect 282458 114552 282514 114608
rect 282826 113736 282882 113792
rect 282826 112240 282882 112296
rect 282826 111580 282882 111616
rect 282826 111560 282828 111580
rect 282828 111560 282880 111580
rect 282880 111560 282882 111580
rect 282826 109248 282882 109304
rect 282274 108432 282330 108488
rect 282366 107752 282422 107808
rect 282826 106936 282882 106992
rect 285770 228248 285826 228304
rect 284942 224848 284998 224904
rect 284666 177384 284722 177440
rect 281998 97824 282054 97880
rect 279054 84088 279110 84144
rect 278042 82048 278098 82104
rect 276110 3460 276166 3496
rect 280802 77832 280858 77888
rect 276110 3440 276112 3460
rect 276112 3440 276164 3460
rect 276164 3440 276166 3460
rect 283562 64232 283618 64288
rect 282182 55800 282238 55856
rect 280894 26832 280950 26888
rect 280802 3848 280858 3904
rect 284942 24792 284998 24848
rect 284298 23432 284354 23488
rect 284942 23432 284998 23488
rect 282274 3984 282330 4040
rect 287334 177520 287390 177576
rect 289910 251912 289966 251968
rect 291106 251932 291162 251968
rect 291106 251912 291108 251932
rect 291108 251912 291160 251932
rect 291160 251912 291162 251932
rect 291474 178608 291530 178664
rect 292670 196696 292726 196752
rect 292578 100816 292634 100872
rect 291198 97824 291254 97880
rect 289818 93064 289874 93120
rect 286322 91704 286378 91760
rect 288346 12144 288402 12200
rect 288990 8200 289046 8256
rect 287794 3440 287850 3496
rect 288346 3440 288402 3496
rect 292486 66136 292542 66192
rect 293222 184184 293278 184240
rect 293222 101360 293278 101416
rect 293222 100816 293278 100872
rect 295338 229764 295394 229800
rect 295338 229744 295340 229764
rect 295340 229744 295392 229764
rect 295392 229744 295394 229764
rect 295338 185544 295394 185600
rect 295338 149096 295394 149152
rect 295522 289992 295578 290048
rect 295890 289992 295946 290048
rect 297454 289856 297510 289912
rect 297454 283464 297510 283520
rect 298006 246336 298062 246392
rect 298006 245656 298062 245712
rect 295982 224304 296038 224360
rect 296718 222944 296774 223000
rect 297914 222944 297970 223000
rect 299478 324944 299534 325000
rect 298834 251776 298890 251832
rect 298466 225528 298522 225584
rect 298742 218728 298798 218784
rect 298006 96464 298062 96520
rect 292578 7520 292634 7576
rect 292578 3712 292634 3768
rect 299662 86284 299718 86320
rect 299662 86264 299664 86284
rect 299664 86264 299716 86284
rect 299716 86264 299718 86284
rect 301502 212064 301558 212120
rect 301042 188400 301098 188456
rect 301042 125432 301098 125488
rect 301318 125432 301374 125488
rect 301318 124752 301374 124808
rect 300766 11736 300822 11792
rect 300674 7520 300730 7576
rect 299662 3984 299718 4040
rect 300674 3984 300730 4040
rect 307022 366288 307078 366344
rect 304998 342896 305054 342952
rect 304998 342216 305054 342272
rect 305642 342216 305698 342272
rect 303618 293800 303674 293856
rect 303618 292576 303674 292632
rect 304262 292576 304318 292632
rect 304998 291216 305054 291272
rect 305090 238720 305146 238776
rect 302974 30912 303030 30968
rect 308402 363568 308458 363624
rect 309782 341400 309838 341456
rect 309782 340856 309838 340912
rect 309138 304952 309194 305008
rect 308402 280744 308458 280800
rect 307758 250008 307814 250064
rect 310426 304952 310482 305008
rect 309874 199280 309930 199336
rect 309782 119312 309838 119368
rect 309138 84768 309194 84824
rect 308402 54440 308458 54496
rect 308402 3984 308458 4040
rect 309046 3984 309102 4040
rect 311898 340856 311954 340912
rect 310518 60560 310574 60616
rect 311162 60560 311218 60616
rect 319626 376624 319682 376680
rect 313278 130328 313334 130384
rect 315302 193840 315358 193896
rect 313922 34448 313978 34504
rect 314566 34448 314622 34504
rect 316130 230288 316186 230344
rect 316682 230288 316738 230344
rect 316774 200776 316830 200832
rect 316682 189760 316738 189816
rect 319442 243480 319498 243536
rect 320270 349016 320326 349072
rect 320822 349016 320878 349072
rect 320822 347792 320878 347848
rect 320178 221856 320234 221912
rect 320638 221856 320694 221912
rect 322202 298152 322258 298208
rect 320914 204992 320970 205048
rect 324318 345616 324374 345672
rect 324962 308352 325018 308408
rect 323674 277480 323730 277536
rect 322294 239400 322350 239456
rect 322294 237360 322350 237416
rect 323582 224168 323638 224224
rect 316682 14456 316738 14512
rect 324318 234540 324320 234560
rect 324320 234540 324372 234560
rect 324372 234540 324374 234560
rect 324318 234504 324374 234540
rect 331862 354592 331918 354648
rect 328458 351872 328514 351928
rect 329102 351872 329158 351928
rect 326342 337320 326398 337376
rect 327722 337320 327778 337376
rect 324962 108296 325018 108352
rect 327078 135904 327134 135960
rect 328366 135924 328422 135960
rect 328366 135904 328368 135924
rect 328368 135904 328420 135924
rect 328420 135904 328422 135924
rect 326342 88984 326398 89040
rect 322294 3712 322350 3768
rect 325054 37848 325110 37904
rect 324410 26152 324466 26208
rect 324962 26152 325018 26208
rect 329102 68176 329158 68232
rect 332598 288396 332600 288416
rect 332600 288396 332652 288416
rect 332652 288396 332654 288416
rect 332598 288360 332654 288396
rect 332598 284300 332654 284336
rect 332598 284280 332600 284300
rect 332600 284280 332652 284300
rect 332652 284280 332654 284300
rect 339498 375264 339554 375320
rect 337382 357992 337438 358048
rect 336002 354728 336058 354784
rect 334806 283464 334862 283520
rect 334714 184320 334770 184376
rect 338762 285640 338818 285696
rect 340142 329840 340198 329896
rect 338854 215872 338910 215928
rect 341522 362208 341578 362264
rect 340878 317328 340934 317384
rect 340234 126248 340290 126304
rect 344006 376896 344062 376952
rect 342902 375264 342958 375320
rect 342902 374720 342958 374776
rect 342994 239400 343050 239456
rect 342902 237224 342958 237280
rect 341614 234640 341670 234696
rect 342994 139984 343050 140040
rect 348422 376488 348478 376544
rect 352562 377440 352618 377496
rect 351090 374584 351146 374640
rect 345754 211928 345810 211984
rect 351182 356632 351238 356688
rect 350446 346432 350502 346488
rect 353942 375944 353998 376000
rect 349802 142160 349858 142216
rect 342166 3304 342222 3360
rect 352562 306448 352618 306504
rect 351182 195200 351238 195256
rect 354034 374040 354090 374096
rect 352654 232464 352710 232520
rect 352746 124072 352802 124128
rect 352562 90344 352618 90400
rect 351642 3848 351698 3904
rect 350446 3440 350502 3496
rect 354678 375672 354734 375728
rect 354678 367648 354734 367704
rect 354034 246336 354090 246392
rect 356242 423680 356298 423736
rect 356150 377440 356206 377496
rect 356334 394440 356390 394496
rect 356426 387096 356482 387152
rect 356426 373360 356482 373416
rect 358726 455912 358782 455968
rect 358726 453464 358782 453520
rect 358726 451016 358782 451072
rect 358726 448588 358782 448624
rect 358726 448568 358728 448588
rect 358728 448568 358780 448588
rect 358780 448568 358782 448588
rect 358726 446120 358782 446176
rect 358726 443672 358782 443728
rect 358726 438932 358782 438968
rect 358726 438912 358728 438932
rect 358728 438912 358780 438932
rect 358780 438912 358782 438932
rect 358726 436328 358782 436384
rect 358726 433880 358782 433936
rect 358726 428984 358782 429040
rect 358726 426536 358782 426592
rect 357530 421640 357586 421696
rect 357438 371864 357494 371920
rect 356794 370504 356850 370560
rect 358726 419192 358782 419248
rect 358726 416780 358728 416800
rect 358728 416780 358780 416800
rect 358780 416780 358782 416800
rect 358726 416744 358782 416780
rect 358726 414296 358782 414352
rect 358726 411848 358782 411904
rect 358726 406952 358782 407008
rect 358726 404232 358782 404288
rect 358726 401784 358782 401840
rect 358634 399336 358690 399392
rect 357622 391992 357678 392048
rect 357714 389544 357770 389600
rect 357898 384648 357954 384704
rect 357898 379752 357954 379808
rect 358082 371320 358138 371376
rect 357530 357992 357586 358048
rect 354034 124072 354090 124128
rect 359094 441224 359150 441280
rect 359002 431432 359058 431488
rect 358082 137672 358138 137728
rect 352562 3440 352618 3496
rect 359462 289040 359518 289096
rect 360842 543768 360898 543824
rect 360934 143520 360990 143576
rect 362958 538464 363014 538520
rect 361854 375944 361910 376000
rect 364430 370504 364486 370560
rect 365718 291760 365774 291816
rect 366362 282104 366418 282160
rect 361578 119992 361634 120048
rect 361578 119312 361634 119368
rect 371330 362344 371386 362400
rect 371330 323584 371386 323640
rect 370502 280744 370558 280800
rect 369122 200640 369178 200696
rect 372710 329024 372766 329080
rect 374642 373360 374698 373416
rect 373262 231104 373318 231160
rect 371882 166232 371938 166288
rect 371238 126248 371294 126304
rect 370502 103128 370558 103184
rect 374734 190440 374790 190496
rect 376758 369008 376814 369064
rect 376022 99320 376078 99376
rect 376114 12280 376170 12336
rect 378138 193160 378194 193216
rect 378874 193160 378930 193216
rect 378874 132368 378930 132424
rect 388442 541048 388498 541104
rect 381542 374720 381598 374776
rect 380162 104080 380218 104136
rect 381634 102720 381690 102776
rect 381542 97688 381598 97744
rect 378874 93744 378930 93800
rect 377402 9560 377458 9616
rect 387062 312432 387118 312488
rect 383014 138624 383070 138680
rect 389178 535472 389234 535528
rect 388442 148280 388498 148336
rect 389178 140664 389234 140720
rect 389178 139984 389234 140040
rect 392674 192480 392730 192536
rect 390558 132368 390614 132424
rect 390558 131144 390614 131200
rect 389914 129920 389970 129976
rect 388442 40568 388498 40624
rect 393410 182960 393466 183016
rect 395342 142704 395398 142760
rect 393410 138760 393466 138816
rect 393410 131280 393466 131336
rect 394606 128696 394662 128752
rect 397366 266328 397422 266384
rect 396814 262792 396870 262848
rect 397366 262792 397422 262848
rect 396722 210296 396778 210352
rect 395986 146240 396042 146296
rect 397458 226888 397514 226944
rect 396814 125976 396870 126032
rect 397550 137536 397606 137592
rect 397550 136720 397606 136776
rect 397642 135496 397698 135552
rect 398654 134816 398710 134872
rect 397550 134000 397606 134056
rect 397642 133456 397698 133512
rect 397550 132096 397606 132152
rect 397550 130600 397606 130656
rect 397550 129240 397606 129296
rect 397550 127880 397606 127936
rect 398102 126656 398158 126712
rect 397550 125160 397606 125216
rect 400218 214648 400274 214704
rect 399574 146240 399630 146296
rect 399482 142296 399538 142352
rect 398838 126656 398894 126712
rect 398746 124616 398802 124672
rect 397550 123800 397606 123856
rect 397642 123256 397698 123312
rect 397550 122440 397606 122496
rect 397734 121080 397790 121136
rect 397642 120536 397698 120592
rect 397734 119992 397790 120048
rect 397642 119856 397698 119912
rect 397550 119176 397606 119232
rect 397642 118360 397698 118416
rect 397550 117816 397606 117872
rect 397550 117136 397606 117192
rect 397550 115776 397606 115832
rect 397642 115096 397698 115152
rect 397550 114452 397552 114472
rect 397552 114452 397604 114472
rect 397604 114452 397606 114472
rect 397550 114416 397606 114452
rect 397642 113736 397698 113792
rect 398746 112920 398802 112976
rect 397550 112376 397606 112432
rect 397458 111732 397460 111752
rect 397460 111732 397512 111752
rect 397512 111732 397514 111752
rect 397458 111696 397514 111732
rect 397550 110200 397606 110256
rect 397458 108996 397514 109032
rect 397458 108976 397460 108996
rect 397460 108976 397512 108996
rect 397512 108976 397514 108996
rect 398194 111016 398250 111072
rect 397642 108316 397698 108352
rect 397642 108296 397644 108316
rect 397644 108296 397696 108316
rect 397696 108296 397698 108316
rect 397458 107480 397514 107536
rect 397550 106800 397606 106856
rect 397458 106120 397514 106176
rect 397458 104796 397460 104816
rect 397460 104796 397512 104816
rect 397512 104796 397514 104816
rect 397458 104760 397514 104796
rect 397550 104216 397606 104272
rect 397458 103436 397460 103456
rect 397460 103436 397512 103456
rect 397512 103436 397514 103456
rect 397458 103400 397514 103436
rect 397458 100816 397514 100872
rect 398654 104080 398710 104136
rect 398194 102040 398250 102096
rect 397918 96328 397974 96384
rect 396906 95104 396962 95160
rect 403622 316104 403678 316160
rect 400310 181328 400366 181384
rect 405002 202136 405058 202192
rect 582654 697176 582710 697232
rect 582562 683848 582618 683904
rect 582470 644000 582526 644056
rect 582378 564304 582434 564360
rect 580262 538192 580318 538248
rect 580170 537784 580226 537840
rect 407854 374584 407910 374640
rect 406014 146920 406070 146976
rect 405738 142296 405794 142352
rect 409878 247560 409934 247616
rect 408590 218592 408646 218648
rect 407946 139984 408002 140040
rect 412546 376760 412602 376816
rect 411258 203632 411314 203688
rect 410522 159296 410578 159352
rect 412638 142704 412694 142760
rect 415398 143384 415454 143440
rect 416134 143384 416190 143440
rect 415490 142704 415546 142760
rect 416134 142160 416190 142216
rect 420182 214512 420238 214568
rect 418894 204856 418950 204912
rect 423678 208392 423734 208448
rect 422942 206216 422998 206272
rect 427818 317464 427874 317520
rect 426438 203496 426494 203552
rect 425150 149096 425206 149152
rect 425058 143384 425114 143440
rect 425794 143384 425850 143440
rect 419630 139440 419686 139496
rect 425518 139440 425574 139496
rect 432602 314744 432658 314800
rect 427082 142160 427138 142216
rect 429198 197920 429254 197976
rect 427450 139440 427506 139496
rect 431314 139440 431370 139496
rect 433522 143520 433578 143576
rect 432602 140800 432658 140856
rect 439134 211792 439190 211848
rect 436374 139440 436430 139496
rect 438858 139304 438914 139360
rect 399850 137672 399906 137728
rect 440238 207032 440294 207088
rect 439594 138488 439650 138544
rect 439502 135768 439558 135824
rect 440238 132776 440294 132832
rect 439410 131688 439466 131744
rect 440238 127880 440294 127936
rect 439410 120808 439466 120864
rect 439410 115912 439466 115968
rect 439318 111832 439374 111888
rect 439318 104352 439374 104408
rect 439410 103808 439466 103864
rect 400034 97824 400090 97880
rect 400862 96872 400918 96928
rect 404542 99320 404598 99376
rect 402610 96872 402666 96928
rect 405738 96328 405794 96384
rect 406474 96328 406530 96384
rect 409694 93744 409750 93800
rect 408498 92520 408554 92576
rect 409694 92520 409750 92576
rect 410982 89664 411038 89720
rect 413558 99864 413614 99920
rect 412270 93064 412326 93120
rect 414846 99864 414902 99920
rect 414662 97144 414718 97200
rect 418710 96464 418766 96520
rect 418066 91704 418122 91760
rect 419998 99048 420054 99104
rect 421930 99184 421986 99240
rect 421286 91024 421342 91080
rect 423862 97144 423918 97200
rect 425702 97008 425758 97064
rect 427726 97008 427782 97064
rect 427082 96872 427138 96928
rect 427910 96872 427966 96928
rect 431590 97688 431646 97744
rect 433522 99864 433578 99920
rect 434810 99864 434866 99920
rect 434810 97824 434866 97880
rect 437386 97824 437442 97880
rect 439318 101632 439374 101688
rect 438674 95104 438730 95160
rect 439502 102312 439558 102368
rect 440422 137400 440478 137456
rect 440330 121896 440386 121952
rect 440422 119040 440478 119096
rect 440330 114960 440386 115016
rect 441710 179968 441766 180024
rect 441710 136176 441766 136232
rect 441894 138896 441950 138952
rect 441986 138080 442042 138136
rect 442906 136740 442962 136776
rect 442906 136720 442908 136740
rect 442908 136720 442960 136740
rect 442960 136720 442962 136740
rect 442906 134816 442962 134872
rect 442906 133456 442962 133512
rect 441802 132096 441858 132152
rect 442906 130772 442908 130792
rect 442908 130772 442960 130792
rect 442960 130772 442962 130792
rect 442906 130736 442962 130772
rect 442906 129920 442962 129976
rect 442170 129240 442226 129296
rect 442906 127220 442962 127256
rect 442906 127200 442908 127220
rect 442908 127200 442960 127220
rect 442960 127200 442962 127220
rect 442906 126656 442962 126712
rect 442814 125976 442870 126032
rect 442906 124616 442962 124672
rect 441618 123936 441674 123992
rect 442630 123936 442686 123992
rect 441894 122612 441896 122632
rect 441896 122612 441948 122632
rect 441948 122612 441950 122632
rect 441894 122576 441950 122612
rect 441618 120400 441674 120456
rect 440882 114416 440938 114472
rect 442906 118532 442908 118552
rect 442908 118532 442960 118552
rect 442960 118532 442962 118552
rect 442906 118496 442962 118532
rect 442906 117136 442962 117192
rect 444378 220088 444434 220144
rect 443090 188264 443146 188320
rect 443182 148280 443238 148336
rect 443090 125160 443146 125216
rect 442906 116340 442962 116376
rect 442906 116320 442908 116340
rect 442908 116320 442960 116340
rect 442960 116320 442962 116340
rect 442906 115812 442908 115832
rect 442908 115812 442960 115832
rect 442960 115812 442962 115832
rect 442906 115776 442962 115812
rect 442906 113600 442962 113656
rect 442906 113092 442908 113112
rect 442908 113092 442960 113112
rect 442960 113092 442962 113112
rect 442906 113056 442962 113092
rect 442170 109520 442226 109576
rect 442446 108996 442502 109032
rect 442446 108976 442448 108996
rect 442448 108976 442500 108996
rect 442500 108976 442502 108996
rect 441710 108160 441766 108216
rect 441618 84768 441674 84824
rect 442906 107480 442962 107536
rect 442354 106120 442410 106176
rect 442722 105576 442778 105632
rect 442170 100816 442226 100872
rect 442906 100136 442962 100192
rect 443182 103400 443238 103456
rect 443090 71712 443146 71768
rect 580354 524456 580410 524512
rect 582378 511264 582434 511320
rect 580262 484608 580318 484664
rect 582378 431568 582434 431624
rect 582378 365064 582434 365120
rect 582378 335960 582434 336016
rect 582378 333240 582434 333296
rect 445942 182824 445998 182880
rect 445850 177248 445906 177304
rect 382922 3984 382978 4040
rect 358082 3304 358138 3360
rect 446034 109792 446090 109848
rect 449162 246200 449218 246256
rect 447230 119312 447286 119368
rect 449990 189624 450046 189680
rect 448610 97824 448666 97880
rect 449990 109792 450046 109848
rect 580906 165824 580962 165880
rect 580170 139304 580226 139360
rect 580262 125976 580318 126032
rect 580170 99456 580226 99512
rect 582562 458088 582618 458144
rect 583206 670656 583262 670712
rect 582746 630808 582802 630864
rect 582930 617480 582986 617536
rect 582838 577632 582894 577688
rect 582746 553968 582802 554024
rect 582654 404912 582710 404968
rect 583022 590960 583078 591016
rect 583114 559000 583170 559056
rect 583022 471416 583078 471472
rect 582930 404912 582986 404968
rect 582838 376624 582894 376680
rect 583114 458088 583170 458144
rect 583298 418240 583354 418296
rect 583206 377304 583262 377360
rect 583022 364248 583078 364304
rect 582838 351872 582894 351928
rect 583022 325216 583078 325272
rect 582838 310936 582894 310992
rect 582746 298696 582802 298752
rect 582930 298696 582986 298752
rect 582746 272176 582802 272232
rect 582838 258848 582894 258904
rect 583298 312024 583354 312080
rect 583114 310936 583170 310992
rect 583114 310528 583170 310584
rect 583022 247560 583078 247616
rect 583022 245520 583078 245576
rect 582654 146920 582710 146976
rect 582470 97144 582526 97200
rect 582470 72936 582526 72992
rect 583206 266328 583262 266384
rect 583206 232328 583262 232384
rect 583574 222808 583630 222864
rect 583298 219000 583354 219056
rect 583206 192480 583262 192536
rect 583022 112784 583078 112840
rect 583390 205672 583446 205728
rect 583482 178608 583538 178664
rect 582746 86128 582802 86184
rect 582654 59608 582710 59664
rect 583114 93064 583170 93120
rect 583022 46280 583078 46336
rect 582838 33088 582894 33144
rect 582562 19760 582618 19816
rect 583114 6568 583170 6624
rect 583758 196560 583814 196616
rect 583666 152224 583722 152280
rect 583666 99048 583722 99104
<< metal3 >>
rect 69606 702476 69612 702540
rect 69676 702538 69682 702540
rect 154113 702538 154179 702541
rect 69676 702536 154179 702538
rect 69676 702480 154118 702536
rect 154174 702480 154179 702536
rect 69676 702478 154179 702480
rect 69676 702476 69682 702478
rect 154113 702475 154179 702478
rect -960 697220 480 697460
rect 582649 697234 582715 697237
rect 583520 697234 584960 697324
rect 582649 697232 584960 697234
rect 582649 697176 582654 697232
rect 582710 697176 584960 697232
rect 582649 697174 584960 697176
rect 582649 697171 582715 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 582557 683906 582623 683909
rect 583520 683906 584960 683996
rect 582557 683904 584960 683906
rect 582557 683848 582562 683904
rect 582618 683848 584960 683904
rect 582557 683846 584960 683848
rect 582557 683843 582623 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 583201 670714 583267 670717
rect 583520 670714 584960 670804
rect 583201 670712 584960 670714
rect 583201 670656 583206 670712
rect 583262 670656 584960 670712
rect 583201 670654 584960 670656
rect 583201 670651 583267 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 2773 658202 2839 658205
rect -960 658200 2839 658202
rect -960 658144 2778 658200
rect 2834 658144 2839 658200
rect -960 658142 2839 658144
rect -960 658052 480 658142
rect 2773 658139 2839 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 582465 644058 582531 644061
rect 583520 644058 584960 644148
rect 582465 644056 584960 644058
rect 582465 644000 582470 644056
rect 582526 644000 584960 644056
rect 582465 643998 584960 644000
rect 582465 643995 582531 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 582741 630866 582807 630869
rect 583520 630866 584960 630956
rect 582741 630864 584960 630866
rect 582741 630808 582746 630864
rect 582802 630808 584960 630864
rect 582741 630806 584960 630808
rect 582741 630803 582807 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 582925 617538 582991 617541
rect 583520 617538 584960 617628
rect 582925 617536 584960 617538
rect 582925 617480 582930 617536
rect 582986 617480 584960 617536
rect 582925 617478 584960 617480
rect 582925 617475 582991 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect 76741 593466 76807 593469
rect 100753 593466 100819 593469
rect 76741 593464 100819 593466
rect 76741 593408 76746 593464
rect 76802 593408 100758 593464
rect 100814 593408 100819 593464
rect 76741 593406 100819 593408
rect 76741 593403 76807 593406
rect 100753 593403 100819 593406
rect -960 592908 480 593148
rect 73981 592106 74047 592109
rect 95877 592106 95943 592109
rect 73981 592104 95943 592106
rect 73981 592048 73986 592104
rect 74042 592048 95882 592104
rect 95938 592048 95943 592104
rect 73981 592046 95943 592048
rect 73981 592043 74047 592046
rect 95877 592043 95943 592046
rect 82261 591018 82327 591021
rect 104157 591018 104223 591021
rect 82261 591016 104223 591018
rect 82261 590960 82266 591016
rect 82322 590960 104162 591016
rect 104218 590960 104223 591016
rect 82261 590958 104223 590960
rect 82261 590955 82327 590958
rect 104157 590955 104223 590958
rect 583017 591018 583083 591021
rect 583520 591018 584960 591108
rect 583017 591016 584960 591018
rect 583017 590960 583022 591016
rect 583078 590960 584960 591016
rect 583017 590958 584960 590960
rect 583017 590955 583083 590958
rect 86861 590882 86927 590885
rect 97257 590882 97323 590885
rect 86861 590880 97323 590882
rect 86861 590824 86866 590880
rect 86922 590824 97262 590880
rect 97318 590824 97323 590880
rect 583520 590868 584960 590958
rect 86861 590822 97323 590824
rect 86861 590819 86927 590822
rect 97257 590819 97323 590822
rect 65977 590746 66043 590749
rect 70301 590746 70367 590749
rect 71129 590746 71195 590749
rect 65977 590744 71195 590746
rect 65977 590688 65982 590744
rect 66038 590688 70306 590744
rect 70362 590688 71134 590744
rect 71190 590688 71195 590744
rect 65977 590686 71195 590688
rect 65977 590683 66043 590686
rect 70301 590683 70367 590686
rect 71129 590683 71195 590686
rect 73061 590746 73127 590749
rect 81893 590746 81959 590749
rect 73061 590744 81959 590746
rect 73061 590688 73066 590744
rect 73122 590688 81898 590744
rect 81954 590688 81959 590744
rect 73061 590686 81959 590688
rect 73061 590683 73127 590686
rect 81893 590683 81959 590686
rect 74441 589930 74507 589933
rect 90357 589930 90423 589933
rect 74441 589928 90423 589930
rect 74441 589872 74446 589928
rect 74502 589872 90362 589928
rect 90418 589872 90423 589928
rect 74441 589870 90423 589872
rect 74441 589867 74507 589870
rect 90357 589867 90423 589870
rect 81341 589522 81407 589525
rect 100661 589522 100727 589525
rect 81341 589520 103530 589522
rect 81341 589464 81346 589520
rect 81402 589464 100666 589520
rect 100722 589464 103530 589520
rect 81341 589462 103530 589464
rect 81341 589459 81407 589462
rect 100661 589459 100727 589462
rect 77661 589386 77727 589389
rect 98637 589386 98703 589389
rect 77661 589384 98703 589386
rect 77661 589328 77666 589384
rect 77722 589328 98642 589384
rect 98698 589328 98703 589384
rect 77661 589326 98703 589328
rect 103470 589386 103530 589462
rect 255957 589386 256023 589389
rect 103470 589384 256023 589386
rect 103470 589328 255962 589384
rect 256018 589328 256023 589384
rect 103470 589326 256023 589328
rect 77661 589323 77727 589326
rect 98637 589323 98703 589326
rect 255957 589323 256023 589326
rect 79685 588706 79751 588709
rect 105537 588706 105603 588709
rect 79685 588704 105603 588706
rect 79685 588648 79690 588704
rect 79746 588648 105542 588704
rect 105598 588648 105603 588704
rect 79685 588646 105603 588648
rect 79685 588643 79751 588646
rect 105537 588643 105603 588646
rect 88057 588570 88123 588573
rect 88190 588570 88196 588572
rect 88057 588568 88196 588570
rect 88057 588512 88062 588568
rect 88118 588512 88196 588568
rect 88057 588510 88196 588512
rect 88057 588507 88123 588510
rect 88190 588508 88196 588510
rect 88260 588508 88266 588572
rect 66805 588434 66871 588437
rect 66805 588432 68908 588434
rect 66805 588376 66810 588432
rect 66866 588376 68908 588432
rect 66805 588374 68908 588376
rect 66805 588371 66871 588374
rect 91093 587618 91159 587621
rect 88596 587616 91159 587618
rect 88596 587560 91098 587616
rect 91154 587560 91159 587616
rect 88596 587558 91159 587560
rect 91093 587555 91159 587558
rect 66253 586530 66319 586533
rect 66253 586528 66362 586530
rect 66253 586472 66258 586528
rect 66314 586472 66362 586528
rect 66253 586467 66362 586472
rect 66302 586394 66362 586467
rect 68878 586394 68938 587044
rect 66302 586334 68938 586394
rect 89713 586258 89779 586261
rect 88596 586256 89779 586258
rect 88596 586200 89718 586256
rect 89774 586200 89779 586256
rect 88596 586198 89779 586200
rect 89713 586195 89779 586198
rect 66897 585714 66963 585717
rect 66897 585712 68908 585714
rect 66897 585656 66902 585712
rect 66958 585656 68908 585712
rect 66897 585654 68908 585656
rect 66897 585651 66963 585654
rect 88190 585652 88196 585716
rect 88260 585714 88266 585716
rect 118693 585714 118759 585717
rect 88260 585712 118759 585714
rect 88260 585656 118698 585712
rect 118754 585656 118759 585712
rect 88260 585654 118759 585656
rect 88260 585652 88266 585654
rect 118693 585651 118759 585654
rect 91277 584898 91343 584901
rect 88596 584896 91343 584898
rect 88596 584840 91282 584896
rect 91338 584840 91343 584896
rect 88596 584838 91343 584840
rect 91277 584835 91343 584838
rect 67725 584354 67791 584357
rect 67725 584352 68908 584354
rect 67725 584296 67730 584352
rect 67786 584296 68908 584352
rect 67725 584294 68908 584296
rect 67725 584291 67791 584294
rect 91829 583674 91895 583677
rect 88596 583672 91895 583674
rect 88596 583616 91834 583672
rect 91890 583616 91895 583672
rect 88596 583614 91895 583616
rect 91829 583611 91895 583614
rect 66805 582994 66871 582997
rect 66805 582992 68908 582994
rect 66805 582936 66810 582992
rect 66866 582936 68908 582992
rect 66805 582934 68908 582936
rect 66805 582931 66871 582934
rect 69422 582252 69428 582316
rect 69492 582252 69498 582316
rect 66529 581770 66595 581773
rect 69430 581770 69490 582252
rect 91277 582178 91343 582181
rect 88596 582176 91343 582178
rect 88596 582120 91282 582176
rect 91338 582120 91343 582176
rect 88596 582118 91343 582120
rect 91277 582115 91343 582118
rect 66529 581768 69490 581770
rect 66529 581712 66534 581768
rect 66590 581740 69490 581768
rect 66590 581712 69460 581740
rect 66529 581710 69460 581712
rect 66529 581707 66595 581710
rect 66805 580274 66871 580277
rect 66805 580272 68908 580274
rect 66805 580216 66810 580272
rect 66866 580216 68908 580272
rect 66805 580214 68908 580216
rect 66805 580211 66871 580214
rect -960 580002 480 580092
rect 3049 580002 3115 580005
rect -960 580000 3115 580002
rect -960 579944 3054 580000
rect 3110 579944 3115 580000
rect -960 579942 3115 579944
rect -960 579852 480 579942
rect 3049 579939 3115 579942
rect 88566 579730 88626 580788
rect 119470 579730 119476 579732
rect 88566 579670 119476 579730
rect 119470 579668 119476 579670
rect 119540 579668 119546 579732
rect 67766 578852 67772 578916
rect 67836 578914 67842 578916
rect 67836 578854 68908 578914
rect 67836 578852 67842 578854
rect 88566 578370 88626 579428
rect 120022 578370 120028 578372
rect 88566 578310 120028 578370
rect 120022 578308 120028 578310
rect 120092 578308 120098 578372
rect 91277 578098 91343 578101
rect 88596 578096 91343 578098
rect 88596 578040 91282 578096
rect 91338 578040 91343 578096
rect 88596 578038 91343 578040
rect 91277 578035 91343 578038
rect 582833 577690 582899 577693
rect 583520 577690 584960 577780
rect 582833 577688 584960 577690
rect 582833 577632 582838 577688
rect 582894 577632 584960 577688
rect 582833 577630 584960 577632
rect 582833 577627 582899 577630
rect 67817 577554 67883 577557
rect 67817 577552 68908 577554
rect 67817 577496 67822 577552
rect 67878 577496 68908 577552
rect 583520 577540 584960 577630
rect 67817 577494 68908 577496
rect 67817 577491 67883 577494
rect 91185 576738 91251 576741
rect 88596 576736 91251 576738
rect 88596 576680 91190 576736
rect 91246 576680 91251 576736
rect 88596 576678 91251 576680
rect 91185 576675 91251 576678
rect 66805 576194 66871 576197
rect 66805 576192 68908 576194
rect 66805 576136 66810 576192
rect 66866 576136 68908 576192
rect 66805 576134 68908 576136
rect 66805 576131 66871 576134
rect 91737 575378 91803 575381
rect 88596 575376 91803 575378
rect 88596 575320 91742 575376
rect 91798 575320 91803 575376
rect 88596 575318 91803 575320
rect 91737 575315 91803 575318
rect 67357 574970 67423 574973
rect 67357 574968 68908 574970
rect 67357 574912 67362 574968
rect 67418 574912 68908 574968
rect 67357 574910 68908 574912
rect 67357 574907 67423 574910
rect 91737 574018 91803 574021
rect 88596 574016 91803 574018
rect 88596 573960 91742 574016
rect 91798 573960 91803 574016
rect 88596 573958 91803 573960
rect 91737 573955 91803 573958
rect 65885 573474 65951 573477
rect 65885 573472 68908 573474
rect 65885 573416 65890 573472
rect 65946 573416 68908 573472
rect 65885 573414 68908 573416
rect 65885 573411 65951 573414
rect 91737 572658 91803 572661
rect 88596 572656 91803 572658
rect 88596 572600 91742 572656
rect 91798 572600 91803 572656
rect 88596 572598 91803 572600
rect 91737 572595 91803 572598
rect 66805 572114 66871 572117
rect 66805 572112 68908 572114
rect 66805 572056 66810 572112
rect 66866 572056 68908 572112
rect 66805 572054 68908 572056
rect 66805 572051 66871 572054
rect 91185 571434 91251 571437
rect 88596 571432 91251 571434
rect 88596 571376 91190 571432
rect 91246 571376 91251 571432
rect 88596 571374 91251 571376
rect 91185 571371 91251 571374
rect 67081 570754 67147 570757
rect 67449 570754 67515 570757
rect 67081 570752 68908 570754
rect 67081 570696 67086 570752
rect 67142 570696 67454 570752
rect 67510 570696 68908 570752
rect 67081 570694 68908 570696
rect 67081 570691 67147 570694
rect 67449 570691 67515 570694
rect 93117 570074 93183 570077
rect 88596 570072 93183 570074
rect 88596 570016 93122 570072
rect 93178 570016 93183 570072
rect 88596 570014 93183 570016
rect 93117 570011 93183 570014
rect 67357 569394 67423 569397
rect 67357 569392 68908 569394
rect 67357 569336 67362 569392
rect 67418 569336 68908 569392
rect 67357 569334 68908 569336
rect 67357 569331 67423 569334
rect 91737 568714 91803 568717
rect 88596 568712 91803 568714
rect 88596 568656 91742 568712
rect 91798 568656 91803 568712
rect 88596 568654 91803 568656
rect 91737 568651 91803 568654
rect 66805 568034 66871 568037
rect 66805 568032 68908 568034
rect 66805 567976 66810 568032
rect 66866 567976 68908 568032
rect 66805 567974 68908 567976
rect 66805 567971 66871 567974
rect 89805 567354 89871 567357
rect 88596 567352 89871 567354
rect 88596 567296 89810 567352
rect 89866 567296 89871 567352
rect 88596 567294 89871 567296
rect 89805 567291 89871 567294
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 67633 566674 67699 566677
rect 67633 566672 68908 566674
rect 67633 566616 67638 566672
rect 67694 566616 68908 566672
rect 67633 566614 68908 566616
rect 67633 566611 67699 566614
rect 91553 565858 91619 565861
rect 88596 565856 91619 565858
rect 88596 565800 91558 565856
rect 91614 565800 91619 565856
rect 88596 565798 91619 565800
rect 91553 565795 91619 565798
rect 66805 565042 66871 565045
rect 66805 565040 68908 565042
rect 66805 564984 66810 565040
rect 66866 564984 68908 565040
rect 66805 564982 68908 564984
rect 66805 564979 66871 564982
rect 91553 564498 91619 564501
rect 88596 564496 91619 564498
rect 88596 564440 91558 564496
rect 91614 564440 91619 564496
rect 88596 564438 91619 564440
rect 91553 564435 91619 564438
rect 582373 564362 582439 564365
rect 583520 564362 584960 564452
rect 582373 564360 584960 564362
rect 582373 564304 582378 564360
rect 582434 564304 584960 564360
rect 582373 564302 584960 564304
rect 582373 564299 582439 564302
rect 583520 564212 584960 564302
rect 66805 563682 66871 563685
rect 66805 563680 68908 563682
rect 66805 563624 66810 563680
rect 66866 563624 68908 563680
rect 66805 563622 68908 563624
rect 66805 563619 66871 563622
rect 91553 563138 91619 563141
rect 88596 563136 91619 563138
rect 88596 563080 91558 563136
rect 91614 563080 91619 563136
rect 88596 563078 91619 563080
rect 91553 563075 91619 563078
rect 66805 562322 66871 562325
rect 66805 562320 68908 562322
rect 66805 562264 66810 562320
rect 66866 562264 68908 562320
rect 66805 562262 68908 562264
rect 66805 562259 66871 562262
rect 91185 561506 91251 561509
rect 88596 561504 91251 561506
rect 88596 561448 91190 561504
rect 91246 561448 91251 561504
rect 88596 561446 91251 561448
rect 91185 561443 91251 561446
rect 66805 560962 66871 560965
rect 66805 560960 68908 560962
rect 66805 560904 66810 560960
rect 66866 560904 68908 560960
rect 66805 560902 68908 560904
rect 66805 560899 66871 560902
rect 88885 560146 88951 560149
rect 89621 560146 89687 560149
rect 88596 560144 89687 560146
rect 88596 560088 88890 560144
rect 88946 560088 89626 560144
rect 89682 560088 89687 560144
rect 88596 560086 89687 560088
rect 88885 560083 88951 560086
rect 89621 560083 89687 560086
rect 66069 559602 66135 559605
rect 66069 559600 68908 559602
rect 66069 559544 66074 559600
rect 66130 559544 68908 559600
rect 66069 559542 68908 559544
rect 66069 559539 66135 559542
rect 205633 559058 205699 559061
rect 583109 559058 583175 559061
rect 205633 559056 583175 559058
rect 205633 559000 205638 559056
rect 205694 559000 583114 559056
rect 583170 559000 583175 559056
rect 205633 558998 583175 559000
rect 205633 558995 205699 558998
rect 583109 558995 583175 558998
rect 92289 558786 92355 558789
rect 88596 558784 92355 558786
rect 88596 558728 92294 558784
rect 92350 558728 92355 558784
rect 88596 558726 92355 558728
rect 92289 558723 92355 558726
rect 66805 558242 66871 558245
rect 66805 558240 68908 558242
rect 66805 558184 66810 558240
rect 66866 558184 68908 558240
rect 66805 558182 68908 558184
rect 66805 558179 66871 558182
rect 166206 557500 166212 557564
rect 166276 557562 166282 557564
rect 231853 557562 231919 557565
rect 166276 557560 231919 557562
rect 166276 557504 231858 557560
rect 231914 557504 231919 557560
rect 166276 557502 231919 557504
rect 166276 557500 166282 557502
rect 231853 557499 231919 557502
rect 91093 557426 91159 557429
rect 88596 557424 91159 557426
rect 88596 557368 91098 557424
rect 91154 557368 91159 557424
rect 88596 557366 91159 557368
rect 91093 557363 91159 557366
rect 66662 556820 66668 556884
rect 66732 556882 66738 556884
rect 66732 556822 68908 556882
rect 66732 556820 66738 556822
rect 187049 556202 187115 556205
rect 243537 556202 243603 556205
rect 187049 556200 243603 556202
rect 187049 556144 187054 556200
rect 187110 556144 243542 556200
rect 243598 556144 243603 556200
rect 187049 556142 243603 556144
rect 187049 556139 187115 556142
rect 243537 556139 243603 556142
rect 91093 556066 91159 556069
rect 88596 556064 91159 556066
rect 88596 556008 91098 556064
rect 91154 556008 91159 556064
rect 88596 556006 91159 556008
rect 91093 556003 91159 556006
rect 66805 555522 66871 555525
rect 66805 555520 68908 555522
rect 66805 555464 66810 555520
rect 66866 555464 68908 555520
rect 66805 555462 68908 555464
rect 66805 555459 66871 555462
rect 184841 554842 184907 554845
rect 240225 554842 240291 554845
rect 184841 554840 240291 554842
rect 184841 554784 184846 554840
rect 184902 554784 240230 554840
rect 240286 554784 240291 554840
rect 184841 554782 240291 554784
rect 184841 554779 184907 554782
rect 240225 554779 240291 554782
rect 66621 554162 66687 554165
rect 67541 554162 67607 554165
rect 66621 554160 68908 554162
rect 66621 554104 66626 554160
rect 66682 554104 67546 554160
rect 67602 554104 68908 554160
rect 66621 554102 68908 554104
rect 66621 554099 66687 554102
rect 67541 554099 67607 554102
rect -960 553890 480 553980
rect 2773 553890 2839 553893
rect -960 553888 2839 553890
rect -960 553832 2778 553888
rect 2834 553832 2839 553888
rect -960 553830 2839 553832
rect 88566 553890 88626 554676
rect 198549 554026 198615 554029
rect 582741 554026 582807 554029
rect 198549 554024 582807 554026
rect 198549 553968 198554 554024
rect 198610 553968 582746 554024
rect 582802 553968 582807 554024
rect 198549 553966 582807 553968
rect 198549 553963 198615 553966
rect 582741 553963 582807 553966
rect 88566 553830 93870 553890
rect -960 553740 480 553830
rect 2773 553827 2839 553830
rect 93810 553482 93870 553830
rect 115054 553482 115060 553484
rect 93810 553422 115060 553482
rect 115054 553420 115060 553422
rect 115124 553420 115130 553484
rect 91369 553346 91435 553349
rect 88596 553344 91435 553346
rect 88596 553288 91374 553344
rect 91430 553288 91435 553344
rect 88596 553286 91435 553288
rect 91369 553283 91435 553286
rect 67449 552802 67515 552805
rect 67449 552800 68908 552802
rect 67449 552744 67454 552800
rect 67510 552744 68908 552800
rect 67449 552742 68908 552744
rect 67449 552739 67515 552742
rect 91093 552122 91159 552125
rect 88596 552120 91159 552122
rect 88596 552064 91098 552120
rect 91154 552064 91159 552120
rect 88596 552062 91159 552064
rect 91093 552059 91159 552062
rect 169109 552122 169175 552125
rect 290089 552122 290155 552125
rect 169109 552120 290155 552122
rect 169109 552064 169114 552120
rect 169170 552064 290094 552120
rect 290150 552064 290155 552120
rect 169109 552062 290155 552064
rect 169109 552059 169175 552062
rect 290089 552059 290155 552062
rect 67541 551442 67607 551445
rect 67541 551440 68908 551442
rect 67541 551384 67546 551440
rect 67602 551384 68908 551440
rect 67541 551382 68908 551384
rect 67541 551379 67607 551382
rect 583520 551020 584960 551260
rect 191189 550898 191255 550901
rect 205633 550898 205699 550901
rect 191189 550896 205699 550898
rect 191189 550840 191194 550896
rect 191250 550840 205638 550896
rect 205694 550840 205699 550896
rect 191189 550838 205699 550840
rect 191189 550835 191255 550838
rect 205633 550835 205699 550838
rect 91093 550762 91159 550765
rect 88596 550760 91159 550762
rect 88596 550704 91098 550760
rect 91154 550704 91159 550760
rect 88596 550702 91159 550704
rect 91093 550699 91159 550702
rect 193949 550762 194015 550765
rect 253933 550762 253999 550765
rect 193949 550760 253999 550762
rect 193949 550704 193954 550760
rect 194010 550704 253938 550760
rect 253994 550704 253999 550760
rect 193949 550702 253999 550704
rect 193949 550699 194015 550702
rect 253933 550699 253999 550702
rect 66805 550082 66871 550085
rect 66805 550080 68908 550082
rect 66805 550024 66810 550080
rect 66866 550024 68908 550080
rect 66805 550022 68908 550024
rect 66805 550019 66871 550022
rect 91093 549402 91159 549405
rect 88596 549400 91159 549402
rect 88596 549344 91098 549400
rect 91154 549344 91159 549400
rect 88596 549342 91159 549344
rect 91093 549339 91159 549342
rect 185669 549402 185735 549405
rect 304993 549402 305059 549405
rect 185669 549400 305059 549402
rect 185669 549344 185674 549400
rect 185730 549344 304998 549400
rect 305054 549344 305059 549400
rect 185669 549342 305059 549344
rect 185669 549339 185735 549342
rect 304993 549339 305059 549342
rect 66805 548722 66871 548725
rect 66805 548720 68908 548722
rect 66805 548664 66810 548720
rect 66866 548664 68908 548720
rect 66805 548662 68908 548664
rect 66805 548659 66871 548662
rect 91277 547906 91343 547909
rect 88596 547904 91343 547906
rect 88596 547848 91282 547904
rect 91338 547848 91343 547904
rect 88596 547846 91343 547848
rect 91142 547773 91202 547846
rect 91277 547843 91343 547846
rect 160686 547844 160692 547908
rect 160756 547906 160762 547908
rect 328453 547906 328519 547909
rect 160756 547904 328519 547906
rect 160756 547848 328458 547904
rect 328514 547848 328519 547904
rect 160756 547846 328519 547848
rect 160756 547844 160762 547846
rect 328453 547843 328519 547846
rect 91093 547768 91202 547773
rect 91093 547712 91098 547768
rect 91154 547712 91202 547768
rect 91093 547710 91202 547712
rect 91093 547707 91159 547710
rect 66805 547362 66871 547365
rect 66805 547360 68908 547362
rect 66805 547304 66810 547360
rect 66866 547304 68908 547360
rect 66805 547302 68908 547304
rect 66805 547299 66871 547302
rect 201033 546682 201099 546685
rect 273253 546682 273319 546685
rect 201033 546680 273319 546682
rect 201033 546624 201038 546680
rect 201094 546624 273258 546680
rect 273314 546624 273319 546680
rect 201033 546622 273319 546624
rect 201033 546619 201099 546622
rect 273253 546619 273319 546622
rect 295333 546682 295399 546685
rect 353334 546682 353340 546684
rect 295333 546680 353340 546682
rect 295333 546624 295338 546680
rect 295394 546624 353340 546680
rect 295333 546622 353340 546624
rect 295333 546619 295399 546622
rect 353334 546620 353340 546622
rect 353404 546620 353410 546684
rect 91502 546546 91508 546548
rect 88596 546486 91508 546546
rect 91502 546484 91508 546486
rect 91572 546484 91578 546548
rect 126881 546546 126947 546549
rect 339953 546546 340019 546549
rect 126881 546544 340019 546546
rect 126881 546488 126886 546544
rect 126942 546488 339958 546544
rect 340014 546488 340019 546544
rect 126881 546486 340019 546488
rect 126881 546483 126947 546486
rect 339953 546483 340019 546486
rect 66805 546002 66871 546005
rect 66805 546000 68908 546002
rect 66805 545944 66810 546000
rect 66866 545944 68908 546000
rect 66805 545942 68908 545944
rect 66805 545939 66871 545942
rect 191046 545260 191052 545324
rect 191116 545322 191122 545324
rect 225321 545322 225387 545325
rect 191116 545320 225387 545322
rect 191116 545264 225326 545320
rect 225382 545264 225387 545320
rect 191116 545262 225387 545264
rect 191116 545260 191122 545262
rect 225321 545259 225387 545262
rect 91553 545186 91619 545189
rect 88596 545184 91619 545186
rect 88596 545128 91558 545184
rect 91614 545128 91619 545184
rect 88596 545126 91619 545128
rect 91553 545123 91619 545126
rect 200798 545124 200804 545188
rect 200868 545186 200874 545188
rect 255313 545186 255379 545189
rect 200868 545184 255379 545186
rect 200868 545128 255318 545184
rect 255374 545128 255379 545184
rect 200868 545126 255379 545128
rect 200868 545124 200874 545126
rect 255313 545123 255379 545126
rect 66805 544642 66871 544645
rect 66805 544640 68908 544642
rect 66805 544584 66810 544640
rect 66866 544584 68908 544640
rect 66805 544582 68908 544584
rect 66805 544579 66871 544582
rect 298369 544098 298435 544101
rect 352046 544098 352052 544100
rect 298369 544096 352052 544098
rect 298369 544040 298374 544096
rect 298430 544040 352052 544096
rect 298369 544038 352052 544040
rect 298369 544035 298435 544038
rect 352046 544036 352052 544038
rect 352116 544036 352122 544100
rect 181294 543900 181300 543964
rect 181364 543962 181370 543964
rect 306649 543962 306715 543965
rect 181364 543960 306715 543962
rect 181364 543904 306654 543960
rect 306710 543904 306715 543960
rect 181364 543902 306715 543904
rect 181364 543900 181370 543902
rect 306649 543899 306715 543902
rect 93761 543826 93827 543829
rect 357617 543826 357683 543829
rect 360837 543826 360903 543829
rect 88596 543824 360903 543826
rect 88596 543768 93766 543824
rect 93822 543768 357622 543824
rect 357678 543768 360842 543824
rect 360898 543768 360903 543824
rect 88596 543766 360903 543768
rect 93761 543763 93827 543766
rect 357617 543763 357683 543766
rect 360837 543763 360903 543766
rect 66805 543282 66871 543285
rect 66805 543280 68908 543282
rect 66805 543224 66810 543280
rect 66866 543224 68908 543280
rect 66805 543222 68908 543224
rect 66805 543219 66871 543222
rect 67357 543010 67423 543013
rect 68686 543010 68692 543012
rect 67357 543008 68692 543010
rect 67357 542952 67362 543008
rect 67418 542952 68692 543008
rect 67357 542950 68692 542952
rect 67357 542947 67423 542950
rect 68686 542948 68692 542950
rect 68756 542948 68762 543012
rect 195237 542738 195303 542741
rect 261753 542738 261819 542741
rect 195237 542736 261819 542738
rect 195237 542680 195242 542736
rect 195298 542680 261758 542736
rect 261814 542680 261819 542736
rect 195237 542678 261819 542680
rect 195237 542675 195303 542678
rect 261753 542675 261819 542678
rect 142061 542602 142127 542605
rect 283465 542602 283531 542605
rect 142061 542600 283531 542602
rect 142061 542544 142066 542600
rect 142122 542544 283470 542600
rect 283526 542544 283531 542600
rect 142061 542542 283531 542544
rect 142061 542539 142127 542542
rect 283465 542539 283531 542542
rect 91553 542466 91619 542469
rect 88596 542464 91619 542466
rect 88596 542408 91558 542464
rect 91614 542408 91619 542464
rect 88596 542406 91619 542408
rect 91553 542403 91619 542406
rect 161238 542404 161244 542468
rect 161308 542466 161314 542468
rect 348233 542466 348299 542469
rect 161308 542464 348299 542466
rect 161308 542408 348238 542464
rect 348294 542408 348299 542464
rect 161308 542406 348299 542408
rect 161308 542404 161314 542406
rect 348233 542403 348299 542406
rect 356053 542468 356119 542469
rect 356053 542464 356100 542468
rect 356164 542466 356170 542468
rect 356053 542408 356058 542464
rect 356053 542404 356100 542408
rect 356164 542406 356210 542466
rect 356164 542404 356170 542406
rect 356053 542403 356119 542404
rect 66989 541922 67055 541925
rect 66989 541920 68908 541922
rect 66989 541864 66994 541920
rect 67050 541864 68908 541920
rect 66989 541862 68908 541864
rect 66989 541859 67055 541862
rect 88190 541452 88196 541516
rect 88260 541514 88266 541516
rect 323577 541514 323643 541517
rect 88260 541512 323643 541514
rect 88260 541456 323582 541512
rect 323638 541456 323643 541512
rect 88260 541454 323643 541456
rect 88260 541452 88266 541454
rect 323577 541451 323643 541454
rect 91502 541180 91508 541244
rect 91572 541242 91578 541244
rect 91572 541182 93870 541242
rect 91572 541180 91578 541182
rect 91921 541106 91987 541109
rect 88596 541104 91987 541106
rect 88596 541048 91926 541104
rect 91982 541048 91987 541104
rect 88596 541046 91987 541048
rect 93810 541106 93870 541182
rect 197854 541180 197860 541244
rect 197924 541242 197930 541244
rect 262213 541242 262279 541245
rect 197924 541240 262279 541242
rect 197924 541184 262218 541240
rect 262274 541184 262279 541240
rect 197924 541182 262279 541184
rect 197924 541180 197930 541182
rect 262213 541179 262279 541182
rect 318241 541242 318307 541245
rect 352230 541242 352236 541244
rect 318241 541240 352236 541242
rect 318241 541184 318246 541240
rect 318302 541184 352236 541240
rect 318241 541182 352236 541184
rect 318241 541179 318307 541182
rect 352230 541180 352236 541182
rect 352300 541180 352306 541244
rect 94589 541106 94655 541109
rect 93810 541104 94655 541106
rect 93810 541048 94594 541104
rect 94650 541048 94655 541104
rect 93810 541046 94655 541048
rect 91921 541043 91987 541046
rect 94589 541043 94655 541046
rect 196709 541106 196775 541109
rect 203609 541106 203675 541109
rect 196709 541104 203675 541106
rect 196709 541048 196714 541104
rect 196770 541048 203614 541104
rect 203670 541048 203675 541104
rect 196709 541046 203675 541048
rect 196709 541043 196775 541046
rect 203609 541043 203675 541046
rect 349981 541106 350047 541109
rect 388437 541106 388503 541109
rect 349981 541104 388503 541106
rect 349981 541048 349986 541104
rect 350042 541048 388442 541104
rect 388498 541048 388503 541104
rect 349981 541046 388503 541048
rect 349981 541043 350047 541046
rect 388437 541043 388503 541046
rect -960 540684 480 540924
rect 67541 540562 67607 540565
rect 67541 540560 68908 540562
rect 67541 540504 67546 540560
rect 67602 540504 68908 540560
rect 67541 540502 68908 540504
rect 67541 540499 67607 540502
rect 88793 540154 88859 540157
rect 357525 540154 357591 540157
rect 88793 540152 357591 540154
rect 88793 540096 88798 540152
rect 88854 540096 357530 540152
rect 357586 540096 357591 540152
rect 88793 540094 357591 540096
rect 88793 540091 88859 540094
rect 357525 540091 357591 540094
rect 184197 539882 184263 539885
rect 280613 539882 280679 539885
rect 184197 539880 280679 539882
rect 184197 539824 184202 539880
rect 184258 539824 280618 539880
rect 280674 539824 280679 539880
rect 184197 539822 280679 539824
rect 184197 539819 184263 539822
rect 280613 539819 280679 539822
rect 93117 539746 93183 539749
rect 88596 539744 93183 539746
rect 88596 539688 93122 539744
rect 93178 539688 93183 539744
rect 88596 539686 93183 539688
rect 93117 539683 93183 539686
rect 159214 539684 159220 539748
rect 159284 539746 159290 539748
rect 322013 539746 322079 539749
rect 159284 539744 322079 539746
rect 159284 539688 322018 539744
rect 322074 539688 322079 539744
rect 159284 539686 322079 539688
rect 159284 539684 159290 539686
rect 322013 539683 322079 539686
rect 48221 539610 48287 539613
rect 67541 539610 67607 539613
rect 48221 539608 67607 539610
rect 48221 539552 48226 539608
rect 48282 539552 67546 539608
rect 67602 539552 67607 539608
rect 48221 539550 67607 539552
rect 48221 539547 48287 539550
rect 67541 539547 67607 539550
rect 270677 539610 270743 539613
rect 273989 539610 274055 539613
rect 270677 539608 274055 539610
rect 270677 539552 270682 539608
rect 270738 539552 273994 539608
rect 274050 539552 274055 539608
rect 270677 539550 274055 539552
rect 270677 539547 270743 539550
rect 273989 539547 274055 539550
rect 67357 539474 67423 539477
rect 169109 539474 169175 539477
rect 67357 539472 169175 539474
rect 67357 539416 67362 539472
rect 67418 539416 169114 539472
rect 169170 539416 169175 539472
rect 67357 539414 169175 539416
rect 67357 539411 67423 539414
rect 169109 539411 169175 539414
rect 92381 538930 92447 538933
rect 99966 538930 99972 538932
rect 92381 538928 99972 538930
rect 92381 538872 92386 538928
rect 92442 538872 99972 538928
rect 92381 538870 99972 538872
rect 92381 538867 92447 538870
rect 99966 538868 99972 538870
rect 100036 538868 100042 538932
rect 93761 538794 93827 538797
rect 106406 538794 106412 538796
rect 93761 538792 106412 538794
rect 93761 538736 93766 538792
rect 93822 538736 106412 538792
rect 93761 538734 106412 538736
rect 93761 538731 93827 538734
rect 106406 538732 106412 538734
rect 106476 538732 106482 538796
rect 195094 538460 195100 538524
rect 195164 538522 195170 538524
rect 222469 538522 222535 538525
rect 195164 538520 222535 538522
rect 195164 538464 222474 538520
rect 222530 538464 222535 538520
rect 195164 538462 222535 538464
rect 195164 538460 195170 538462
rect 222469 538459 222535 538462
rect 223205 538522 223271 538525
rect 265525 538522 265591 538525
rect 223205 538520 265591 538522
rect 223205 538464 223210 538520
rect 223266 538464 265530 538520
rect 265586 538464 265591 538520
rect 223205 538462 265591 538464
rect 223205 538459 223271 538462
rect 265525 538459 265591 538462
rect 337101 538522 337167 538525
rect 362953 538522 363019 538525
rect 337101 538520 363019 538522
rect 337101 538464 337106 538520
rect 337162 538464 362958 538520
rect 363014 538464 363019 538520
rect 337101 538462 363019 538464
rect 337101 538459 337167 538462
rect 362953 538459 363019 538462
rect 198733 538386 198799 538389
rect 356237 538386 356303 538389
rect 198733 538384 356303 538386
rect 198733 538328 198738 538384
rect 198794 538328 356242 538384
rect 356298 538328 356303 538384
rect 198733 538326 356303 538328
rect 198733 538323 198799 538326
rect 356237 538323 356303 538326
rect 188889 538250 188955 538253
rect 217501 538250 217567 538253
rect 188889 538248 217567 538250
rect 188889 538192 188894 538248
rect 188950 538192 217506 538248
rect 217562 538192 217567 538248
rect 188889 538190 217567 538192
rect 188889 538187 188955 538190
rect 217501 538187 217567 538190
rect 221089 538250 221155 538253
rect 580257 538250 580323 538253
rect 221089 538248 580323 538250
rect 221089 538192 221094 538248
rect 221150 538192 580262 538248
rect 580318 538192 580323 538248
rect 221089 538190 580323 538192
rect 221089 538187 221155 538190
rect 580257 538187 580323 538190
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 192569 537162 192635 537165
rect 335445 537162 335511 537165
rect 192569 537160 335511 537162
rect 192569 537104 192574 537160
rect 192630 537104 335450 537160
rect 335506 537104 335511 537160
rect 192569 537102 335511 537104
rect 192569 537099 192635 537102
rect 335445 537099 335511 537102
rect 177297 537026 177363 537029
rect 333789 537026 333855 537029
rect 177297 537024 333855 537026
rect 177297 536968 177302 537024
rect 177358 536968 333794 537024
rect 333850 536968 333855 537024
rect 177297 536966 333855 536968
rect 177297 536963 177363 536966
rect 333789 536963 333855 536966
rect 130469 536890 130535 536893
rect 353661 536890 353727 536893
rect 130469 536888 353727 536890
rect 130469 536832 130474 536888
rect 130530 536832 353666 536888
rect 353722 536832 353727 536888
rect 130469 536830 353727 536832
rect 130469 536827 130535 536830
rect 353661 536827 353727 536830
rect 72601 536754 72667 536757
rect 88190 536754 88196 536756
rect 72601 536752 88196 536754
rect 72601 536696 72606 536752
rect 72662 536696 88196 536752
rect 72601 536694 88196 536696
rect 72601 536691 72667 536694
rect 88190 536692 88196 536694
rect 88260 536692 88266 536756
rect 22737 536074 22803 536077
rect 44081 536074 44147 536077
rect 73153 536074 73219 536077
rect 22737 536072 73219 536074
rect 22737 536016 22742 536072
rect 22798 536016 44086 536072
rect 44142 536016 73158 536072
rect 73214 536016 73219 536072
rect 22737 536014 73219 536016
rect 22737 536011 22803 536014
rect 44081 536011 44147 536014
rect 73153 536011 73219 536014
rect 80053 535802 80119 535805
rect 308397 535802 308463 535805
rect 80053 535800 308463 535802
rect 80053 535744 80058 535800
rect 80114 535744 308402 535800
rect 308458 535744 308463 535800
rect 80053 535742 308463 535744
rect 80053 535739 80119 535742
rect 308397 535739 308463 535742
rect 173249 535666 173315 535669
rect 276013 535666 276079 535669
rect 276933 535666 276999 535669
rect 173249 535664 276999 535666
rect 173249 535608 173254 535664
rect 173310 535608 276018 535664
rect 276074 535608 276938 535664
rect 276994 535608 276999 535664
rect 173249 535606 276999 535608
rect 173249 535603 173315 535606
rect 276013 535603 276079 535606
rect 276933 535603 276999 535606
rect 69565 535532 69631 535533
rect 69565 535530 69612 535532
rect 69520 535528 69612 535530
rect 69520 535472 69570 535528
rect 69520 535470 69612 535472
rect 69565 535468 69612 535470
rect 69676 535468 69682 535532
rect 199326 535468 199332 535532
rect 199396 535530 199402 535532
rect 208669 535530 208735 535533
rect 199396 535528 208735 535530
rect 199396 535472 208674 535528
rect 208730 535472 208735 535528
rect 199396 535470 208735 535472
rect 199396 535468 199402 535470
rect 69565 535467 69631 535468
rect 208669 535467 208735 535470
rect 304073 535530 304139 535533
rect 389173 535530 389239 535533
rect 304073 535528 389239 535530
rect 304073 535472 304078 535528
rect 304134 535472 389178 535528
rect 389234 535472 389239 535528
rect 304073 535470 389239 535472
rect 304073 535467 304139 535470
rect 389173 535467 389239 535470
rect 67766 535332 67772 535396
rect 67836 535394 67842 535396
rect 76557 535394 76623 535397
rect 67836 535392 76623 535394
rect 67836 535336 76562 535392
rect 76618 535336 76623 535392
rect 67836 535334 76623 535336
rect 67836 535332 67842 535334
rect 76557 535331 76623 535334
rect 199745 535394 199811 535397
rect 200389 535394 200455 535397
rect 201033 535394 201099 535397
rect 221089 535394 221155 535397
rect 199745 535392 200455 535394
rect 199745 535336 199750 535392
rect 199806 535336 200394 535392
rect 200450 535336 200455 535392
rect 199745 535334 200455 535336
rect 199745 535331 199811 535334
rect 200389 535331 200455 535334
rect 200622 535392 201099 535394
rect 200622 535336 201038 535392
rect 201094 535336 201099 535392
rect 200622 535334 201099 535336
rect 199878 535196 199884 535260
rect 199948 535258 199954 535260
rect 200622 535258 200682 535334
rect 201033 535331 201099 535334
rect 209730 535392 221155 535394
rect 209730 535336 221094 535392
rect 221150 535336 221155 535392
rect 209730 535334 221155 535336
rect 199948 535198 200682 535258
rect 199948 535196 199954 535198
rect 191741 534986 191807 534989
rect 209730 534986 209790 535334
rect 221089 535331 221155 535334
rect 191741 534984 209790 534986
rect 191741 534928 191746 534984
rect 191802 534928 209790 534984
rect 191741 534926 209790 534928
rect 191741 534923 191807 534926
rect 4797 534714 4863 534717
rect 94589 534714 94655 534717
rect 357617 534714 357683 534717
rect 4797 534712 94655 534714
rect 4797 534656 4802 534712
rect 4858 534656 94594 534712
rect 94650 534656 94655 534712
rect 4797 534654 94655 534656
rect 356132 534712 357683 534714
rect 356132 534656 357622 534712
rect 357678 534656 357683 534712
rect 356132 534654 357683 534656
rect 4797 534651 4863 534654
rect 94589 534651 94655 534654
rect 357617 534651 357683 534654
rect 188981 534170 189047 534173
rect 200070 534170 200130 534548
rect 188981 534168 200130 534170
rect 188981 534112 188986 534168
rect 189042 534112 200130 534168
rect 188981 534110 200130 534112
rect 188981 534107 189047 534110
rect 182817 533354 182883 533357
rect 199745 533354 199811 533357
rect 182817 533352 199811 533354
rect 182817 533296 182822 533352
rect 182878 533296 199750 533352
rect 199806 533296 199811 533352
rect 182817 533294 199811 533296
rect 182817 533291 182883 533294
rect 199745 533291 199811 533294
rect 197445 532266 197511 532269
rect 197445 532264 200100 532266
rect 197445 532208 197450 532264
rect 197506 532208 200100 532264
rect 197445 532206 200100 532208
rect 197445 532203 197511 532206
rect 358721 532130 358787 532133
rect 356132 532128 358787 532130
rect 356132 532072 358726 532128
rect 358782 532072 358787 532128
rect 356132 532070 358787 532072
rect 358721 532067 358787 532070
rect 197445 529818 197511 529821
rect 198549 529818 198615 529821
rect 197445 529816 200100 529818
rect 197445 529760 197450 529816
rect 197506 529760 198554 529816
rect 198610 529760 200100 529816
rect 197445 529758 200100 529760
rect 197445 529755 197511 529758
rect 198549 529755 198615 529758
rect 358721 529682 358787 529685
rect 356132 529680 358787 529682
rect 356132 529624 358726 529680
rect 358782 529624 358787 529680
rect 356132 529622 358787 529624
rect 358721 529619 358787 529622
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 170397 527778 170463 527781
rect 199326 527778 199332 527780
rect 170397 527776 199332 527778
rect 170397 527720 170402 527776
rect 170458 527720 199332 527776
rect 170397 527718 199332 527720
rect 170397 527715 170463 527718
rect 199326 527716 199332 527718
rect 199396 527716 199402 527780
rect 197445 527370 197511 527373
rect 197445 527368 200100 527370
rect 197445 527312 197450 527368
rect 197506 527312 200100 527368
rect 197445 527310 200100 527312
rect 197445 527307 197511 527310
rect 358721 527234 358787 527237
rect 356132 527232 358787 527234
rect 356132 527176 358726 527232
rect 358782 527176 358787 527232
rect 356132 527174 358787 527176
rect 358721 527171 358787 527174
rect 175774 526356 175780 526420
rect 175844 526418 175850 526420
rect 197854 526418 197860 526420
rect 175844 526358 197860 526418
rect 175844 526356 175850 526358
rect 197854 526356 197860 526358
rect 197924 526356 197930 526420
rect 197537 524786 197603 524789
rect 358721 524786 358787 524789
rect 197537 524784 200100 524786
rect 197537 524728 197542 524784
rect 197598 524728 200100 524784
rect 197537 524726 200100 524728
rect 356132 524784 358787 524786
rect 356132 524728 358726 524784
rect 358782 524728 358787 524784
rect 356132 524726 358787 524728
rect 197537 524723 197603 524726
rect 358721 524723 358787 524726
rect 580349 524514 580415 524517
rect 583520 524514 584960 524604
rect 580349 524512 584960 524514
rect 580349 524456 580354 524512
rect 580410 524456 584960 524512
rect 580349 524454 584960 524456
rect 580349 524451 580415 524454
rect 583520 524364 584960 524454
rect 197445 522338 197511 522341
rect 357433 522338 357499 522341
rect 358721 522338 358787 522341
rect 197445 522336 200100 522338
rect 197445 522280 197450 522336
rect 197506 522280 200100 522336
rect 197445 522278 200100 522280
rect 356132 522336 358787 522338
rect 356132 522280 357438 522336
rect 357494 522280 358726 522336
rect 358782 522280 358787 522336
rect 356132 522278 358787 522280
rect 197445 522275 197511 522278
rect 357433 522275 357499 522278
rect 358721 522275 358787 522278
rect 356329 519890 356395 519893
rect 358629 519890 358695 519893
rect 356132 519888 358695 519890
rect 163446 518876 163452 518940
rect 163516 518938 163522 518940
rect 200070 518938 200130 519860
rect 356132 519832 356334 519888
rect 356390 519832 358634 519888
rect 358690 519832 358695 519888
rect 356132 519830 358695 519832
rect 356329 519827 356395 519830
rect 358629 519827 358695 519830
rect 163516 518878 200130 518938
rect 163516 518876 163522 518878
rect 197445 517442 197511 517445
rect 358721 517442 358787 517445
rect 197445 517440 200100 517442
rect 197445 517384 197450 517440
rect 197506 517384 200100 517440
rect 197445 517382 200100 517384
rect 356132 517440 358787 517442
rect 356132 517384 358726 517440
rect 358782 517384 358787 517440
rect 356132 517382 358787 517384
rect 197445 517379 197511 517382
rect 358721 517379 358787 517382
rect 360142 514994 360148 514996
rect -960 514858 480 514948
rect 180750 514934 200100 514994
rect 356132 514934 360148 514994
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 161974 514796 161980 514860
rect 162044 514858 162050 514860
rect 180750 514858 180810 514934
rect 360142 514932 360148 514934
rect 360212 514932 360218 514996
rect 162044 514798 180810 514858
rect 162044 514796 162050 514798
rect 357525 512682 357591 512685
rect 356132 512680 357591 512682
rect 356132 512624 357530 512680
rect 357586 512624 357591 512680
rect 356132 512622 357591 512624
rect 357525 512619 357591 512622
rect 198590 512484 198596 512548
rect 198660 512546 198666 512548
rect 198660 512486 200100 512546
rect 198660 512484 198666 512486
rect 582373 511322 582439 511325
rect 583520 511322 584960 511412
rect 582373 511320 584960 511322
rect 582373 511264 582378 511320
rect 582434 511264 584960 511320
rect 582373 511262 584960 511264
rect 582373 511259 582439 511262
rect 583520 511172 584960 511262
rect 197445 510234 197511 510237
rect 197445 510232 200100 510234
rect 197445 510176 197450 510232
rect 197506 510176 200100 510232
rect 197445 510174 200100 510176
rect 197445 510171 197511 510174
rect 358077 510098 358143 510101
rect 356132 510096 358143 510098
rect 356132 510040 358082 510096
rect 358138 510040 358143 510096
rect 356132 510038 358143 510040
rect 358077 510035 358143 510038
rect 197445 507650 197511 507653
rect 358721 507650 358787 507653
rect 197445 507648 200100 507650
rect 197445 507592 197450 507648
rect 197506 507592 200100 507648
rect 197445 507590 200100 507592
rect 356132 507648 358787 507650
rect 356132 507592 358726 507648
rect 358782 507592 358787 507648
rect 356132 507590 358787 507592
rect 197445 507587 197511 507590
rect 358721 507587 358787 507590
rect 199009 505202 199075 505205
rect 358721 505202 358787 505205
rect 199009 505200 200100 505202
rect 199009 505144 199014 505200
rect 199070 505144 200100 505200
rect 199009 505142 200100 505144
rect 356132 505200 358787 505202
rect 356132 505144 358726 505200
rect 358782 505144 358787 505200
rect 356132 505142 358787 505144
rect 199009 505139 199075 505142
rect 358721 505139 358787 505142
rect 197445 502754 197511 502757
rect 358721 502754 358787 502757
rect 197445 502752 200100 502754
rect 197445 502696 197450 502752
rect 197506 502696 200100 502752
rect 197445 502694 200100 502696
rect 356132 502752 358787 502754
rect 356132 502696 358726 502752
rect 358782 502696 358787 502752
rect 356132 502694 358787 502696
rect 197445 502691 197511 502694
rect 358721 502691 358787 502694
rect -960 501802 480 501892
rect 2773 501802 2839 501805
rect -960 501800 2839 501802
rect -960 501744 2778 501800
rect 2834 501744 2839 501800
rect -960 501742 2839 501744
rect -960 501652 480 501742
rect 2773 501739 2839 501742
rect 197445 500442 197511 500445
rect 198641 500442 198707 500445
rect 197445 500440 200100 500442
rect 197445 500384 197450 500440
rect 197506 500384 198646 500440
rect 198702 500384 200100 500440
rect 197445 500382 200100 500384
rect 197445 500379 197511 500382
rect 198641 500379 198707 500382
rect 356102 499898 356162 500276
rect 356278 499898 356284 499900
rect 356102 499838 356284 499898
rect 356278 499836 356284 499838
rect 356348 499836 356354 499900
rect 358721 497858 358787 497861
rect 356132 497856 358787 497858
rect 168966 496844 168972 496908
rect 169036 496906 169042 496908
rect 200070 496906 200130 497828
rect 356132 497800 358726 497856
rect 358782 497800 358787 497856
rect 583520 497844 584960 498084
rect 356132 497798 358787 497800
rect 358721 497795 358787 497798
rect 169036 496846 200130 496906
rect 169036 496844 169042 496846
rect 197445 495546 197511 495549
rect 358629 495546 358695 495549
rect 197445 495544 200100 495546
rect 197445 495488 197450 495544
rect 197506 495488 200100 495544
rect 197445 495486 200100 495488
rect 356132 495544 358695 495546
rect 356132 495488 358634 495544
rect 358690 495488 358695 495544
rect 356132 495486 358695 495488
rect 197445 495483 197511 495486
rect 358629 495483 358695 495486
rect 197445 492962 197511 492965
rect 358721 492962 358787 492965
rect 197445 492960 200100 492962
rect 197445 492904 197450 492960
rect 197506 492904 200100 492960
rect 197445 492902 200100 492904
rect 356132 492960 358787 492962
rect 356132 492904 358726 492960
rect 358782 492904 358787 492960
rect 356132 492902 358787 492904
rect 197445 492899 197511 492902
rect 358721 492899 358787 492902
rect 356237 490922 356303 490925
rect 356102 490920 356303 490922
rect 356102 490864 356242 490920
rect 356298 490864 356303 490920
rect 356102 490862 356303 490864
rect 197445 490514 197511 490517
rect 197445 490512 200100 490514
rect 197445 490456 197450 490512
rect 197506 490456 200100 490512
rect 197445 490454 200100 490456
rect 197445 490451 197511 490454
rect 356102 490348 356162 490862
rect 356237 490859 356303 490862
rect -960 488596 480 488836
rect 197445 488066 197511 488069
rect 197445 488064 200100 488066
rect 197445 488008 197450 488064
rect 197506 488008 200100 488064
rect 197445 488006 200100 488008
rect 197445 488003 197511 488006
rect 358721 487794 358787 487797
rect 356132 487792 358787 487794
rect 356132 487736 358726 487792
rect 358782 487736 358787 487792
rect 356132 487734 358787 487736
rect 358721 487731 358787 487734
rect 197445 485618 197511 485621
rect 197445 485616 200100 485618
rect 197445 485560 197450 485616
rect 197506 485560 200100 485616
rect 197445 485558 200100 485560
rect 197445 485555 197511 485558
rect 358169 485346 358235 485349
rect 356132 485344 358235 485346
rect 356132 485288 358174 485344
rect 358230 485288 358235 485344
rect 356132 485286 358235 485288
rect 358169 485283 358235 485286
rect 580257 484666 580323 484669
rect 583520 484666 584960 484756
rect 580257 484664 584960 484666
rect 580257 484608 580262 484664
rect 580318 484608 584960 484664
rect 580257 484606 584960 484608
rect 580257 484603 580323 484606
rect 583520 484516 584960 484606
rect 197997 483170 198063 483173
rect 197997 483168 200100 483170
rect 197997 483112 198002 483168
rect 198058 483112 200100 483168
rect 197997 483110 200100 483112
rect 197997 483107 198063 483110
rect 357893 482898 357959 482901
rect 356132 482896 357959 482898
rect 356132 482840 357898 482896
rect 357954 482840 357959 482896
rect 356132 482838 357959 482840
rect 357893 482835 357959 482838
rect 197445 480722 197511 480725
rect 197445 480720 200100 480722
rect 197445 480664 197450 480720
rect 197506 480664 200100 480720
rect 197445 480662 200100 480664
rect 197445 480659 197511 480662
rect 356102 480178 356162 480420
rect 356278 480178 356284 480180
rect 356102 480118 356284 480178
rect 356278 480116 356284 480118
rect 356348 480116 356354 480180
rect 197445 478274 197511 478277
rect 197445 478272 200100 478274
rect 197445 478216 197450 478272
rect 197506 478216 200100 478272
rect 197445 478214 200100 478216
rect 197445 478211 197511 478214
rect 357893 478002 357959 478005
rect 356132 478000 357959 478002
rect 356132 477944 357898 478000
rect 357954 477944 357959 478000
rect 356132 477942 357959 477944
rect 357893 477939 357959 477942
rect 197445 475826 197511 475829
rect 197445 475824 200100 475826
rect -960 475690 480 475780
rect 197445 475768 197450 475824
rect 197506 475768 200100 475824
rect 197445 475766 200100 475768
rect 197445 475763 197511 475766
rect 3509 475690 3575 475693
rect -960 475688 3575 475690
rect -960 475632 3514 475688
rect 3570 475632 3575 475688
rect -960 475630 3575 475632
rect -960 475540 480 475630
rect 3509 475627 3575 475630
rect 358721 475554 358787 475557
rect 356132 475552 358787 475554
rect 356132 475496 358726 475552
rect 358782 475496 358787 475552
rect 356132 475494 358787 475496
rect 358721 475491 358787 475494
rect 197445 473378 197511 473381
rect 197445 473376 200100 473378
rect 197445 473320 197450 473376
rect 197506 473320 200100 473376
rect 197445 473318 200100 473320
rect 197445 473315 197511 473318
rect 358721 473106 358787 473109
rect 356132 473104 358787 473106
rect 356132 473048 358726 473104
rect 358782 473048 358787 473104
rect 356132 473046 358787 473048
rect 358721 473043 358787 473046
rect 583017 471474 583083 471477
rect 583520 471474 584960 471564
rect 583017 471472 584960 471474
rect 583017 471416 583022 471472
rect 583078 471416 584960 471472
rect 583017 471414 584960 471416
rect 583017 471411 583083 471414
rect 583520 471324 584960 471414
rect 95969 471202 96035 471205
rect 104934 471202 104940 471204
rect 95969 471200 104940 471202
rect 95969 471144 95974 471200
rect 96030 471144 104940 471200
rect 95969 471142 104940 471144
rect 95969 471139 96035 471142
rect 104934 471140 104940 471142
rect 105004 471140 105010 471204
rect 197077 470930 197143 470933
rect 197077 470928 200100 470930
rect 197077 470872 197082 470928
rect 197138 470872 200100 470928
rect 197077 470870 200100 470872
rect 197077 470867 197143 470870
rect 358721 470658 358787 470661
rect 356132 470656 358787 470658
rect 356132 470600 358726 470656
rect 358782 470600 358787 470656
rect 356132 470598 358787 470600
rect 358721 470595 358787 470598
rect 83457 469842 83523 469845
rect 89662 469842 89668 469844
rect 83457 469840 89668 469842
rect 83457 469784 83462 469840
rect 83518 469784 89668 469840
rect 83457 469782 89668 469784
rect 83457 469779 83523 469782
rect 89662 469780 89668 469782
rect 89732 469780 89738 469844
rect 108389 469842 108455 469845
rect 117998 469842 118004 469844
rect 108389 469840 118004 469842
rect 108389 469784 108394 469840
rect 108450 469784 118004 469840
rect 108389 469782 118004 469784
rect 108389 469779 108455 469782
rect 117998 469780 118004 469782
rect 118068 469780 118074 469844
rect 90541 468482 90607 468485
rect 100702 468482 100708 468484
rect 90541 468480 100708 468482
rect 90541 468424 90546 468480
rect 90602 468424 100708 468480
rect 90541 468422 100708 468424
rect 90541 468419 90607 468422
rect 100702 468420 100708 468422
rect 100772 468420 100778 468484
rect 101397 468482 101463 468485
rect 115974 468482 115980 468484
rect 101397 468480 115980 468482
rect 101397 468424 101402 468480
rect 101458 468424 115980 468480
rect 101397 468422 115980 468424
rect 101397 468419 101463 468422
rect 115974 468420 115980 468422
rect 116044 468420 116050 468484
rect 197445 468482 197511 468485
rect 197445 468480 200100 468482
rect 197445 468424 197450 468480
rect 197506 468424 200100 468480
rect 197445 468422 200100 468424
rect 197445 468419 197511 468422
rect 356102 467938 356162 468180
rect 356237 467938 356303 467941
rect 356102 467936 356303 467938
rect 356102 467880 356242 467936
rect 356298 467880 356303 467936
rect 356102 467878 356303 467880
rect 356237 467875 356303 467878
rect 94589 467122 94655 467125
rect 108982 467122 108988 467124
rect 94589 467120 108988 467122
rect 94589 467064 94594 467120
rect 94650 467064 108988 467120
rect 94589 467062 108988 467064
rect 94589 467059 94655 467062
rect 108982 467060 108988 467062
rect 109052 467060 109058 467124
rect 197445 466034 197511 466037
rect 197445 466032 200100 466034
rect 197445 465976 197450 466032
rect 197506 465976 200100 466032
rect 197445 465974 200100 465976
rect 197445 465971 197511 465974
rect 86861 465762 86927 465765
rect 96654 465762 96660 465764
rect 86861 465760 96660 465762
rect 86861 465704 86866 465760
rect 86922 465704 96660 465760
rect 86861 465702 96660 465704
rect 86861 465699 86927 465702
rect 96654 465700 96660 465702
rect 96724 465700 96730 465764
rect 97257 465762 97323 465765
rect 107694 465762 107700 465764
rect 97257 465760 107700 465762
rect 97257 465704 97262 465760
rect 97318 465704 107700 465760
rect 97257 465702 107700 465704
rect 97257 465699 97323 465702
rect 107694 465700 107700 465702
rect 107764 465700 107770 465764
rect 358721 465762 358787 465765
rect 356132 465760 358787 465762
rect 356132 465704 358726 465760
rect 358782 465704 358787 465760
rect 356132 465702 358787 465704
rect 358721 465699 358787 465702
rect 156597 465220 156663 465221
rect 156597 465216 156644 465220
rect 156708 465218 156714 465220
rect 156597 465160 156602 465216
rect 156597 465156 156644 465160
rect 156708 465158 156754 465218
rect 156708 465156 156714 465158
rect 156597 465155 156663 465156
rect 197445 463314 197511 463317
rect 198825 463314 198891 463317
rect 358629 463314 358695 463317
rect 197445 463312 200100 463314
rect 197445 463256 197450 463312
rect 197506 463256 198830 463312
rect 198886 463256 200100 463312
rect 197445 463254 200100 463256
rect 356132 463312 358695 463314
rect 356132 463256 358634 463312
rect 358690 463256 358695 463312
rect 356132 463254 358695 463256
rect 197445 463251 197511 463254
rect 198825 463251 198891 463254
rect 358629 463251 358695 463254
rect 93117 462906 93183 462909
rect 102174 462906 102180 462908
rect 93117 462904 102180 462906
rect 93117 462848 93122 462904
rect 93178 462848 102180 462904
rect 93117 462846 102180 462848
rect 93117 462843 93183 462846
rect 102174 462844 102180 462846
rect 102244 462844 102250 462908
rect -960 462634 480 462724
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 197445 460866 197511 460869
rect 358721 460866 358787 460869
rect 197445 460864 200100 460866
rect 197445 460808 197450 460864
rect 197506 460808 200100 460864
rect 197445 460806 200100 460808
rect 356132 460864 358787 460866
rect 356132 460808 358726 460864
rect 358782 460808 358787 460864
rect 356132 460806 358787 460808
rect 197445 460803 197511 460806
rect 358721 460803 358787 460806
rect 81433 458962 81499 458965
rect 91134 458962 91140 458964
rect 81433 458960 91140 458962
rect 81433 458904 81438 458960
rect 81494 458904 91140 458960
rect 81433 458902 91140 458904
rect 81433 458899 81499 458902
rect 91134 458900 91140 458902
rect 91204 458900 91210 458964
rect 198774 458418 198780 458420
rect 180750 458358 198780 458418
rect 128997 458282 129063 458285
rect 180750 458282 180810 458358
rect 198774 458356 198780 458358
rect 198844 458418 198850 458420
rect 357433 458418 357499 458421
rect 198844 458358 200100 458418
rect 356132 458416 357499 458418
rect 356132 458360 357438 458416
rect 357494 458360 357499 458416
rect 356132 458358 357499 458360
rect 198844 458356 198850 458358
rect 357433 458355 357499 458358
rect 128997 458280 180810 458282
rect 128997 458224 129002 458280
rect 129058 458224 180810 458280
rect 128997 458222 180810 458224
rect 128997 458219 129063 458222
rect 582557 458146 582623 458149
rect 583109 458146 583175 458149
rect 583520 458146 584960 458236
rect 582557 458144 584960 458146
rect 582557 458088 582562 458144
rect 582618 458088 583114 458144
rect 583170 458088 584960 458144
rect 582557 458086 584960 458088
rect 582557 458083 582623 458086
rect 583109 458083 583175 458086
rect 583520 457996 584960 458086
rect 86953 457602 87019 457605
rect 98126 457602 98132 457604
rect 86953 457600 98132 457602
rect 86953 457544 86958 457600
rect 87014 457544 98132 457600
rect 86953 457542 98132 457544
rect 86953 457539 87019 457542
rect 98126 457540 98132 457542
rect 98196 457540 98202 457604
rect 97901 457466 97967 457469
rect 111742 457466 111748 457468
rect 97901 457464 111748 457466
rect 97901 457408 97906 457464
rect 97962 457408 111748 457464
rect 97901 457406 111748 457408
rect 97901 457403 97967 457406
rect 111742 457404 111748 457406
rect 111812 457404 111818 457468
rect 61837 456106 61903 456109
rect 71998 456106 72004 456108
rect 61837 456104 72004 456106
rect 61837 456048 61842 456104
rect 61898 456048 72004 456104
rect 61837 456046 72004 456048
rect 61837 456043 61903 456046
rect 71998 456044 72004 456046
rect 72068 456044 72074 456108
rect 82813 456106 82879 456109
rect 92606 456106 92612 456108
rect 82813 456104 92612 456106
rect 82813 456048 82818 456104
rect 82874 456048 92612 456104
rect 82813 456046 92612 456048
rect 82813 456043 82879 456046
rect 92606 456044 92612 456046
rect 92676 456044 92682 456108
rect 197445 455970 197511 455973
rect 358721 455970 358787 455973
rect 197445 455968 200100 455970
rect 197445 455912 197450 455968
rect 197506 455912 200100 455968
rect 197445 455910 200100 455912
rect 356132 455968 358787 455970
rect 356132 455912 358726 455968
rect 358782 455912 358787 455968
rect 356132 455910 358787 455912
rect 197445 455907 197511 455910
rect 358721 455907 358787 455910
rect 64689 454746 64755 454749
rect 72601 454746 72667 454749
rect 64689 454744 72667 454746
rect 64689 454688 64694 454744
rect 64750 454688 72606 454744
rect 72662 454688 72667 454744
rect 64689 454686 72667 454688
rect 64689 454683 64755 454686
rect 72601 454683 72667 454686
rect 198089 453522 198155 453525
rect 358721 453522 358787 453525
rect 198089 453520 200100 453522
rect 198089 453464 198094 453520
rect 198150 453464 200100 453520
rect 198089 453462 200100 453464
rect 356132 453520 358787 453522
rect 356132 453464 358726 453520
rect 358782 453464 358787 453520
rect 356132 453462 358787 453464
rect 198089 453459 198155 453462
rect 358721 453459 358787 453462
rect 66897 452570 66963 452573
rect 69054 452570 69060 452572
rect 66897 452568 69060 452570
rect 66897 452512 66902 452568
rect 66958 452512 69060 452568
rect 66897 452510 69060 452512
rect 66897 452507 66963 452510
rect 69054 452508 69060 452510
rect 69124 452508 69130 452572
rect 69054 451828 69060 451892
rect 69124 451890 69130 451892
rect 192661 451890 192727 451893
rect 69124 451888 192727 451890
rect 69124 451832 192666 451888
rect 192722 451832 192727 451888
rect 69124 451830 192727 451832
rect 69124 451828 69130 451830
rect 192661 451827 192727 451830
rect 358721 451074 358787 451077
rect 356132 451072 358787 451074
rect 98729 449986 98795 449989
rect 171869 449986 171935 449989
rect 98729 449984 171935 449986
rect 98729 449928 98734 449984
rect 98790 449928 171874 449984
rect 171930 449928 171935 449984
rect 98729 449926 171935 449928
rect 98729 449923 98795 449926
rect 171869 449923 171935 449926
rect 184790 449924 184796 449988
rect 184860 449986 184866 449988
rect 200070 449986 200130 451044
rect 356132 451016 358726 451072
rect 358782 451016 358787 451072
rect 356132 451014 358787 451016
rect 358721 451011 358787 451014
rect 184860 449926 200130 449986
rect 184860 449924 184866 449926
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 89069 449170 89135 449173
rect 93894 449170 93900 449172
rect 89069 449168 93900 449170
rect 89069 449112 89074 449168
rect 89130 449112 93900 449168
rect 89069 449110 93900 449112
rect 89069 449107 89135 449110
rect 93894 449108 93900 449110
rect 93964 449108 93970 449172
rect 111057 449170 111123 449173
rect 122598 449170 122604 449172
rect 111057 449168 122604 449170
rect 111057 449112 111062 449168
rect 111118 449112 122604 449168
rect 111057 449110 122604 449112
rect 111057 449107 111123 449110
rect 122598 449108 122604 449110
rect 122668 449108 122674 449172
rect 116117 448626 116183 448629
rect 155309 448626 155375 448629
rect 116117 448624 155375 448626
rect 116117 448568 116122 448624
rect 116178 448568 155314 448624
rect 155370 448568 155375 448624
rect 116117 448566 155375 448568
rect 116117 448563 116183 448566
rect 155309 448563 155375 448566
rect 197353 448626 197419 448629
rect 358721 448626 358787 448629
rect 197353 448624 200100 448626
rect 197353 448568 197358 448624
rect 197414 448568 200100 448624
rect 197353 448566 200100 448568
rect 356132 448624 358787 448626
rect 356132 448568 358726 448624
rect 358782 448568 358787 448624
rect 356132 448566 358787 448568
rect 197353 448563 197419 448566
rect 358721 448563 358787 448566
rect 57881 447810 57947 447813
rect 82813 447810 82879 447813
rect 57881 447808 82879 447810
rect 57881 447752 57886 447808
rect 57942 447752 82818 447808
rect 82874 447752 82879 447808
rect 57881 447750 82879 447752
rect 57881 447747 57947 447750
rect 82813 447747 82879 447750
rect 84193 447810 84259 447813
rect 95182 447810 95188 447812
rect 84193 447808 95188 447810
rect 84193 447752 84198 447808
rect 84254 447752 95188 447808
rect 84193 447750 95188 447752
rect 84193 447747 84259 447750
rect 95182 447748 95188 447750
rect 95252 447748 95258 447812
rect 105537 447130 105603 447133
rect 184841 447130 184907 447133
rect 186998 447130 187004 447132
rect 105537 447128 187004 447130
rect 105537 447072 105542 447128
rect 105598 447072 184846 447128
rect 184902 447072 187004 447128
rect 105537 447070 187004 447072
rect 105537 447067 105603 447070
rect 184841 447067 184907 447070
rect 186998 447068 187004 447070
rect 187068 447068 187074 447132
rect 92473 446994 92539 446997
rect 93025 446994 93091 446997
rect 130469 446994 130535 446997
rect 92473 446992 130535 446994
rect 92473 446936 92478 446992
rect 92534 446936 93030 446992
rect 93086 446936 130474 446992
rect 130530 446936 130535 446992
rect 92473 446934 130535 446936
rect 92473 446931 92539 446934
rect 93025 446931 93091 446934
rect 130469 446931 130535 446934
rect 70393 446450 70459 446453
rect 71814 446450 71820 446452
rect 70393 446448 71820 446450
rect 70393 446392 70398 446448
rect 70454 446392 71820 446448
rect 70393 446390 71820 446392
rect 70393 446387 70459 446390
rect 71814 446388 71820 446390
rect 71884 446388 71890 446452
rect 197353 446178 197419 446181
rect 358721 446178 358787 446181
rect 197353 446176 200100 446178
rect 197353 446120 197358 446176
rect 197414 446120 200100 446176
rect 197353 446118 200100 446120
rect 356132 446176 358787 446178
rect 356132 446120 358726 446176
rect 358782 446120 358787 446176
rect 356132 446118 358787 446120
rect 197353 446115 197419 446118
rect 358721 446115 358787 446118
rect 71773 445906 71839 445909
rect 71998 445906 72004 445908
rect 71773 445904 72004 445906
rect 71773 445848 71778 445904
rect 71834 445848 72004 445904
rect 71773 445846 72004 445848
rect 71773 445843 71839 445846
rect 71998 445844 72004 445846
rect 72068 445906 72074 445908
rect 72734 445906 72740 445908
rect 72068 445846 72740 445906
rect 72068 445844 72074 445846
rect 72734 445844 72740 445846
rect 72804 445844 72810 445908
rect 93710 445844 93716 445908
rect 93780 445906 93786 445908
rect 96613 445906 96679 445909
rect 97625 445906 97691 445909
rect 93780 445904 97691 445906
rect 93780 445848 96618 445904
rect 96674 445848 97630 445904
rect 97686 445848 97691 445904
rect 93780 445846 97691 445848
rect 93780 445844 93786 445846
rect 96613 445843 96679 445846
rect 97625 445843 97691 445846
rect 39941 445770 40007 445773
rect 93025 445770 93091 445773
rect 39941 445768 93091 445770
rect 39941 445712 39946 445768
rect 40002 445712 93030 445768
rect 93086 445712 93091 445768
rect 39941 445710 93091 445712
rect 39941 445707 40007 445710
rect 93025 445707 93091 445710
rect 100477 445772 100543 445773
rect 100477 445768 100524 445772
rect 100588 445770 100594 445772
rect 113173 445770 113239 445773
rect 114369 445772 114435 445773
rect 114318 445770 114324 445772
rect 100477 445712 100482 445768
rect 100477 445708 100524 445712
rect 100588 445710 100634 445770
rect 113173 445768 114324 445770
rect 114388 445768 114435 445772
rect 113173 445712 113178 445768
rect 113234 445712 114324 445768
rect 114430 445712 114435 445768
rect 113173 445710 114324 445712
rect 100588 445708 100594 445710
rect 100477 445707 100543 445708
rect 113173 445707 113239 445710
rect 114318 445708 114324 445710
rect 114388 445708 114435 445712
rect 114369 445707 114435 445708
rect 117589 445770 117655 445773
rect 118509 445772 118575 445773
rect 118509 445770 118556 445772
rect 117589 445768 118556 445770
rect 118620 445770 118626 445772
rect 168465 445770 168531 445773
rect 169017 445770 169083 445773
rect 117589 445712 117594 445768
rect 117650 445712 118514 445768
rect 117589 445710 118556 445712
rect 117589 445707 117655 445710
rect 118509 445708 118556 445710
rect 118620 445710 118702 445770
rect 168465 445768 169083 445770
rect 168465 445712 168470 445768
rect 168526 445712 169022 445768
rect 169078 445712 169083 445768
rect 168465 445710 169083 445712
rect 118620 445708 118626 445710
rect 118509 445707 118575 445708
rect 168465 445707 168531 445710
rect 169017 445707 169083 445710
rect 87597 444954 87663 444957
rect 87597 444952 103530 444954
rect 87597 444896 87602 444952
rect 87658 444896 103530 444952
rect 87597 444894 103530 444896
rect 87597 444891 87663 444894
rect 94497 444820 94563 444821
rect 94446 444818 94452 444820
rect 94406 444758 94452 444818
rect 94516 444816 94563 444820
rect 94558 444760 94563 444816
rect 94446 444756 94452 444758
rect 94516 444756 94563 444760
rect 103470 444818 103530 444894
rect 109534 444892 109540 444956
rect 109604 444954 109610 444956
rect 109677 444954 109743 444957
rect 109604 444952 109743 444954
rect 109604 444896 109682 444952
rect 109738 444896 109743 444952
rect 109604 444894 109743 444896
rect 109604 444892 109610 444894
rect 109677 444891 109743 444894
rect 111558 444892 111564 444956
rect 111628 444954 111634 444956
rect 111701 444954 111767 444957
rect 111628 444952 111767 444954
rect 111628 444896 111706 444952
rect 111762 444896 111767 444952
rect 111628 444894 111767 444896
rect 111628 444892 111634 444894
rect 111701 444891 111767 444894
rect 121545 444818 121611 444821
rect 103470 444816 121611 444818
rect 103470 444760 121550 444816
rect 121606 444760 121611 444816
rect 103470 444758 121611 444760
rect 94497 444755 94563 444756
rect 121545 444755 121611 444758
rect 90357 444682 90423 444685
rect 141417 444682 141483 444685
rect 90357 444680 141483 444682
rect 90357 444624 90362 444680
rect 90418 444624 141422 444680
rect 141478 444624 141483 444680
rect 583520 444668 584960 444908
rect 90357 444622 141483 444624
rect 90357 444619 90423 444622
rect 141417 444619 141483 444622
rect 55121 444546 55187 444549
rect 79409 444546 79475 444549
rect 55121 444544 79475 444546
rect 55121 444488 55126 444544
rect 55182 444488 79414 444544
rect 79470 444488 79475 444544
rect 55121 444486 79475 444488
rect 55121 444483 55187 444486
rect 79409 444483 79475 444486
rect 82813 444546 82879 444549
rect 83825 444546 83891 444549
rect 168465 444546 168531 444549
rect 82813 444544 168531 444546
rect 82813 444488 82818 444544
rect 82874 444488 83830 444544
rect 83886 444488 168470 444544
rect 168526 444488 168531 444544
rect 82813 444486 168531 444488
rect 82813 444483 82879 444486
rect 83825 444483 83891 444486
rect 168465 444483 168531 444486
rect 121545 444410 121611 444413
rect 122281 444410 122347 444413
rect 130377 444410 130443 444413
rect 121545 444408 130443 444410
rect 121545 444352 121550 444408
rect 121606 444352 122286 444408
rect 122342 444352 130382 444408
rect 130438 444352 130443 444408
rect 121545 444350 130443 444352
rect 121545 444347 121611 444350
rect 122281 444347 122347 444350
rect 130377 444347 130443 444350
rect 124121 444274 124187 444277
rect 120612 444272 124187 444274
rect 120612 444216 124126 444272
rect 124182 444216 124187 444272
rect 120612 444214 124187 444216
rect 124121 444211 124187 444214
rect 197353 443730 197419 443733
rect 358721 443730 358787 443733
rect 197353 443728 200100 443730
rect 197353 443672 197358 443728
rect 197414 443672 200100 443728
rect 197353 443670 200100 443672
rect 356132 443728 358787 443730
rect 356132 443672 358726 443728
rect 358782 443672 358787 443728
rect 356132 443670 358787 443672
rect 197353 443667 197419 443670
rect 358721 443667 358787 443670
rect 120901 442914 120967 442917
rect 120901 442912 122850 442914
rect 120901 442856 120906 442912
rect 120962 442856 122850 442912
rect 120901 442854 122850 442856
rect 120901 442851 120967 442854
rect 122790 442370 122850 442854
rect 154062 442370 154068 442372
rect 122790 442310 154068 442370
rect 154062 442308 154068 442310
rect 154132 442308 154138 442372
rect 67725 442234 67791 442237
rect 67725 442232 68908 442234
rect 67725 442176 67730 442232
rect 67786 442176 68908 442232
rect 67725 442174 68908 442176
rect 67725 442171 67791 442174
rect 124121 442098 124187 442101
rect 120612 442096 124187 442098
rect 120612 442040 124126 442096
rect 124182 442040 124187 442096
rect 120612 442038 124187 442040
rect 124121 442035 124187 442038
rect 197721 441418 197787 441421
rect 197721 441416 200100 441418
rect 197721 441360 197726 441416
rect 197782 441360 200100 441416
rect 197721 441358 200100 441360
rect 197721 441355 197787 441358
rect 359089 441282 359155 441285
rect 356132 441280 359155 441282
rect 356132 441224 359094 441280
rect 359150 441224 359155 441280
rect 356132 441222 359155 441224
rect 359089 441219 359155 441222
rect 66897 440058 66963 440061
rect 121453 440058 121519 440061
rect 66897 440056 68908 440058
rect 66897 440000 66902 440056
rect 66958 440000 68908 440056
rect 66897 439998 68908 440000
rect 120612 440056 121519 440058
rect 120612 440000 121458 440056
rect 121514 440000 121519 440056
rect 120612 439998 121519 440000
rect 66897 439995 66963 439998
rect 121453 439995 121519 439998
rect 196566 438908 196572 438972
rect 196636 438970 196642 438972
rect 357566 438970 357572 438972
rect 196636 438910 200100 438970
rect 356132 438910 357572 438970
rect 196636 438908 196642 438910
rect 357566 438908 357572 438910
rect 357636 438970 357642 438972
rect 358721 438970 358787 438973
rect 357636 438968 358787 438970
rect 357636 438912 358726 438968
rect 358782 438912 358787 438968
rect 357636 438910 358787 438912
rect 357636 438908 357642 438910
rect 358721 438907 358787 438910
rect 124121 437882 124187 437885
rect 120612 437880 124187 437882
rect 120612 437824 124126 437880
rect 124182 437824 124187 437880
rect 120612 437822 124187 437824
rect 124121 437819 124187 437822
rect 66897 437746 66963 437749
rect 66897 437744 68908 437746
rect 66897 437688 66902 437744
rect 66958 437688 68908 437744
rect 66897 437686 68908 437688
rect 66897 437683 66963 437686
rect -960 436508 480 436748
rect 197353 436386 197419 436389
rect 358721 436386 358787 436389
rect 197353 436384 200100 436386
rect 197353 436328 197358 436384
rect 197414 436328 200100 436384
rect 197353 436326 200100 436328
rect 356132 436384 358787 436386
rect 356132 436328 358726 436384
rect 358782 436328 358787 436384
rect 356132 436326 358787 436328
rect 197353 436323 197419 436326
rect 358721 436323 358787 436326
rect 120717 435978 120783 435981
rect 120582 435976 120783 435978
rect 120582 435920 120722 435976
rect 120778 435920 120783 435976
rect 120582 435918 120783 435920
rect 120582 435404 120642 435918
rect 120717 435915 120783 435918
rect 66897 435298 66963 435301
rect 66897 435296 68908 435298
rect 66897 435240 66902 435296
rect 66958 435240 68908 435296
rect 66897 435238 68908 435240
rect 66897 435235 66963 435238
rect 197353 433938 197419 433941
rect 358721 433938 358787 433941
rect 197353 433936 200100 433938
rect 197353 433880 197358 433936
rect 197414 433880 200100 433936
rect 197353 433878 200100 433880
rect 356132 433936 358787 433938
rect 356132 433880 358726 433936
rect 358782 433880 358787 433936
rect 356132 433878 358787 433880
rect 197353 433875 197419 433878
rect 358721 433875 358787 433878
rect 66805 433258 66871 433261
rect 124121 433258 124187 433261
rect 66805 433256 68908 433258
rect 66805 433200 66810 433256
rect 66866 433200 68908 433256
rect 66805 433198 68908 433200
rect 120612 433256 124187 433258
rect 120612 433200 124126 433256
rect 124182 433200 124187 433256
rect 120612 433198 124187 433200
rect 66805 433195 66871 433198
rect 124121 433195 124187 433198
rect 582373 431626 582439 431629
rect 583520 431626 584960 431716
rect 582373 431624 584960 431626
rect 582373 431568 582378 431624
rect 582434 431568 584960 431624
rect 582373 431566 584960 431568
rect 582373 431563 582439 431566
rect 358997 431490 359063 431493
rect 356132 431488 359063 431490
rect 66529 431082 66595 431085
rect 66529 431080 68908 431082
rect 66529 431024 66534 431080
rect 66590 431024 68908 431080
rect 66529 431022 68908 431024
rect 66529 431019 66595 431022
rect 120214 430674 120274 430916
rect 124121 430674 124187 430677
rect 120214 430672 124187 430674
rect 120214 430642 124126 430672
rect 120206 430578 120212 430642
rect 120276 430616 124126 430642
rect 124182 430616 124187 430672
rect 120276 430614 124187 430616
rect 120276 430578 120282 430614
rect 124121 430611 124187 430614
rect 177798 430612 177804 430676
rect 177868 430674 177874 430676
rect 200070 430674 200130 431460
rect 356132 431432 359002 431488
rect 359058 431432 359063 431488
rect 583520 431476 584960 431566
rect 356132 431430 359063 431432
rect 358997 431427 359063 431430
rect 177868 430614 200130 430674
rect 177868 430612 177874 430614
rect 197353 429042 197419 429045
rect 358721 429042 358787 429045
rect 197353 429040 200100 429042
rect 197353 428984 197358 429040
rect 197414 428984 200100 429040
rect 197353 428982 200100 428984
rect 356132 429040 358787 429042
rect 356132 428984 358726 429040
rect 358782 428984 358787 429040
rect 356132 428982 358787 428984
rect 197353 428979 197419 428982
rect 358721 428979 358787 428982
rect 120390 428708 120396 428772
rect 120460 428708 120466 428772
rect 66713 428634 66779 428637
rect 66713 428632 68908 428634
rect 66713 428576 66718 428632
rect 66774 428576 68908 428632
rect 66713 428574 68908 428576
rect 66713 428571 66779 428574
rect 120398 428498 120458 428708
rect 121453 428498 121519 428501
rect 120398 428496 121519 428498
rect 120398 428468 121458 428496
rect 120428 428440 121458 428468
rect 121514 428440 121519 428496
rect 120428 428438 121519 428440
rect 121453 428435 121519 428438
rect 197353 426594 197419 426597
rect 358721 426594 358787 426597
rect 197353 426592 200100 426594
rect 197353 426536 197358 426592
rect 197414 426536 200100 426592
rect 197353 426534 200100 426536
rect 356132 426592 358787 426594
rect 356132 426536 358726 426592
rect 358782 426536 358787 426592
rect 356132 426534 358787 426536
rect 197353 426531 197419 426534
rect 358721 426531 358787 426534
rect 66253 426322 66319 426325
rect 121678 426322 121684 426324
rect 66253 426320 68908 426322
rect 66253 426264 66258 426320
rect 66314 426264 68908 426320
rect 66253 426262 68908 426264
rect 120612 426262 121684 426322
rect 66253 426259 66319 426262
rect 121678 426260 121684 426262
rect 121748 426322 121754 426324
rect 122598 426322 122604 426324
rect 121748 426262 122604 426322
rect 121748 426260 121754 426262
rect 122598 426260 122604 426262
rect 122668 426260 122674 426324
rect 66069 424282 66135 424285
rect 66069 424280 68908 424282
rect 66069 424224 66074 424280
rect 66130 424224 68908 424280
rect 66069 424222 68908 424224
rect 66069 424219 66135 424222
rect 197353 424146 197419 424149
rect 197353 424144 200100 424146
rect 120582 423738 120642 424116
rect 197353 424088 197358 424144
rect 197414 424088 200100 424144
rect 197353 424086 200100 424088
rect 197353 424083 197419 424086
rect 122833 423738 122899 423741
rect 123477 423738 123543 423741
rect 120582 423736 123543 423738
rect -960 423602 480 423692
rect 120582 423680 122838 423736
rect 122894 423680 123482 423736
rect 123538 423680 123543 423736
rect 120582 423678 123543 423680
rect 356102 423738 356162 424116
rect 356237 423738 356303 423741
rect 356102 423736 356303 423738
rect 356102 423680 356242 423736
rect 356298 423680 356303 423736
rect 356102 423678 356303 423680
rect 122833 423675 122899 423678
rect 123477 423675 123543 423678
rect 356237 423675 356303 423678
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 124121 422106 124187 422109
rect 120612 422104 124187 422106
rect 120612 422048 124126 422104
rect 124182 422048 124187 422104
rect 120612 422046 124187 422048
rect 124121 422043 124187 422046
rect 66253 421970 66319 421973
rect 66253 421968 68908 421970
rect 66253 421912 66258 421968
rect 66314 421912 68908 421968
rect 66253 421910 68908 421912
rect 66253 421907 66319 421910
rect 198641 421698 198707 421701
rect 357525 421698 357591 421701
rect 198641 421696 200100 421698
rect 198641 421640 198646 421696
rect 198702 421640 200100 421696
rect 198641 421638 200100 421640
rect 356132 421696 357591 421698
rect 356132 421640 357530 421696
rect 357586 421640 357591 421696
rect 356132 421638 357591 421640
rect 198641 421635 198707 421638
rect 357525 421635 357591 421638
rect 66662 419596 66668 419660
rect 66732 419658 66738 419660
rect 67766 419658 67772 419660
rect 66732 419598 67772 419658
rect 66732 419596 66738 419598
rect 67766 419596 67772 419598
rect 67836 419658 67842 419660
rect 121494 419658 121500 419660
rect 67836 419598 68908 419658
rect 120612 419598 121500 419658
rect 67836 419596 67842 419598
rect 121494 419596 121500 419598
rect 121564 419658 121570 419660
rect 123017 419658 123083 419661
rect 121564 419656 123083 419658
rect 121564 419600 123022 419656
rect 123078 419600 123083 419656
rect 121564 419598 123083 419600
rect 121564 419596 121570 419598
rect 123017 419595 123083 419598
rect 197353 419250 197419 419253
rect 358721 419250 358787 419253
rect 197353 419248 200100 419250
rect 197353 419192 197358 419248
rect 197414 419192 200100 419248
rect 197353 419190 200100 419192
rect 356132 419248 358787 419250
rect 356132 419192 358726 419248
rect 358782 419192 358787 419248
rect 356132 419190 358787 419192
rect 197353 419187 197419 419190
rect 358721 419187 358787 419190
rect 583293 418298 583359 418301
rect 583520 418298 584960 418388
rect 583293 418296 584960 418298
rect 583293 418240 583298 418296
rect 583354 418240 584960 418296
rect 583293 418238 584960 418240
rect 583293 418235 583359 418238
rect 583520 418148 584960 418238
rect 122189 418026 122255 418029
rect 120582 418024 122255 418026
rect 120582 417968 122194 418024
rect 122250 417968 122255 418024
rect 120582 417966 122255 417968
rect 66897 417346 66963 417349
rect 66897 417344 68908 417346
rect 66897 417288 66902 417344
rect 66958 417288 68908 417344
rect 66897 417286 68908 417288
rect 66897 417283 66963 417286
rect 120582 417074 120642 417966
rect 122189 417963 122255 417966
rect 120717 417074 120783 417077
rect 120582 417072 120783 417074
rect 120582 417016 120722 417072
rect 120778 417016 120783 417072
rect 120582 417014 120783 417016
rect 120717 417011 120783 417014
rect 198917 416802 198983 416805
rect 358721 416802 358787 416805
rect 198917 416800 200100 416802
rect 198917 416744 198922 416800
rect 198978 416744 200100 416800
rect 198917 416742 200100 416744
rect 356132 416800 358787 416802
rect 356132 416744 358726 416800
rect 358782 416744 358787 416800
rect 356132 416742 358787 416744
rect 198917 416739 198983 416742
rect 358721 416739 358787 416742
rect 66253 415170 66319 415173
rect 124121 415170 124187 415173
rect 66253 415168 68908 415170
rect 66253 415112 66258 415168
rect 66314 415112 68908 415168
rect 66253 415110 68908 415112
rect 120612 415168 124187 415170
rect 120612 415112 124126 415168
rect 124182 415112 124187 415168
rect 120612 415110 124187 415112
rect 66253 415107 66319 415110
rect 124121 415107 124187 415110
rect 197353 414354 197419 414357
rect 358721 414354 358787 414357
rect 197353 414352 200100 414354
rect 197353 414296 197358 414352
rect 197414 414296 200100 414352
rect 197353 414294 200100 414296
rect 356132 414352 358787 414354
rect 356132 414296 358726 414352
rect 358782 414296 358787 414352
rect 356132 414294 358787 414296
rect 197353 414291 197419 414294
rect 358721 414291 358787 414294
rect 67449 412858 67515 412861
rect 122833 412858 122899 412861
rect 67449 412856 68908 412858
rect 67449 412800 67454 412856
rect 67510 412800 68908 412856
rect 67449 412798 68908 412800
rect 120612 412856 122899 412858
rect 120612 412800 122838 412856
rect 122894 412800 122899 412856
rect 120612 412798 122899 412800
rect 67449 412795 67515 412798
rect 122833 412795 122899 412798
rect 197353 411906 197419 411909
rect 358721 411906 358787 411909
rect 197353 411904 200100 411906
rect 197353 411848 197358 411904
rect 197414 411848 200100 411904
rect 197353 411846 200100 411848
rect 356132 411904 358787 411906
rect 356132 411848 358726 411904
rect 358782 411848 358787 411904
rect 356132 411846 358787 411848
rect 197353 411843 197419 411846
rect 358721 411843 358787 411846
rect 120625 411090 120691 411093
rect 120582 411088 120691 411090
rect 120582 411032 120630 411088
rect 120686 411032 120691 411088
rect 120582 411027 120691 411032
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 67357 410546 67423 410549
rect 120582 410546 120642 411027
rect 121177 410546 121243 410549
rect 67357 410544 69092 410546
rect 67357 410488 67362 410544
rect 67418 410516 69092 410544
rect 120582 410544 121243 410546
rect 120582 410516 121182 410544
rect 67418 410488 69122 410516
rect 67357 410486 69122 410488
rect 120612 410488 121182 410516
rect 121238 410488 121243 410544
rect 120612 410486 121243 410488
rect 67357 410483 67423 410486
rect 69062 410004 69122 410486
rect 121177 410483 121243 410486
rect 69054 409940 69060 410004
rect 69124 409940 69130 410004
rect 197353 409594 197419 409597
rect 197353 409592 200100 409594
rect 197353 409536 197358 409592
rect 197414 409536 200100 409592
rect 197353 409534 200100 409536
rect 197353 409531 197419 409534
rect 358854 409458 358860 409460
rect 356132 409398 358860 409458
rect 358854 409396 358860 409398
rect 358924 409396 358930 409460
rect 124121 408506 124187 408509
rect 120612 408504 124187 408506
rect 120612 408448 124126 408504
rect 124182 408448 124187 408504
rect 120612 408446 124187 408448
rect 124121 408443 124187 408446
rect 66345 408370 66411 408373
rect 66345 408368 68908 408370
rect 66345 408312 66350 408368
rect 66406 408312 68908 408368
rect 66345 408310 68908 408312
rect 66345 408307 66411 408310
rect 197353 407010 197419 407013
rect 358721 407010 358787 407013
rect 197353 407008 200100 407010
rect 197353 406952 197358 407008
rect 197414 406952 200100 407008
rect 197353 406950 200100 406952
rect 356132 407008 358787 407010
rect 356132 406952 358726 407008
rect 358782 406952 358787 407008
rect 356132 406950 358787 406952
rect 197353 406947 197419 406950
rect 358721 406947 358787 406950
rect 124305 406330 124371 406333
rect 120612 406328 124371 406330
rect 120612 406272 124310 406328
rect 124366 406272 124371 406328
rect 120612 406270 124371 406272
rect 124305 406267 124371 406270
rect 66805 406194 66871 406197
rect 66805 406192 68908 406194
rect 66805 406136 66810 406192
rect 66866 406136 68908 406192
rect 66805 406134 68908 406136
rect 66805 406131 66871 406134
rect 582649 404970 582715 404973
rect 582925 404970 582991 404973
rect 583520 404970 584960 405060
rect 582649 404968 584960 404970
rect 582649 404912 582654 404968
rect 582710 404912 582930 404968
rect 582986 404912 584960 404968
rect 582649 404910 584960 404912
rect 582649 404907 582715 404910
rect 582925 404907 582991 404910
rect 583520 404820 584960 404910
rect 197353 404562 197419 404565
rect 197353 404560 200100 404562
rect 197353 404504 197358 404560
rect 197414 404504 200100 404560
rect 197353 404502 200100 404504
rect 197353 404499 197419 404502
rect 358721 404290 358787 404293
rect 356132 404288 358787 404290
rect 356132 404232 358726 404288
rect 358782 404232 358787 404288
rect 356132 404230 358787 404232
rect 358721 404227 358787 404230
rect 66621 403746 66687 403749
rect 122925 403746 122991 403749
rect 66621 403744 68908 403746
rect 66621 403688 66626 403744
rect 66682 403688 68908 403744
rect 66621 403686 68908 403688
rect 120612 403744 122991 403746
rect 120612 403688 122930 403744
rect 122986 403688 122991 403744
rect 120612 403686 122991 403688
rect 66621 403683 66687 403686
rect 122925 403683 122991 403686
rect 173014 401644 173020 401708
rect 173084 401706 173090 401708
rect 200070 401706 200130 402084
rect 358721 401842 358787 401845
rect 356132 401840 358787 401842
rect 356132 401784 358726 401840
rect 358782 401784 358787 401840
rect 356132 401782 358787 401784
rect 358721 401779 358787 401782
rect 173084 401646 200130 401706
rect 173084 401644 173090 401646
rect 66805 401570 66871 401573
rect 123937 401570 124003 401573
rect 66805 401568 68908 401570
rect 66805 401512 66810 401568
rect 66866 401512 68908 401568
rect 66805 401510 68908 401512
rect 120612 401568 124003 401570
rect 120612 401512 123942 401568
rect 123998 401512 124003 401568
rect 120612 401510 124003 401512
rect 66805 401507 66871 401510
rect 123937 401507 124003 401510
rect 197353 399666 197419 399669
rect 197353 399664 200100 399666
rect 197353 399608 197358 399664
rect 197414 399608 200100 399664
rect 197353 399606 200100 399608
rect 197353 399603 197419 399606
rect 66805 399530 66871 399533
rect 124121 399530 124187 399533
rect 66805 399528 68908 399530
rect 66805 399472 66810 399528
rect 66866 399472 68908 399528
rect 66805 399470 68908 399472
rect 120612 399528 124187 399530
rect 120612 399472 124126 399528
rect 124182 399472 124187 399528
rect 120612 399470 124187 399472
rect 66805 399467 66871 399470
rect 124121 399467 124187 399470
rect 358629 399394 358695 399397
rect 356132 399392 358695 399394
rect 356132 399336 358634 399392
rect 358690 399336 358695 399392
rect 356132 399334 358695 399336
rect 358629 399331 358695 399334
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 66989 396946 67055 396949
rect 67357 396946 67423 396949
rect 124121 396946 124187 396949
rect 66989 396944 68908 396946
rect 66989 396888 66994 396944
rect 67050 396888 67362 396944
rect 67418 396888 68908 396944
rect 66989 396886 68908 396888
rect 120612 396944 124187 396946
rect 120612 396888 124126 396944
rect 124182 396888 124187 396944
rect 120612 396886 124187 396888
rect 66989 396883 67055 396886
rect 67357 396883 67423 396886
rect 124121 396883 124187 396886
rect 173198 396068 173204 396132
rect 173268 396130 173274 396132
rect 200070 396130 200130 397188
rect 360326 396946 360332 396948
rect 356132 396886 360332 396946
rect 360326 396884 360332 396886
rect 360396 396884 360402 396948
rect 173268 396070 200130 396130
rect 173268 396068 173274 396070
rect 67265 395994 67331 395997
rect 67541 395994 67607 395997
rect 67265 395992 67607 395994
rect 67265 395936 67270 395992
rect 67326 395936 67546 395992
rect 67602 395936 67607 395992
rect 67265 395934 67607 395936
rect 67265 395931 67331 395934
rect 67541 395931 67607 395934
rect 67541 394906 67607 394909
rect 67541 394904 68908 394906
rect 67541 394848 67546 394904
rect 67602 394848 68908 394904
rect 67541 394846 68908 394848
rect 67541 394843 67607 394846
rect 122782 394770 122788 394772
rect 120612 394710 122788 394770
rect 122782 394708 122788 394710
rect 122852 394708 122858 394772
rect 197353 394770 197419 394773
rect 197353 394768 200100 394770
rect 197353 394712 197358 394768
rect 197414 394712 200100 394768
rect 197353 394710 200100 394712
rect 197353 394707 197419 394710
rect 356329 394498 356395 394501
rect 356132 394496 356395 394498
rect 356132 394440 356334 394496
rect 356390 394440 356395 394496
rect 356132 394438 356395 394440
rect 356329 394435 356395 394438
rect 65793 393274 65859 393277
rect 65926 393274 65932 393276
rect 65793 393272 65932 393274
rect 65793 393216 65798 393272
rect 65854 393216 65932 393272
rect 65793 393214 65932 393216
rect 65793 393211 65859 393214
rect 65926 393212 65932 393214
rect 65996 393274 66002 393276
rect 65996 393214 68938 393274
rect 65996 393212 66002 393214
rect 68878 392700 68938 393214
rect 122925 392594 122991 392597
rect 123753 392594 123819 392597
rect 120612 392592 123819 392594
rect 120612 392536 122930 392592
rect 122986 392536 123758 392592
rect 123814 392536 123819 392592
rect 120612 392534 123819 392536
rect 122925 392531 122991 392534
rect 123753 392531 123819 392534
rect 198549 392322 198615 392325
rect 180750 392320 200100 392322
rect 180750 392264 198554 392320
rect 198610 392264 200100 392320
rect 180750 392262 200100 392264
rect 119470 392124 119476 392188
rect 119540 392186 119546 392188
rect 180750 392186 180810 392262
rect 198549 392259 198615 392262
rect 119540 392126 180810 392186
rect 119540 392124 119546 392126
rect 357617 392050 357683 392053
rect 356132 392048 357683 392050
rect 356132 391992 357622 392048
rect 357678 391992 357683 392048
rect 356132 391990 357683 391992
rect 357617 391987 357683 391990
rect 583520 391628 584960 391868
rect 61745 391370 61811 391373
rect 80462 391370 80468 391372
rect 61745 391368 80468 391370
rect 61745 391312 61750 391368
rect 61806 391312 80468 391368
rect 61745 391310 80468 391312
rect 61745 391307 61811 391310
rect 80462 391308 80468 391310
rect 80532 391308 80538 391372
rect 63217 391234 63283 391237
rect 142797 391234 142863 391237
rect 63217 391232 64890 391234
rect 63217 391176 63222 391232
rect 63278 391176 64890 391232
rect 63217 391174 64890 391176
rect 63217 391171 63283 391174
rect 64830 391098 64890 391174
rect 93810 391232 142863 391234
rect 93810 391176 142802 391232
rect 142858 391176 142863 391232
rect 93810 391174 142863 391176
rect 85849 391098 85915 391101
rect 93810 391098 93870 391174
rect 142797 391171 142863 391174
rect 64830 391096 93870 391098
rect 64830 391040 85854 391096
rect 85910 391040 93870 391096
rect 64830 391038 93870 391040
rect 85849 391035 85915 391038
rect 104934 391036 104940 391100
rect 105004 391098 105010 391100
rect 105077 391098 105143 391101
rect 105004 391096 105143 391098
rect 105004 391040 105082 391096
rect 105138 391040 105143 391096
rect 105004 391038 105143 391040
rect 105004 391036 105010 391038
rect 105077 391035 105143 391038
rect 80053 390962 80119 390965
rect 80462 390962 80468 390964
rect 80053 390960 80468 390962
rect 80053 390904 80058 390960
rect 80114 390904 80468 390960
rect 80053 390902 80468 390904
rect 80053 390899 80119 390902
rect 80462 390900 80468 390902
rect 80532 390962 80538 390964
rect 80605 390962 80671 390965
rect 80532 390960 80671 390962
rect 80532 390904 80610 390960
rect 80666 390904 80671 390960
rect 80532 390902 80671 390904
rect 80532 390900 80538 390902
rect 80605 390899 80671 390902
rect 115749 390690 115815 390693
rect 121494 390690 121500 390692
rect 115749 390688 121500 390690
rect 115749 390632 115754 390688
rect 115810 390632 121500 390688
rect 115749 390630 121500 390632
rect 115749 390627 115815 390630
rect 121494 390628 121500 390630
rect 121564 390628 121570 390692
rect 71865 390556 71931 390557
rect 71814 390554 71820 390556
rect 71774 390494 71820 390554
rect 71884 390552 71931 390556
rect 71926 390496 71931 390552
rect 71814 390492 71820 390494
rect 71884 390492 71931 390496
rect 108982 390492 108988 390556
rect 109052 390554 109058 390556
rect 109677 390554 109743 390557
rect 109052 390552 109743 390554
rect 109052 390496 109682 390552
rect 109738 390496 109743 390552
rect 109052 390494 109743 390496
rect 109052 390492 109058 390494
rect 71865 390491 71931 390492
rect 109677 390491 109743 390494
rect 69606 390356 69612 390420
rect 69676 390418 69682 390420
rect 69933 390418 69999 390421
rect 69676 390416 69999 390418
rect 69676 390360 69938 390416
rect 69994 390360 69999 390416
rect 69676 390358 69999 390360
rect 69676 390356 69682 390358
rect 69933 390355 69999 390358
rect 89662 390356 89668 390420
rect 89732 390418 89738 390420
rect 89805 390418 89871 390421
rect 89732 390416 89871 390418
rect 89732 390360 89810 390416
rect 89866 390360 89871 390416
rect 89732 390358 89871 390360
rect 89732 390356 89738 390358
rect 89805 390355 89871 390358
rect 91134 390356 91140 390420
rect 91204 390418 91210 390420
rect 91277 390418 91343 390421
rect 91204 390416 91343 390418
rect 91204 390360 91282 390416
rect 91338 390360 91343 390416
rect 91204 390358 91343 390360
rect 91204 390356 91210 390358
rect 91277 390355 91343 390358
rect 92606 390356 92612 390420
rect 92676 390418 92682 390420
rect 92749 390418 92815 390421
rect 92676 390416 92815 390418
rect 92676 390360 92754 390416
rect 92810 390360 92815 390416
rect 92676 390358 92815 390360
rect 92676 390356 92682 390358
rect 92749 390355 92815 390358
rect 93894 390356 93900 390420
rect 93964 390418 93970 390420
rect 94221 390418 94287 390421
rect 93964 390416 94287 390418
rect 93964 390360 94226 390416
rect 94282 390360 94287 390416
rect 93964 390358 94287 390360
rect 93964 390356 93970 390358
rect 94221 390355 94287 390358
rect 95366 390356 95372 390420
rect 95436 390418 95442 390420
rect 95877 390418 95943 390421
rect 95436 390416 95943 390418
rect 95436 390360 95882 390416
rect 95938 390360 95943 390416
rect 95436 390358 95943 390360
rect 95436 390356 95442 390358
rect 95877 390355 95943 390358
rect 96654 390356 96660 390420
rect 96724 390418 96730 390420
rect 97349 390418 97415 390421
rect 96724 390416 97415 390418
rect 96724 390360 97354 390416
rect 97410 390360 97415 390416
rect 96724 390358 97415 390360
rect 96724 390356 96730 390358
rect 97349 390355 97415 390358
rect 98126 390356 98132 390420
rect 98196 390418 98202 390420
rect 98821 390418 98887 390421
rect 98196 390416 98887 390418
rect 98196 390360 98826 390416
rect 98882 390360 98887 390416
rect 98196 390358 98887 390360
rect 98196 390356 98202 390358
rect 98821 390355 98887 390358
rect 100661 390420 100727 390421
rect 102133 390420 102199 390421
rect 100661 390416 100708 390420
rect 100772 390418 100778 390420
rect 100661 390360 100666 390416
rect 100661 390356 100708 390360
rect 100772 390358 100818 390418
rect 102133 390416 102180 390420
rect 102244 390418 102250 390420
rect 102133 390360 102138 390416
rect 100772 390356 100778 390358
rect 102133 390356 102180 390360
rect 102244 390358 102290 390418
rect 102244 390356 102250 390358
rect 106406 390356 106412 390420
rect 106476 390418 106482 390420
rect 106549 390418 106615 390421
rect 106476 390416 106615 390418
rect 106476 390360 106554 390416
rect 106610 390360 106615 390416
rect 106476 390358 106615 390360
rect 106476 390356 106482 390358
rect 100661 390355 100727 390356
rect 102133 390355 102199 390356
rect 106549 390355 106615 390358
rect 107694 390356 107700 390420
rect 107764 390418 107770 390420
rect 108021 390418 108087 390421
rect 107764 390416 108087 390418
rect 107764 390360 108026 390416
rect 108082 390360 108087 390416
rect 107764 390358 108087 390360
rect 107764 390356 107770 390358
rect 108021 390355 108087 390358
rect 115933 390420 115999 390421
rect 115933 390416 115980 390420
rect 116044 390418 116050 390420
rect 117865 390418 117931 390421
rect 117998 390418 118004 390420
rect 115933 390360 115938 390416
rect 115933 390356 115980 390360
rect 116044 390358 116090 390418
rect 117865 390416 118004 390418
rect 117865 390360 117870 390416
rect 117926 390360 118004 390416
rect 117865 390358 118004 390360
rect 116044 390356 116050 390358
rect 115933 390355 115999 390356
rect 117865 390355 117931 390358
rect 117998 390356 118004 390358
rect 118068 390356 118074 390420
rect 68553 390282 68619 390285
rect 76414 390282 76420 390284
rect 68553 390280 76420 390282
rect 68553 390224 68558 390280
rect 68614 390224 76420 390280
rect 68553 390222 76420 390224
rect 68553 390219 68619 390222
rect 76414 390220 76420 390222
rect 76484 390220 76490 390284
rect 197353 390010 197419 390013
rect 197353 390008 200100 390010
rect 197353 389952 197358 390008
rect 197414 389952 200100 390008
rect 197353 389950 200100 389952
rect 197353 389947 197419 389950
rect 357709 389602 357775 389605
rect 356132 389600 357775 389602
rect 356132 389544 357714 389600
rect 357770 389544 357775 389600
rect 356132 389542 357775 389544
rect 357709 389539 357775 389542
rect 3417 389194 3483 389197
rect 89662 389194 89668 389196
rect 3417 389192 89668 389194
rect 3417 389136 3422 389192
rect 3478 389136 89668 389192
rect 3417 389134 89668 389136
rect 3417 389131 3483 389134
rect 89662 389132 89668 389134
rect 89732 389132 89738 389196
rect 109769 389194 109835 389197
rect 166257 389194 166323 389197
rect 109769 389192 166323 389194
rect 109769 389136 109774 389192
rect 109830 389136 166262 389192
rect 166318 389136 166323 389192
rect 109769 389134 166323 389136
rect 109769 389131 109835 389134
rect 166257 389131 166323 389134
rect 100845 389058 100911 389061
rect 101857 389058 101923 389061
rect 100845 389056 101923 389058
rect 100845 389000 100850 389056
rect 100906 389000 101862 389056
rect 101918 389000 101923 389056
rect 100845 388998 101923 389000
rect 100845 388995 100911 388998
rect 101857 388995 101923 388998
rect 102317 389058 102383 389061
rect 103329 389058 103395 389061
rect 102317 389056 103395 389058
rect 102317 389000 102322 389056
rect 102378 389000 103334 389056
rect 103390 389000 103395 389056
rect 102317 388998 103395 389000
rect 102317 388995 102383 388998
rect 103329 388995 103395 388998
rect 111742 388996 111748 389060
rect 111812 389058 111818 389060
rect 112897 389058 112963 389061
rect 111812 389056 112963 389058
rect 111812 389000 112902 389056
rect 112958 389000 112963 389056
rect 111812 388998 112963 389000
rect 111812 388996 111818 388998
rect 112897 388995 112963 388998
rect 116117 389058 116183 389061
rect 117129 389058 117195 389061
rect 116117 389056 117195 389058
rect 116117 389000 116122 389056
rect 116178 389000 117134 389056
rect 117190 389000 117195 389056
rect 116117 388998 117195 389000
rect 116117 388995 116183 388998
rect 117129 388995 117195 388998
rect 64689 388922 64755 388925
rect 74533 388922 74599 388925
rect 64689 388920 74599 388922
rect 64689 388864 64694 388920
rect 64750 388864 74538 388920
rect 74594 388864 74599 388920
rect 64689 388862 74599 388864
rect 64689 388859 64755 388862
rect 74533 388859 74599 388862
rect 99966 388860 99972 388924
rect 100036 388922 100042 388924
rect 103697 388922 103763 388925
rect 100036 388920 103763 388922
rect 100036 388864 103702 388920
rect 103758 388864 103763 388920
rect 100036 388862 103763 388864
rect 100036 388860 100042 388862
rect 103697 388859 103763 388862
rect 115054 388860 115060 388924
rect 115124 388922 115130 388924
rect 117313 388922 117379 388925
rect 118969 388922 119035 388925
rect 115124 388920 119035 388922
rect 115124 388864 117318 388920
rect 117374 388864 118974 388920
rect 119030 388864 119035 388920
rect 115124 388862 119035 388864
rect 115124 388860 115130 388862
rect 117313 388859 117379 388862
rect 118969 388859 119035 388862
rect 83917 388788 83983 388789
rect 83917 388786 83964 388788
rect 83836 388784 83964 388786
rect 84028 388786 84034 388788
rect 135253 388786 135319 388789
rect 84028 388784 135319 388786
rect 83836 388728 83922 388784
rect 84028 388728 135258 388784
rect 135314 388728 135319 388784
rect 83836 388726 83964 388728
rect 83917 388724 83964 388726
rect 84028 388726 135319 388728
rect 84028 388724 84034 388726
rect 83917 388723 83983 388724
rect 135253 388723 135319 388726
rect 95182 387772 95188 387836
rect 95252 387834 95258 387836
rect 96245 387834 96311 387837
rect 95252 387832 96311 387834
rect 95252 387776 96250 387832
rect 96306 387776 96311 387832
rect 95252 387774 96311 387776
rect 95252 387772 95258 387774
rect 96245 387771 96311 387774
rect 100477 387836 100543 387837
rect 100477 387832 100524 387836
rect 100588 387834 100594 387836
rect 100477 387776 100482 387832
rect 100477 387772 100524 387776
rect 100588 387774 100634 387834
rect 100588 387772 100594 387774
rect 100477 387771 100543 387772
rect 66161 387698 66227 387701
rect 79317 387698 79383 387701
rect 66161 387696 79383 387698
rect 66161 387640 66166 387696
rect 66222 387640 79322 387696
rect 79378 387640 79383 387696
rect 66161 387638 79383 387640
rect 66161 387635 66227 387638
rect 79317 387635 79383 387638
rect 197353 387426 197419 387429
rect 197353 387424 200100 387426
rect 197353 387368 197358 387424
rect 197414 387368 200100 387424
rect 197353 387366 200100 387368
rect 197353 387363 197419 387366
rect 356421 387154 356487 387157
rect 356132 387152 356487 387154
rect 356132 387096 356426 387152
rect 356482 387096 356487 387152
rect 356132 387094 356487 387096
rect 356421 387091 356487 387094
rect 97717 387018 97783 387021
rect 158069 387018 158135 387021
rect 97717 387016 158135 387018
rect 97717 386960 97722 387016
rect 97778 386960 158074 387016
rect 158130 386960 158135 387016
rect 97717 386958 158135 386960
rect 97717 386955 97783 386958
rect 158069 386955 158135 386958
rect 105537 386474 105603 386477
rect 192334 386474 192340 386476
rect 105537 386472 192340 386474
rect 105537 386416 105542 386472
rect 105598 386416 192340 386472
rect 105537 386414 192340 386416
rect 105537 386411 105603 386414
rect 192334 386412 192340 386414
rect 192404 386412 192410 386476
rect 113173 386338 113239 386341
rect 114369 386338 114435 386341
rect 124213 386338 124279 386341
rect 113173 386336 124279 386338
rect 113173 386280 113178 386336
rect 113234 386280 114374 386336
rect 114430 386280 124218 386336
rect 124274 386280 124279 386336
rect 113173 386278 124279 386280
rect 113173 386275 113239 386278
rect 114369 386275 114435 386278
rect 124213 386275 124279 386278
rect 91645 385794 91711 385797
rect 119981 385794 120047 385797
rect 91645 385792 120047 385794
rect 91645 385736 91650 385792
rect 91706 385736 119986 385792
rect 120042 385736 120047 385792
rect 91645 385734 120047 385736
rect 91645 385731 91711 385734
rect 119981 385731 120047 385734
rect 4797 385658 4863 385661
rect 95182 385658 95188 385660
rect 4797 385656 95188 385658
rect 4797 385600 4802 385656
rect 4858 385600 95188 385656
rect 4797 385598 95188 385600
rect 4797 385595 4863 385598
rect 95182 385596 95188 385598
rect 95252 385596 95258 385660
rect 104157 385658 104223 385661
rect 134517 385658 134583 385661
rect 104157 385656 134583 385658
rect 104157 385600 104162 385656
rect 104218 385600 134522 385656
rect 134578 385600 134583 385656
rect 104157 385598 134583 385600
rect 104157 385595 104223 385598
rect 134517 385595 134583 385598
rect 197353 385114 197419 385117
rect 198590 385114 198596 385116
rect 197353 385112 198596 385114
rect 197353 385056 197358 385112
rect 197414 385056 198596 385112
rect 197353 385054 198596 385056
rect 197353 385051 197419 385054
rect 198590 385052 198596 385054
rect 198660 385052 198666 385116
rect 196709 384978 196775 384981
rect 196709 384976 200100 384978
rect 196709 384920 196714 384976
rect 196770 384920 200100 384976
rect 196709 384918 200100 384920
rect 196709 384915 196775 384918
rect 357893 384706 357959 384709
rect 356132 384704 357959 384706
rect 356132 384648 357898 384704
rect 357954 384648 357959 384704
rect 356132 384646 357959 384648
rect 357893 384643 357959 384646
rect -960 384284 480 384524
rect 91093 384298 91159 384301
rect 120206 384298 120212 384300
rect 91093 384296 120212 384298
rect 91093 384240 91098 384296
rect 91154 384240 120212 384296
rect 91093 384238 120212 384240
rect 91093 384235 91159 384238
rect 120206 384236 120212 384238
rect 120276 384236 120282 384300
rect 103421 383074 103487 383077
rect 155217 383074 155283 383077
rect 103421 383072 155283 383074
rect 103421 383016 103426 383072
rect 103482 383016 155222 383072
rect 155278 383016 155283 383072
rect 103421 383014 155283 383016
rect 103421 383011 103487 383014
rect 155217 383011 155283 383014
rect 43989 382938 44055 382941
rect 122598 382938 122604 382940
rect 43989 382936 122604 382938
rect 43989 382880 43994 382936
rect 44050 382880 122604 382936
rect 43989 382878 122604 382880
rect 43989 382875 44055 382878
rect 122598 382876 122604 382878
rect 122668 382876 122674 382940
rect 356094 382604 356100 382668
rect 356164 382666 356170 382668
rect 356462 382666 356468 382668
rect 356164 382606 356468 382666
rect 356164 382604 356170 382606
rect 356462 382604 356468 382606
rect 356532 382604 356538 382668
rect 198825 382530 198891 382533
rect 198825 382528 200100 382530
rect 198825 382472 198830 382528
rect 198886 382472 200100 382528
rect 198825 382470 200100 382472
rect 198825 382467 198891 382470
rect 173801 382394 173867 382397
rect 193121 382394 193187 382397
rect 173801 382392 193187 382394
rect 173801 382336 173806 382392
rect 173862 382336 193126 382392
rect 193182 382336 193187 382392
rect 173801 382334 193187 382336
rect 173801 382331 173867 382334
rect 193121 382331 193187 382334
rect 356102 381988 356162 382228
rect 356094 381924 356100 381988
rect 356164 381924 356170 381988
rect 80053 381578 80119 381581
rect 194542 381578 194548 381580
rect 80053 381576 194548 381578
rect 80053 381520 80058 381576
rect 80114 381520 194548 381576
rect 80053 381518 194548 381520
rect 80053 381515 80119 381518
rect 194542 381516 194548 381518
rect 194612 381516 194618 381580
rect 69657 380218 69723 380221
rect 195237 380218 195303 380221
rect 69657 380216 195303 380218
rect 69657 380160 69662 380216
rect 69718 380160 195242 380216
rect 195298 380160 195303 380216
rect 69657 380158 195303 380160
rect 69657 380155 69723 380158
rect 195237 380155 195303 380158
rect 197353 380218 197419 380221
rect 197353 380216 200100 380218
rect 197353 380160 197358 380216
rect 197414 380160 200100 380216
rect 197353 380158 200100 380160
rect 197353 380155 197419 380158
rect 357893 379810 357959 379813
rect 356132 379808 357959 379810
rect 356132 379752 357898 379808
rect 357954 379752 357959 379808
rect 356132 379750 357959 379752
rect 357893 379747 357959 379750
rect 55029 379402 55095 379405
rect 178033 379402 178099 379405
rect 178401 379402 178467 379405
rect 55029 379400 178467 379402
rect 55029 379344 55034 379400
rect 55090 379344 178038 379400
rect 178094 379344 178406 379400
rect 178462 379344 178467 379400
rect 55029 379342 178467 379344
rect 55029 379339 55095 379342
rect 178033 379339 178099 379342
rect 178401 379339 178467 379342
rect 67766 378660 67772 378724
rect 67836 378722 67842 378724
rect 124949 378722 125015 378725
rect 67836 378720 125015 378722
rect 67836 378664 124954 378720
rect 125010 378664 125015 378720
rect 67836 378662 125015 378664
rect 67836 378660 67842 378662
rect 124949 378659 125015 378662
rect 178401 378722 178467 378725
rect 195237 378722 195303 378725
rect 178401 378720 195303 378722
rect 178401 378664 178406 378720
rect 178462 378664 195242 378720
rect 195298 378664 195303 378720
rect 178401 378662 195303 378664
rect 178401 378659 178467 378662
rect 195237 378659 195303 378662
rect 583520 378450 584960 378540
rect 567150 378390 584960 378450
rect 136633 378178 136699 378181
rect 137921 378178 137987 378181
rect 136633 378176 200130 378178
rect 136633 378120 136638 378176
rect 136694 378120 137926 378176
rect 137982 378120 200130 378176
rect 136633 378118 200130 378120
rect 136633 378115 136699 378118
rect 137921 378115 137987 378118
rect 90357 378042 90423 378045
rect 90357 378040 122850 378042
rect 90357 377984 90362 378040
rect 90418 377984 122850 378040
rect 90357 377982 122850 377984
rect 90357 377979 90423 377982
rect 116577 377906 116643 377909
rect 117129 377906 117195 377909
rect 116577 377904 117195 377906
rect 116577 377848 116582 377904
rect 116638 377848 117134 377904
rect 117190 377848 117195 377904
rect 116577 377846 117195 377848
rect 122790 377906 122850 377982
rect 132493 377906 132559 377909
rect 122790 377904 132559 377906
rect 122790 377848 132498 377904
rect 132554 377848 132559 377904
rect 122790 377846 132559 377848
rect 116577 377843 116643 377846
rect 117129 377843 117195 377846
rect 132493 377843 132559 377846
rect 200070 377634 200130 378118
rect 359406 378116 359412 378180
rect 359476 378178 359482 378180
rect 567150 378178 567210 378390
rect 583520 378300 584960 378390
rect 359476 378118 567210 378178
rect 359476 378116 359482 378118
rect 201309 377634 201375 377637
rect 200070 377632 201375 377634
rect 200070 377576 201314 377632
rect 201370 377576 201375 377632
rect 200070 377574 201375 377576
rect 201309 377571 201375 377574
rect 194501 377498 194567 377501
rect 201585 377498 201651 377501
rect 194501 377496 201651 377498
rect 194501 377440 194506 377496
rect 194562 377440 201590 377496
rect 201646 377440 201651 377496
rect 194501 377438 201651 377440
rect 194501 377435 194567 377438
rect 201585 377435 201651 377438
rect 352557 377498 352623 377501
rect 356145 377498 356211 377501
rect 352557 377496 356211 377498
rect 352557 377440 352562 377496
rect 352618 377440 356150 377496
rect 356206 377440 356211 377496
rect 352557 377438 356211 377440
rect 352557 377435 352623 377438
rect 356145 377435 356211 377438
rect 179270 377300 179276 377364
rect 179340 377362 179346 377364
rect 187141 377362 187207 377365
rect 583201 377362 583267 377365
rect 179340 377360 187207 377362
rect 179340 377304 187146 377360
rect 187202 377304 187207 377360
rect 179340 377302 187207 377304
rect 179340 377300 179346 377302
rect 187141 377299 187207 377302
rect 412590 377360 583267 377362
rect 412590 377304 583206 377360
rect 583262 377304 583267 377360
rect 412590 377302 583267 377304
rect 116577 376954 116643 376957
rect 272701 376954 272767 376957
rect 116577 376952 272767 376954
rect 116577 376896 116582 376952
rect 116638 376896 272706 376952
rect 272762 376896 272767 376952
rect 116577 376894 272767 376896
rect 116577 376891 116643 376894
rect 272701 376891 272767 376894
rect 344001 376954 344067 376957
rect 359406 376954 359412 376956
rect 344001 376952 359412 376954
rect 344001 376896 344006 376952
rect 344062 376896 359412 376952
rect 344001 376894 359412 376896
rect 344001 376891 344067 376894
rect 359406 376892 359412 376894
rect 359476 376892 359482 376956
rect 412590 376821 412650 377302
rect 583201 377299 583267 377302
rect 129089 376818 129155 376821
rect 129641 376818 129707 376821
rect 176101 376818 176167 376821
rect 129089 376816 176167 376818
rect 129089 376760 129094 376816
rect 129150 376760 129646 376816
rect 129702 376760 176106 376816
rect 176162 376760 176167 376816
rect 129089 376758 176167 376760
rect 129089 376755 129155 376758
rect 129641 376755 129707 376758
rect 176101 376755 176167 376758
rect 192661 376818 192727 376821
rect 218237 376818 218303 376821
rect 281349 376818 281415 376821
rect 412541 376818 412650 376821
rect 192661 376816 218303 376818
rect 192661 376760 192666 376816
rect 192722 376760 218242 376816
rect 218298 376760 218303 376816
rect 192661 376758 218303 376760
rect 192661 376755 192727 376758
rect 218237 376755 218303 376758
rect 281214 376816 412650 376818
rect 281214 376760 281354 376816
rect 281410 376760 412546 376816
rect 412602 376760 412650 376816
rect 281214 376758 412650 376760
rect 65885 376682 65951 376685
rect 280153 376682 280219 376685
rect 281214 376682 281274 376758
rect 281349 376755 281415 376758
rect 412541 376755 412607 376758
rect 65885 376680 281274 376682
rect 65885 376624 65890 376680
rect 65946 376624 280158 376680
rect 280214 376624 281274 376680
rect 65885 376622 281274 376624
rect 319621 376682 319687 376685
rect 582833 376682 582899 376685
rect 319621 376680 582899 376682
rect 319621 376624 319626 376680
rect 319682 376624 582838 376680
rect 582894 376624 582899 376680
rect 319621 376622 582899 376624
rect 65885 376619 65951 376622
rect 280153 376619 280219 376622
rect 319621 376619 319687 376622
rect 582833 376619 582899 376622
rect 199878 376484 199884 376548
rect 199948 376546 199954 376548
rect 200021 376546 200087 376549
rect 199948 376544 200087 376546
rect 199948 376488 200026 376544
rect 200082 376488 200087 376544
rect 199948 376486 200087 376488
rect 199948 376484 199954 376486
rect 200021 376483 200087 376486
rect 348417 376546 348483 376549
rect 352230 376546 352236 376548
rect 348417 376544 352236 376546
rect 348417 376488 348422 376544
rect 348478 376488 352236 376544
rect 348417 376486 352236 376488
rect 348417 376483 348483 376486
rect 352230 376484 352236 376486
rect 352300 376484 352306 376548
rect 195881 376138 195947 376141
rect 205725 376138 205791 376141
rect 195881 376136 205791 376138
rect 195881 376080 195886 376136
rect 195942 376080 205730 376136
rect 205786 376080 205791 376136
rect 195881 376078 205791 376080
rect 195881 376075 195947 376078
rect 205725 376075 205791 376078
rect 185577 376002 185643 376005
rect 202229 376002 202295 376005
rect 185577 376000 202295 376002
rect 185577 375944 185582 376000
rect 185638 375944 202234 376000
rect 202290 375944 202295 376000
rect 185577 375942 202295 375944
rect 185577 375939 185643 375942
rect 202229 375939 202295 375942
rect 353937 376002 354003 376005
rect 361849 376002 361915 376005
rect 353937 376000 361915 376002
rect 353937 375944 353942 376000
rect 353998 375944 361854 376000
rect 361910 375944 361915 376000
rect 353937 375942 361915 375944
rect 353937 375939 354003 375942
rect 361849 375939 361915 375942
rect 354673 375732 354739 375733
rect 354622 375668 354628 375732
rect 354692 375730 354739 375732
rect 354692 375728 354784 375730
rect 354734 375672 354784 375728
rect 354692 375670 354784 375672
rect 354692 375668 354739 375670
rect 354673 375667 354739 375668
rect 71681 375458 71747 375461
rect 178861 375458 178927 375461
rect 71681 375456 178927 375458
rect 71681 375400 71686 375456
rect 71742 375400 178866 375456
rect 178922 375400 178927 375456
rect 71681 375398 178927 375400
rect 71681 375395 71747 375398
rect 178861 375395 178927 375398
rect 194542 375260 194548 375324
rect 194612 375322 194618 375324
rect 241421 375322 241487 375325
rect 194612 375320 241487 375322
rect 194612 375264 241426 375320
rect 241482 375264 241487 375320
rect 194612 375262 241487 375264
rect 194612 375260 194618 375262
rect 241421 375259 241487 375262
rect 288750 375260 288756 375324
rect 288820 375322 288826 375324
rect 289629 375322 289695 375325
rect 288820 375320 289695 375322
rect 288820 375264 289634 375320
rect 289690 375264 289695 375320
rect 288820 375262 289695 375264
rect 288820 375260 288826 375262
rect 289629 375259 289695 375262
rect 339493 375322 339559 375325
rect 342897 375322 342963 375325
rect 339493 375320 342963 375322
rect 339493 375264 339498 375320
rect 339554 375264 342902 375320
rect 342958 375264 342963 375320
rect 339493 375262 342963 375264
rect 339493 375259 339559 375262
rect 342897 375259 342963 375262
rect 215201 375186 215267 375189
rect 218237 375186 218303 375189
rect 215201 375184 218303 375186
rect 215201 375128 215206 375184
rect 215262 375128 218242 375184
rect 218298 375128 218303 375184
rect 215201 375126 218303 375128
rect 215201 375123 215267 375126
rect 218237 375123 218303 375126
rect 342897 374778 342963 374781
rect 381537 374778 381603 374781
rect 342897 374776 381603 374778
rect 342897 374720 342902 374776
rect 342958 374720 381542 374776
rect 381598 374720 381603 374776
rect 342897 374718 381603 374720
rect 342897 374715 342963 374718
rect 381537 374715 381603 374718
rect 274081 374642 274147 374645
rect 287973 374642 288039 374645
rect 274081 374640 288039 374642
rect 274081 374584 274086 374640
rect 274142 374584 287978 374640
rect 288034 374584 288039 374640
rect 274081 374582 288039 374584
rect 274081 374579 274147 374582
rect 287973 374579 288039 374582
rect 351085 374642 351151 374645
rect 407849 374642 407915 374645
rect 351085 374640 407915 374642
rect 351085 374584 351090 374640
rect 351146 374584 407854 374640
rect 407910 374584 407915 374640
rect 351085 374582 407915 374584
rect 351085 374579 351151 374582
rect 407849 374579 407915 374582
rect 60641 374098 60707 374101
rect 214557 374098 214623 374101
rect 60641 374096 214623 374098
rect 60641 374040 60646 374096
rect 60702 374040 214562 374096
rect 214618 374040 214623 374096
rect 60641 374038 214623 374040
rect 60641 374035 60707 374038
rect 214557 374035 214623 374038
rect 241421 374098 241487 374101
rect 248045 374098 248111 374101
rect 241421 374096 248111 374098
rect 241421 374040 241426 374096
rect 241482 374040 248050 374096
rect 248106 374040 248111 374096
rect 241421 374038 248111 374040
rect 241421 374035 241487 374038
rect 248045 374035 248111 374038
rect 264237 374098 264303 374101
rect 273897 374098 273963 374101
rect 264237 374096 273963 374098
rect 264237 374040 264242 374096
rect 264298 374040 273902 374096
rect 273958 374040 273963 374096
rect 264237 374038 273963 374040
rect 264237 374035 264303 374038
rect 273897 374035 273963 374038
rect 354029 374098 354095 374101
rect 356462 374098 356468 374100
rect 354029 374096 356468 374098
rect 354029 374040 354034 374096
rect 354090 374040 356468 374096
rect 354029 374038 356468 374040
rect 354029 374035 354095 374038
rect 356462 374036 356468 374038
rect 356532 374036 356538 374100
rect 114553 373418 114619 373421
rect 356421 373418 356487 373421
rect 374637 373418 374703 373421
rect 114553 373416 374703 373418
rect 114553 373360 114558 373416
rect 114614 373360 356426 373416
rect 356482 373360 374642 373416
rect 374698 373360 374703 373416
rect 114553 373358 374703 373360
rect 114553 373355 114619 373358
rect 356421 373355 356487 373358
rect 374637 373355 374703 373358
rect 56317 373282 56383 373285
rect 357566 373282 357572 373284
rect 56317 373280 357572 373282
rect 56317 373224 56322 373280
rect 56378 373224 357572 373280
rect 56317 373222 357572 373224
rect 56317 373219 56383 373222
rect 357566 373220 357572 373222
rect 357636 373220 357642 373284
rect 180558 371860 180564 371924
rect 180628 371922 180634 371924
rect 357433 371922 357499 371925
rect 180628 371920 357499 371922
rect 180628 371864 357438 371920
rect 357494 371864 357499 371920
rect 180628 371862 357499 371864
rect 180628 371860 180634 371862
rect 357433 371859 357499 371862
rect -960 371378 480 371468
rect 2957 371378 3023 371381
rect -960 371376 3023 371378
rect -960 371320 2962 371376
rect 3018 371320 3023 371376
rect -960 371318 3023 371320
rect -960 371228 480 371318
rect 2957 371315 3023 371318
rect 59261 371378 59327 371381
rect 220813 371378 220879 371381
rect 221457 371378 221523 371381
rect 59261 371376 221523 371378
rect 59261 371320 59266 371376
rect 59322 371320 220818 371376
rect 220874 371320 221462 371376
rect 221518 371320 221523 371376
rect 59261 371318 221523 371320
rect 59261 371315 59327 371318
rect 220813 371315 220879 371318
rect 221457 371315 221523 371318
rect 358077 371378 358143 371381
rect 358854 371378 358860 371380
rect 358077 371376 358860 371378
rect 358077 371320 358082 371376
rect 358138 371320 358860 371376
rect 358077 371318 358860 371320
rect 358077 371315 358143 371318
rect 358854 371316 358860 371318
rect 358924 371316 358930 371380
rect 198774 370772 198780 370836
rect 198844 370834 198850 370836
rect 218697 370834 218763 370837
rect 198844 370832 218763 370834
rect 198844 370776 218702 370832
rect 218758 370776 218763 370832
rect 198844 370774 218763 370776
rect 198844 370772 198850 370774
rect 218697 370771 218763 370774
rect 82670 370636 82676 370700
rect 82740 370698 82746 370700
rect 133137 370698 133203 370701
rect 82740 370696 133203 370698
rect 82740 370640 133142 370696
rect 133198 370640 133203 370696
rect 82740 370638 133203 370640
rect 82740 370636 82746 370638
rect 133137 370635 133203 370638
rect 213678 370636 213684 370700
rect 213748 370698 213754 370700
rect 245653 370698 245719 370701
rect 213748 370696 245719 370698
rect 213748 370640 245658 370696
rect 245714 370640 245719 370696
rect 213748 370638 245719 370640
rect 213748 370636 213754 370638
rect 245653 370635 245719 370638
rect 67766 370500 67772 370564
rect 67836 370562 67842 370564
rect 123477 370562 123543 370565
rect 67836 370560 123543 370562
rect 67836 370504 123482 370560
rect 123538 370504 123543 370560
rect 67836 370502 123543 370504
rect 67836 370500 67842 370502
rect 123477 370499 123543 370502
rect 128997 370562 129063 370565
rect 168557 370562 168623 370565
rect 128997 370560 168623 370562
rect 128997 370504 129002 370560
rect 129058 370504 168562 370560
rect 168618 370504 168623 370560
rect 128997 370502 168623 370504
rect 128997 370499 129063 370502
rect 168557 370499 168623 370502
rect 184381 370562 184447 370565
rect 250294 370562 250300 370564
rect 184381 370560 250300 370562
rect 184381 370504 184386 370560
rect 184442 370504 250300 370560
rect 184381 370502 250300 370504
rect 184381 370499 184447 370502
rect 250294 370500 250300 370502
rect 250364 370500 250370 370564
rect 356789 370562 356855 370565
rect 364425 370562 364491 370565
rect 356789 370560 364491 370562
rect 356789 370504 356794 370560
rect 356850 370504 364430 370560
rect 364486 370504 364491 370560
rect 356789 370502 364491 370504
rect 356789 370499 356855 370502
rect 364425 370499 364491 370502
rect 111057 369882 111123 369885
rect 111558 369882 111564 369884
rect 111057 369880 111564 369882
rect 111057 369824 111062 369880
rect 111118 369824 111564 369880
rect 111057 369822 111564 369824
rect 111057 369819 111123 369822
rect 111558 369820 111564 369822
rect 111628 369882 111634 369884
rect 183093 369882 183159 369885
rect 111628 369880 183159 369882
rect 111628 369824 183098 369880
rect 183154 369824 183159 369880
rect 111628 369822 183159 369824
rect 111628 369820 111634 369822
rect 183093 369819 183159 369822
rect 132401 369202 132467 369205
rect 209129 369202 209195 369205
rect 132401 369200 209195 369202
rect 132401 369144 132406 369200
rect 132462 369144 209134 369200
rect 209190 369144 209195 369200
rect 132401 369142 209195 369144
rect 132401 369139 132467 369142
rect 209129 369139 209195 369142
rect 129733 369066 129799 369069
rect 163497 369066 163563 369069
rect 376753 369066 376819 369069
rect 129733 369064 376819 369066
rect 129733 369008 129738 369064
rect 129794 369008 163502 369064
rect 163558 369008 376758 369064
rect 376814 369008 376819 369064
rect 129733 369006 376819 369008
rect 129733 369003 129799 369006
rect 163497 369003 163563 369006
rect 376753 369003 376819 369006
rect 71037 368522 71103 368525
rect 121678 368522 121684 368524
rect 71037 368520 121684 368522
rect 71037 368464 71042 368520
rect 71098 368464 121684 368520
rect 71037 368462 121684 368464
rect 71037 368459 71103 368462
rect 121678 368460 121684 368462
rect 121748 368460 121754 368524
rect 85573 368386 85639 368389
rect 86217 368386 86283 368389
rect 85573 368384 86283 368386
rect 85573 368328 85578 368384
rect 85634 368328 86222 368384
rect 86278 368328 86283 368384
rect 85573 368326 86283 368328
rect 85573 368323 85639 368326
rect 86217 368323 86283 368326
rect 195881 368386 195947 368389
rect 360326 368386 360332 368388
rect 195881 368384 360332 368386
rect 195881 368328 195886 368384
rect 195942 368328 360332 368384
rect 195881 368326 360332 368328
rect 195881 368323 195947 368326
rect 360326 368324 360332 368326
rect 360396 368324 360402 368388
rect 191097 367842 191163 367845
rect 200205 367842 200271 367845
rect 191097 367840 200271 367842
rect 191097 367784 191102 367840
rect 191158 367784 200210 367840
rect 200266 367784 200271 367840
rect 191097 367782 200271 367784
rect 191097 367779 191163 367782
rect 200205 367779 200271 367782
rect 200798 367780 200804 367844
rect 200868 367842 200874 367844
rect 260833 367842 260899 367845
rect 200868 367840 260899 367842
rect 200868 367784 260838 367840
rect 260894 367784 260899 367840
rect 200868 367782 260899 367784
rect 200868 367780 200874 367782
rect 260833 367779 260899 367782
rect 114461 367706 114527 367709
rect 354673 367706 354739 367709
rect 114461 367704 354739 367706
rect 114461 367648 114466 367704
rect 114522 367648 354678 367704
rect 354734 367648 354739 367704
rect 114461 367646 354739 367648
rect 114461 367643 114527 367646
rect 354673 367643 354739 367646
rect 86217 367162 86283 367165
rect 188429 367162 188495 367165
rect 86217 367160 188495 367162
rect 86217 367104 86222 367160
rect 86278 367104 188434 367160
rect 188490 367104 188495 367160
rect 86217 367102 188495 367104
rect 86217 367099 86283 367102
rect 188429 367099 188495 367102
rect 178769 366482 178835 366485
rect 205817 366482 205883 366485
rect 178769 366480 205883 366482
rect 178769 366424 178774 366480
rect 178830 366424 205822 366480
rect 205878 366424 205883 366480
rect 178769 366422 205883 366424
rect 178769 366419 178835 366422
rect 205817 366419 205883 366422
rect 75821 366346 75887 366349
rect 195094 366346 195100 366348
rect 75821 366344 195100 366346
rect 75821 366288 75826 366344
rect 75882 366288 195100 366344
rect 75821 366286 195100 366288
rect 75821 366283 75887 366286
rect 195094 366284 195100 366286
rect 195164 366284 195170 366348
rect 208393 366346 208459 366349
rect 307017 366346 307083 366349
rect 208393 366344 307083 366346
rect 208393 366288 208398 366344
rect 208454 366288 307022 366344
rect 307078 366288 307083 366344
rect 208393 366286 307083 366288
rect 208393 366283 208459 366286
rect 307017 366283 307083 366286
rect 85481 365802 85547 365805
rect 230473 365802 230539 365805
rect 231117 365802 231183 365805
rect 85481 365800 231183 365802
rect 85481 365744 85486 365800
rect 85542 365744 230478 365800
rect 230534 365744 231122 365800
rect 231178 365744 231183 365800
rect 85481 365742 231183 365744
rect 85481 365739 85547 365742
rect 230473 365739 230539 365742
rect 231117 365739 231183 365742
rect 118601 365668 118667 365669
rect 118550 365604 118556 365668
rect 118620 365666 118667 365668
rect 118620 365664 118712 365666
rect 118662 365608 118712 365664
rect 118620 365606 118712 365608
rect 118620 365604 118667 365606
rect 118601 365603 118667 365604
rect 582373 365122 582439 365125
rect 583520 365122 584960 365212
rect 582373 365120 584960 365122
rect 582373 365064 582378 365120
rect 582434 365064 584960 365120
rect 582373 365062 584960 365064
rect 582373 365059 582439 365062
rect 81014 364924 81020 364988
rect 81084 364986 81090 364988
rect 356278 364986 356284 364988
rect 81084 364926 356284 364986
rect 81084 364924 81090 364926
rect 356278 364924 356284 364926
rect 356348 364924 356354 364988
rect 583520 364972 584960 365062
rect 118601 364442 118667 364445
rect 238017 364442 238083 364445
rect 118601 364440 238083 364442
rect 118601 364384 118606 364440
rect 118662 364384 238022 364440
rect 238078 364384 238083 364440
rect 118601 364382 238083 364384
rect 118601 364379 118667 364382
rect 238017 364379 238083 364382
rect 114318 364244 114324 364308
rect 114388 364306 114394 364308
rect 118509 364306 118575 364309
rect 114388 364304 118575 364306
rect 114388 364248 118514 364304
rect 118570 364248 118575 364304
rect 114388 364246 118575 364248
rect 114388 364244 114394 364246
rect 118509 364243 118575 364246
rect 196709 364306 196775 364309
rect 583017 364306 583083 364309
rect 196709 364304 583083 364306
rect 196709 364248 196714 364304
rect 196770 364248 583022 364304
rect 583078 364248 583083 364304
rect 196709 364246 583083 364248
rect 196709 364243 196775 364246
rect 583017 364243 583083 364246
rect 63309 363762 63375 363765
rect 111742 363762 111748 363764
rect 63309 363760 111748 363762
rect 63309 363704 63314 363760
rect 63370 363704 111748 363760
rect 63309 363702 111748 363704
rect 63309 363699 63375 363702
rect 111742 363700 111748 363702
rect 111812 363700 111818 363764
rect 190310 363700 190316 363764
rect 190380 363762 190386 363764
rect 202873 363762 202939 363765
rect 190380 363760 202939 363762
rect 190380 363704 202878 363760
rect 202934 363704 202939 363760
rect 190380 363702 202939 363704
rect 190380 363700 190386 363702
rect 202873 363699 202939 363702
rect 108941 363626 109007 363629
rect 161473 363626 161539 363629
rect 108941 363624 161539 363626
rect 108941 363568 108946 363624
rect 109002 363568 161478 363624
rect 161534 363568 161539 363624
rect 108941 363566 161539 363568
rect 108941 363563 109007 363566
rect 161473 363563 161539 363566
rect 177389 363626 177455 363629
rect 308397 363626 308463 363629
rect 177389 363624 308463 363626
rect 177389 363568 177394 363624
rect 177450 363568 308402 363624
rect 308458 363568 308463 363624
rect 177389 363566 308463 363568
rect 177389 363563 177455 363566
rect 308397 363563 308463 363566
rect 144729 363218 144795 363221
rect 190310 363218 190316 363220
rect 144729 363216 190316 363218
rect 144729 363160 144734 363216
rect 144790 363160 190316 363216
rect 144729 363158 190316 363160
rect 144729 363155 144795 363158
rect 190310 363156 190316 363158
rect 190380 363156 190386 363220
rect 100661 363082 100727 363085
rect 187141 363082 187207 363085
rect 100661 363080 187207 363082
rect 100661 363024 100666 363080
rect 100722 363024 187146 363080
rect 187202 363024 187207 363080
rect 100661 363022 187207 363024
rect 100661 363019 100727 363022
rect 187141 363019 187207 363022
rect 229093 362538 229159 362541
rect 240358 362538 240364 362540
rect 229093 362536 240364 362538
rect 229093 362480 229098 362536
rect 229154 362480 240364 362536
rect 229093 362478 240364 362480
rect 229093 362475 229159 362478
rect 240358 362476 240364 362478
rect 240428 362476 240434 362540
rect 72734 362340 72740 362404
rect 72804 362402 72810 362404
rect 123477 362402 123543 362405
rect 72804 362400 123543 362402
rect 72804 362344 123482 362400
rect 123538 362344 123543 362400
rect 72804 362342 123543 362344
rect 72804 362340 72810 362342
rect 123477 362339 123543 362342
rect 151077 362402 151143 362405
rect 154614 362402 154620 362404
rect 151077 362400 154620 362402
rect 151077 362344 151082 362400
rect 151138 362344 154620 362400
rect 151077 362342 154620 362344
rect 151077 362339 151143 362342
rect 154614 362340 154620 362342
rect 154684 362340 154690 362404
rect 233141 362402 233207 362405
rect 371325 362402 371391 362405
rect 233141 362400 371391 362402
rect 233141 362344 233146 362400
rect 233202 362344 371330 362400
rect 371386 362344 371391 362400
rect 233141 362342 371391 362344
rect 233141 362339 233207 362342
rect 371325 362339 371391 362342
rect 121678 362204 121684 362268
rect 121748 362266 121754 362268
rect 195237 362266 195303 362269
rect 121748 362264 195303 362266
rect 121748 362208 195242 362264
rect 195298 362208 195303 362264
rect 121748 362206 195303 362208
rect 121748 362204 121754 362206
rect 195237 362203 195303 362206
rect 201401 362266 201467 362269
rect 341517 362266 341583 362269
rect 201401 362264 341583 362266
rect 201401 362208 201406 362264
rect 201462 362208 341522 362264
rect 341578 362208 341583 362264
rect 201401 362206 341583 362208
rect 201401 362203 201467 362206
rect 341517 362203 341583 362206
rect 94497 361722 94563 361725
rect 95049 361722 95115 361725
rect 232497 361722 232563 361725
rect 233141 361722 233207 361725
rect 94497 361720 233207 361722
rect 94497 361664 94502 361720
rect 94558 361664 95054 361720
rect 95110 361664 232502 361720
rect 232558 361664 233146 361720
rect 233202 361664 233207 361720
rect 94497 361662 233207 361664
rect 94497 361659 94563 361662
rect 95049 361659 95115 361662
rect 232497 361659 232563 361662
rect 233141 361659 233207 361662
rect 67950 360844 67956 360908
rect 68020 360906 68026 360908
rect 86217 360906 86283 360909
rect 68020 360904 86283 360906
rect 68020 360848 86222 360904
rect 86278 360848 86283 360904
rect 68020 360846 86283 360848
rect 68020 360844 68026 360846
rect 86217 360843 86283 360846
rect 133781 360498 133847 360501
rect 174537 360498 174603 360501
rect 174721 360498 174787 360501
rect 133781 360496 174787 360498
rect 133781 360440 133786 360496
rect 133842 360440 174542 360496
rect 174598 360440 174726 360496
rect 174782 360440 174787 360496
rect 133781 360438 174787 360440
rect 133781 360435 133847 360438
rect 174537 360435 174603 360438
rect 174721 360435 174787 360438
rect 101949 360362 102015 360365
rect 188337 360362 188403 360365
rect 101949 360360 188403 360362
rect 101949 360304 101954 360360
rect 102010 360304 188342 360360
rect 188398 360304 188403 360360
rect 101949 360302 188403 360304
rect 101949 360299 102015 360302
rect 188337 360299 188403 360302
rect 85389 360226 85455 360229
rect 89662 360226 89668 360228
rect 85389 360224 89668 360226
rect 85389 360168 85394 360224
rect 85450 360168 89668 360224
rect 85389 360166 89668 360168
rect 85389 360163 85455 360166
rect 89662 360164 89668 360166
rect 89732 360164 89738 360228
rect 113173 360226 113239 360229
rect 114461 360226 114527 360229
rect 246297 360226 246363 360229
rect 113173 360224 246363 360226
rect 113173 360168 113178 360224
rect 113234 360168 114466 360224
rect 114522 360168 246302 360224
rect 246358 360168 246363 360224
rect 113173 360166 246363 360168
rect 113173 360163 113239 360166
rect 114461 360163 114527 360166
rect 246297 360163 246363 360166
rect 150341 359546 150407 359549
rect 178677 359546 178743 359549
rect 150341 359544 178743 359546
rect 150341 359488 150346 359544
rect 150402 359488 178682 359544
rect 178738 359488 178743 359544
rect 150341 359486 178743 359488
rect 150341 359483 150407 359486
rect 178677 359483 178743 359486
rect 206870 359484 206876 359548
rect 206940 359546 206946 359548
rect 213269 359546 213335 359549
rect 283557 359546 283623 359549
rect 285581 359546 285647 359549
rect 206940 359544 213335 359546
rect 206940 359488 213274 359544
rect 213330 359488 213335 359544
rect 206940 359486 213335 359488
rect 206940 359484 206946 359486
rect 213269 359483 213335 359486
rect 277350 359544 285647 359546
rect 277350 359488 283562 359544
rect 283618 359488 285586 359544
rect 285642 359488 285647 359544
rect 277350 359486 285647 359488
rect 66110 359348 66116 359412
rect 66180 359410 66186 359412
rect 277350 359410 277410 359486
rect 283557 359483 283623 359486
rect 285581 359483 285647 359486
rect 66180 359350 277410 359410
rect 66180 359348 66186 359350
rect 70577 358866 70643 358869
rect 71589 358866 71655 358869
rect 195513 358866 195579 358869
rect 70577 358864 195579 358866
rect 70577 358808 70582 358864
rect 70638 358808 71594 358864
rect 71650 358808 195518 358864
rect 195574 358808 195579 358864
rect 70577 358806 195579 358808
rect 70577 358803 70643 358806
rect 71589 358803 71655 358806
rect 195513 358803 195579 358806
rect -960 358458 480 358548
rect 3417 358458 3483 358461
rect -960 358456 3483 358458
rect -960 358400 3422 358456
rect 3478 358400 3483 358456
rect -960 358398 3483 358400
rect -960 358308 480 358398
rect 3417 358395 3483 358398
rect 337377 358050 337443 358053
rect 357525 358050 357591 358053
rect 335310 358048 357591 358050
rect 335310 357992 337382 358048
rect 337438 357992 357530 358048
rect 357586 357992 357591 358048
rect 335310 357990 357591 357992
rect 82905 357642 82971 357645
rect 84101 357642 84167 357645
rect 244917 357642 244983 357645
rect 82905 357640 244983 357642
rect 82905 357584 82910 357640
rect 82966 357584 84106 357640
rect 84162 357584 244922 357640
rect 244978 357584 244983 357640
rect 82905 357582 244983 357584
rect 82905 357579 82971 357582
rect 84101 357579 84167 357582
rect 244917 357579 244983 357582
rect 69790 357444 69796 357508
rect 69860 357506 69866 357508
rect 335310 357506 335370 357990
rect 337377 357987 337443 357990
rect 357525 357987 357591 357990
rect 69860 357446 335370 357506
rect 69860 357444 69866 357446
rect 155217 356826 155283 356829
rect 172513 356826 172579 356829
rect 155217 356824 172579 356826
rect 155217 356768 155222 356824
rect 155278 356768 172518 356824
rect 172574 356768 172579 356824
rect 155217 356766 172579 356768
rect 155217 356763 155283 356766
rect 172513 356763 172579 356766
rect 99189 356690 99255 356693
rect 242157 356690 242223 356693
rect 245009 356690 245075 356693
rect 99189 356688 245075 356690
rect 99189 356632 99194 356688
rect 99250 356632 242162 356688
rect 242218 356632 245014 356688
rect 245070 356632 245075 356688
rect 99189 356630 245075 356632
rect 99189 356627 99255 356630
rect 242157 356627 242223 356630
rect 245009 356627 245075 356630
rect 254577 356690 254643 356693
rect 351177 356690 351243 356693
rect 254577 356688 351243 356690
rect 254577 356632 254582 356688
rect 254638 356632 351182 356688
rect 351238 356632 351243 356688
rect 254577 356630 351243 356632
rect 254577 356627 254643 356630
rect 351177 356627 351243 356630
rect 92473 356146 92539 356149
rect 93669 356146 93735 356149
rect 151077 356146 151143 356149
rect 92473 356144 151143 356146
rect 92473 356088 92478 356144
rect 92534 356088 93674 356144
rect 93730 356088 151082 356144
rect 151138 356088 151143 356144
rect 92473 356086 151143 356088
rect 92473 356083 92539 356086
rect 93669 356083 93735 356086
rect 151077 356083 151143 356086
rect 139301 355466 139367 355469
rect 170581 355466 170647 355469
rect 139301 355464 170647 355466
rect 139301 355408 139306 355464
rect 139362 355408 170586 355464
rect 170642 355408 170647 355464
rect 139301 355406 170647 355408
rect 139301 355403 139367 355406
rect 170581 355403 170647 355406
rect 160737 355330 160803 355333
rect 253289 355330 253355 355333
rect 160737 355328 253355 355330
rect 160737 355272 160742 355328
rect 160798 355272 253294 355328
rect 253350 355272 253355 355328
rect 160737 355270 253355 355272
rect 160737 355267 160803 355270
rect 253289 355267 253355 355270
rect 102133 354786 102199 354789
rect 103421 354786 103487 354789
rect 335997 354786 336063 354789
rect 102133 354784 336063 354786
rect 102133 354728 102138 354784
rect 102194 354728 103426 354784
rect 103482 354728 336002 354784
rect 336058 354728 336063 354784
rect 102133 354726 336063 354728
rect 102133 354723 102199 354726
rect 103421 354723 103487 354726
rect 335997 354723 336063 354726
rect 69054 354588 69060 354652
rect 69124 354650 69130 354652
rect 100661 354650 100727 354653
rect 69124 354648 100727 354650
rect 69124 354592 100666 354648
rect 100722 354592 100727 354648
rect 69124 354590 100727 354592
rect 69124 354588 69130 354590
rect 100661 354587 100727 354590
rect 181621 354650 181687 354653
rect 331857 354650 331923 354653
rect 181621 354648 331923 354650
rect 181621 354592 181626 354648
rect 181682 354592 331862 354648
rect 331918 354592 331923 354648
rect 181621 354590 331923 354592
rect 181621 354587 181687 354590
rect 331857 354587 331923 354590
rect 3509 353970 3575 353973
rect 69054 353970 69060 353972
rect 3509 353968 69060 353970
rect 3509 353912 3514 353968
rect 3570 353912 69060 353968
rect 3509 353910 69060 353912
rect 3509 353907 3575 353910
rect 69054 353908 69060 353910
rect 69124 353908 69130 353972
rect 96521 353970 96587 353973
rect 177849 353970 177915 353973
rect 96521 353968 177915 353970
rect 96521 353912 96526 353968
rect 96582 353912 177854 353968
rect 177910 353912 177915 353968
rect 96521 353910 177915 353912
rect 96521 353907 96587 353910
rect 177849 353907 177915 353910
rect 221457 353970 221523 353973
rect 268326 353970 268332 353972
rect 221457 353968 268332 353970
rect 221457 353912 221462 353968
rect 221518 353912 268332 353968
rect 221457 353910 268332 353912
rect 221457 353907 221523 353910
rect 268326 353908 268332 353910
rect 268396 353908 268402 353972
rect 177849 353562 177915 353565
rect 180006 353562 180012 353564
rect 177849 353560 180012 353562
rect 177849 353504 177854 353560
rect 177910 353504 180012 353560
rect 177849 353502 180012 353504
rect 177849 353499 177915 353502
rect 180006 353500 180012 353502
rect 180076 353500 180082 353564
rect 93117 353426 93183 353429
rect 93710 353426 93716 353428
rect 93117 353424 93716 353426
rect 93117 353368 93122 353424
rect 93178 353368 93716 353424
rect 93117 353366 93716 353368
rect 93117 353363 93183 353366
rect 93710 353364 93716 353366
rect 93780 353426 93786 353428
rect 251909 353426 251975 353429
rect 93780 353424 251975 353426
rect 93780 353368 251914 353424
rect 251970 353368 251975 353424
rect 93780 353366 251975 353368
rect 93780 353364 93786 353366
rect 251909 353363 251975 353366
rect 128169 352066 128235 352069
rect 270401 352066 270467 352069
rect 128169 352064 270467 352066
rect 128169 352008 128174 352064
rect 128230 352008 270406 352064
rect 270462 352008 270467 352064
rect 128169 352006 270467 352008
rect 128169 352003 128235 352006
rect 270401 352003 270467 352006
rect 65977 351930 66043 351933
rect 328453 351930 328519 351933
rect 329097 351930 329163 351933
rect 65977 351928 329163 351930
rect 65977 351872 65982 351928
rect 66038 351872 328458 351928
rect 328514 351872 329102 351928
rect 329158 351872 329163 351928
rect 65977 351870 329163 351872
rect 65977 351867 66043 351870
rect 328453 351867 328519 351870
rect 329097 351867 329163 351870
rect 582833 351930 582899 351933
rect 583520 351930 584960 352020
rect 582833 351928 584960 351930
rect 582833 351872 582838 351928
rect 582894 351872 584960 351928
rect 582833 351870 584960 351872
rect 582833 351867 582899 351870
rect 583520 351780 584960 351870
rect 209630 351324 209636 351388
rect 209700 351386 209706 351388
rect 227713 351386 227779 351389
rect 209700 351384 227779 351386
rect 209700 351328 227718 351384
rect 227774 351328 227779 351384
rect 209700 351326 227779 351328
rect 209700 351324 209706 351326
rect 227713 351323 227779 351326
rect 100661 351250 100727 351253
rect 188889 351250 188955 351253
rect 211889 351250 211955 351253
rect 100661 351248 211955 351250
rect 100661 351192 100666 351248
rect 100722 351192 188894 351248
rect 188950 351192 211894 351248
rect 211950 351192 211955 351248
rect 100661 351190 211955 351192
rect 100661 351187 100727 351190
rect 188889 351187 188955 351190
rect 211889 351187 211955 351190
rect 138013 351114 138079 351117
rect 263685 351114 263751 351117
rect 138013 351112 263751 351114
rect 138013 351056 138018 351112
rect 138074 351056 263690 351112
rect 263746 351056 263751 351112
rect 138013 351054 263751 351056
rect 138013 351051 138079 351054
rect 263685 351051 263751 351054
rect 72918 350508 72924 350572
rect 72988 350570 72994 350572
rect 180057 350570 180123 350573
rect 72988 350568 180123 350570
rect 72988 350512 180062 350568
rect 180118 350512 180123 350568
rect 72988 350510 180123 350512
rect 72988 350508 72994 350510
rect 180057 350507 180123 350510
rect 215293 350434 215359 350437
rect 132450 350432 215359 350434
rect 132450 350376 215298 350432
rect 215354 350376 215359 350432
rect 132450 350374 215359 350376
rect 106181 349890 106247 349893
rect 128353 349890 128419 349893
rect 132450 349890 132510 350374
rect 215293 350371 215359 350374
rect 215293 350026 215359 350029
rect 216029 350026 216095 350029
rect 215293 350024 216095 350026
rect 215293 349968 215298 350024
rect 215354 349968 216034 350024
rect 216090 349968 216095 350024
rect 215293 349966 216095 349968
rect 215293 349963 215359 349966
rect 216029 349963 216095 349966
rect 106181 349888 132510 349890
rect 106181 349832 106186 349888
rect 106242 349832 128358 349888
rect 128414 349832 132510 349888
rect 106181 349830 132510 349832
rect 171869 349890 171935 349893
rect 176653 349890 176719 349893
rect 253197 349890 253263 349893
rect 255957 349890 256023 349893
rect 171869 349888 176719 349890
rect 171869 349832 171874 349888
rect 171930 349832 176658 349888
rect 176714 349832 176719 349888
rect 171869 349830 176719 349832
rect 106181 349827 106247 349830
rect 128353 349827 128419 349830
rect 171869 349827 171935 349830
rect 176653 349827 176719 349830
rect 238710 349888 256023 349890
rect 238710 349832 253202 349888
rect 253258 349832 255962 349888
rect 256018 349832 256023 349888
rect 238710 349830 256023 349832
rect 76557 349754 76623 349757
rect 101857 349754 101923 349757
rect 76557 349752 101923 349754
rect 76557 349696 76562 349752
rect 76618 349696 101862 349752
rect 101918 349696 101923 349752
rect 76557 349694 101923 349696
rect 76557 349691 76623 349694
rect 101857 349691 101923 349694
rect 121729 349754 121795 349757
rect 238710 349754 238770 349830
rect 253197 349827 253263 349830
rect 255957 349827 256023 349830
rect 285581 349890 285647 349893
rect 286174 349890 286180 349892
rect 285581 349888 286180 349890
rect 285581 349832 285586 349888
rect 285642 349832 286180 349888
rect 285581 349830 286180 349832
rect 285581 349827 285647 349830
rect 286174 349828 286180 349830
rect 286244 349828 286250 349892
rect 121729 349752 238770 349754
rect 121729 349696 121734 349752
rect 121790 349696 238770 349752
rect 121729 349694 238770 349696
rect 121729 349691 121795 349694
rect 320265 349074 320331 349077
rect 320817 349074 320883 349077
rect 320265 349072 320883 349074
rect 320265 349016 320270 349072
rect 320326 349016 320822 349072
rect 320878 349016 320883 349072
rect 320265 349014 320883 349016
rect 320265 349011 320331 349014
rect 320817 349011 320883 349014
rect 126237 348122 126303 348125
rect 176009 348122 176075 348125
rect 126237 348120 176075 348122
rect 126237 348064 126242 348120
rect 126298 348064 176014 348120
rect 176070 348064 176075 348120
rect 126237 348062 176075 348064
rect 126237 348059 126303 348062
rect 176009 348059 176075 348062
rect 65926 347924 65932 347988
rect 65996 347986 66002 347988
rect 153837 347986 153903 347989
rect 65996 347984 153903 347986
rect 65996 347928 153842 347984
rect 153898 347928 153903 347984
rect 65996 347926 153903 347928
rect 65996 347924 66002 347926
rect 153837 347923 153903 347926
rect 67357 347850 67423 347853
rect 110413 347850 110479 347853
rect 67357 347848 110479 347850
rect 67357 347792 67362 347848
rect 67418 347792 110418 347848
rect 110474 347792 110479 347848
rect 67357 347790 110479 347792
rect 67357 347787 67423 347790
rect 110413 347787 110479 347790
rect 133689 347850 133755 347853
rect 320817 347850 320883 347853
rect 133689 347848 320883 347850
rect 133689 347792 133694 347848
rect 133750 347792 320822 347848
rect 320878 347792 320883 347848
rect 133689 347790 320883 347792
rect 133689 347787 133755 347790
rect 320817 347787 320883 347790
rect 79317 347170 79383 347173
rect 124857 347170 124923 347173
rect 79317 347168 124923 347170
rect 79317 347112 79322 347168
rect 79378 347112 124862 347168
rect 124918 347112 124923 347168
rect 79317 347110 124923 347112
rect 79317 347107 79383 347110
rect 124857 347107 124923 347110
rect 57697 347034 57763 347037
rect 99966 347034 99972 347036
rect 57697 347032 99972 347034
rect 57697 346976 57702 347032
rect 57758 346976 99972 347032
rect 57697 346974 99972 346976
rect 57697 346971 57763 346974
rect 99966 346972 99972 346974
rect 100036 346972 100042 347036
rect 121453 347034 121519 347037
rect 196709 347034 196775 347037
rect 121453 347032 196775 347034
rect 121453 346976 121458 347032
rect 121514 346976 196714 347032
rect 196770 346976 196775 347032
rect 121453 346974 196775 346976
rect 121453 346971 121519 346974
rect 196709 346971 196775 346974
rect 140773 346626 140839 346629
rect 141417 346626 141483 346629
rect 169569 346626 169635 346629
rect 140773 346624 169635 346626
rect 140773 346568 140778 346624
rect 140834 346568 141422 346624
rect 141478 346568 169574 346624
rect 169630 346568 169635 346624
rect 140773 346566 169635 346568
rect 140773 346563 140839 346566
rect 141417 346563 141483 346566
rect 169569 346563 169635 346566
rect 120717 346490 120783 346493
rect 149053 346490 149119 346493
rect 120717 346488 149119 346490
rect 120717 346432 120722 346488
rect 120778 346432 149058 346488
rect 149114 346432 149119 346488
rect 120717 346430 149119 346432
rect 120717 346427 120783 346430
rect 149053 346427 149119 346430
rect 151721 346490 151787 346493
rect 350441 346490 350507 346493
rect 151721 346488 350507 346490
rect 151721 346432 151726 346488
rect 151782 346432 350446 346488
rect 350502 346432 350507 346488
rect 151721 346430 350507 346432
rect 151721 346427 151787 346430
rect 350441 346427 350507 346430
rect 107745 346354 107811 346357
rect 108297 346354 108363 346357
rect 107745 346352 108363 346354
rect 107745 346296 107750 346352
rect 107806 346296 108302 346352
rect 108358 346296 108363 346352
rect 107745 346294 108363 346296
rect 107745 346291 107811 346294
rect 108297 346291 108363 346294
rect 184289 345946 184355 345949
rect 235349 345946 235415 345949
rect 184289 345944 235415 345946
rect 184289 345888 184294 345944
rect 184350 345888 235354 345944
rect 235410 345888 235415 345944
rect 184289 345886 235415 345888
rect 184289 345883 184355 345886
rect 235349 345883 235415 345886
rect 67265 345810 67331 345813
rect 187233 345810 187299 345813
rect 67265 345808 187299 345810
rect 67265 345752 67270 345808
rect 67326 345752 187238 345808
rect 187294 345752 187299 345808
rect 67265 345750 187299 345752
rect 67265 345747 67331 345750
rect 187233 345747 187299 345750
rect 73153 345674 73219 345677
rect 119470 345674 119476 345676
rect 73153 345672 119476 345674
rect 73153 345616 73158 345672
rect 73214 345616 119476 345672
rect 73153 345614 119476 345616
rect 73153 345611 73219 345614
rect 119470 345612 119476 345614
rect 119540 345612 119546 345676
rect 149053 345674 149119 345677
rect 155217 345674 155283 345677
rect 149053 345672 155283 345674
rect 149053 345616 149058 345672
rect 149114 345616 155222 345672
rect 155278 345616 155283 345672
rect 149053 345614 155283 345616
rect 149053 345611 149119 345614
rect 155217 345611 155283 345614
rect 168281 345674 168347 345677
rect 324313 345674 324379 345677
rect 168281 345672 324379 345674
rect 168281 345616 168286 345672
rect 168342 345616 324318 345672
rect 324374 345616 324379 345672
rect 168281 345614 324379 345616
rect 168281 345611 168347 345614
rect 324313 345611 324379 345614
rect -960 345402 480 345492
rect 3601 345402 3667 345405
rect -960 345400 3667 345402
rect -960 345344 3606 345400
rect 3662 345344 3667 345400
rect -960 345342 3667 345344
rect -960 345252 480 345342
rect 3601 345339 3667 345342
rect 107745 345130 107811 345133
rect 174905 345130 174971 345133
rect 107745 345128 174971 345130
rect 107745 345072 107750 345128
rect 107806 345072 174910 345128
rect 174966 345072 174971 345128
rect 107745 345070 174971 345072
rect 107745 345067 107811 345070
rect 174905 345067 174971 345070
rect 66662 344388 66668 344452
rect 66732 344450 66738 344452
rect 174629 344450 174695 344453
rect 66732 344448 174695 344450
rect 66732 344392 174634 344448
rect 174690 344392 174695 344448
rect 66732 344390 174695 344392
rect 66732 344388 66738 344390
rect 174629 344387 174695 344390
rect 210734 344388 210740 344452
rect 210804 344450 210810 344452
rect 237373 344450 237439 344453
rect 210804 344448 237439 344450
rect 210804 344392 237378 344448
rect 237434 344392 237439 344448
rect 210804 344390 237439 344392
rect 210804 344388 210810 344390
rect 237373 344387 237439 344390
rect 245009 344450 245075 344453
rect 291694 344450 291700 344452
rect 245009 344448 291700 344450
rect 245009 344392 245014 344448
rect 245070 344392 291700 344448
rect 245009 344390 291700 344392
rect 245009 344387 245075 344390
rect 291694 344388 291700 344390
rect 291764 344388 291770 344452
rect 69606 344252 69612 344316
rect 69676 344314 69682 344316
rect 116577 344314 116643 344317
rect 69676 344312 116643 344314
rect 69676 344256 116582 344312
rect 116638 344256 116643 344312
rect 69676 344254 116643 344256
rect 69676 344252 69682 344254
rect 116577 344251 116643 344254
rect 119889 344314 119955 344317
rect 264237 344314 264303 344317
rect 286225 344316 286291 344317
rect 119889 344312 264303 344314
rect 119889 344256 119894 344312
rect 119950 344256 264242 344312
rect 264298 344256 264303 344312
rect 119889 344254 264303 344256
rect 119889 344251 119955 344254
rect 264237 344251 264303 344254
rect 286174 344252 286180 344316
rect 286244 344314 286291 344316
rect 286244 344312 286336 344314
rect 286286 344256 286336 344312
rect 286244 344254 286336 344256
rect 286244 344252 286291 344254
rect 286225 344251 286291 344252
rect 156597 343906 156663 343909
rect 156597 343904 161490 343906
rect 156597 343848 156602 343904
rect 156658 343848 161490 343904
rect 156597 343846 161490 343848
rect 156597 343843 156663 343846
rect 118325 343770 118391 343773
rect 156873 343770 156939 343773
rect 118325 343768 156939 343770
rect 118325 343712 118330 343768
rect 118386 343712 156878 343768
rect 156934 343712 156939 343768
rect 118325 343710 156939 343712
rect 161430 343770 161490 343846
rect 161565 343770 161631 343773
rect 222837 343770 222903 343773
rect 161430 343768 222903 343770
rect 161430 343712 161570 343768
rect 161626 343712 222842 343768
rect 222898 343712 222903 343768
rect 161430 343710 222903 343712
rect 118325 343707 118391 343710
rect 156873 343707 156939 343710
rect 161565 343707 161631 343710
rect 222837 343707 222903 343710
rect 48129 343634 48195 343637
rect 115841 343634 115907 343637
rect 48129 343632 115907 343634
rect 48129 343576 48134 343632
rect 48190 343576 115846 343632
rect 115902 343576 115907 343632
rect 48129 343574 115907 343576
rect 48129 343571 48195 343574
rect 115841 343571 115907 343574
rect 107469 343090 107535 343093
rect 157742 343090 157748 343092
rect 107469 343088 157748 343090
rect 107469 343032 107474 343088
rect 107530 343032 157748 343088
rect 107469 343030 157748 343032
rect 107469 343027 107535 343030
rect 157742 343028 157748 343030
rect 157812 343028 157818 343092
rect 115841 342954 115907 342957
rect 304993 342954 305059 342957
rect 115841 342952 305059 342954
rect 115841 342896 115846 342952
rect 115902 342896 304998 342952
rect 305054 342896 305059 342952
rect 115841 342894 305059 342896
rect 115841 342891 115907 342894
rect 304993 342891 305059 342894
rect 81433 342274 81499 342277
rect 230422 342274 230428 342276
rect 81433 342272 230428 342274
rect 81433 342216 81438 342272
rect 81494 342216 230428 342272
rect 81433 342214 230428 342216
rect 81433 342211 81499 342214
rect 230422 342212 230428 342214
rect 230492 342212 230498 342276
rect 304993 342274 305059 342277
rect 305637 342274 305703 342277
rect 304993 342272 305703 342274
rect 304993 342216 304998 342272
rect 305054 342216 305642 342272
rect 305698 342216 305703 342272
rect 304993 342214 305703 342216
rect 304993 342211 305059 342214
rect 305637 342211 305703 342214
rect 159357 341594 159423 341597
rect 167729 341594 167795 341597
rect 159357 341592 167795 341594
rect 159357 341536 159362 341592
rect 159418 341536 167734 341592
rect 167790 341536 167795 341592
rect 159357 341534 167795 341536
rect 159357 341531 159423 341534
rect 167729 341531 167795 341534
rect 287697 341594 287763 341597
rect 354438 341594 354444 341596
rect 287697 341592 354444 341594
rect 287697 341536 287702 341592
rect 287758 341536 354444 341592
rect 287697 341534 354444 341536
rect 287697 341531 287763 341534
rect 354438 341532 354444 341534
rect 354508 341532 354514 341596
rect 111609 341458 111675 341461
rect 309777 341458 309843 341461
rect 111609 341456 309843 341458
rect 111609 341400 111614 341456
rect 111670 341400 309782 341456
rect 309838 341400 309843 341456
rect 111609 341398 309843 341400
rect 111609 341395 111675 341398
rect 309777 341395 309843 341398
rect 141417 341050 141483 341053
rect 142061 341050 142127 341053
rect 157333 341050 157399 341053
rect 141417 341048 157399 341050
rect 141417 340992 141422 341048
rect 141478 340992 142066 341048
rect 142122 340992 157338 341048
rect 157394 340992 157399 341048
rect 141417 340990 157399 340992
rect 141417 340987 141483 340990
rect 142061 340987 142127 340990
rect 157333 340987 157399 340990
rect 71773 340914 71839 340917
rect 73061 340914 73127 340917
rect 189901 340914 189967 340917
rect 71773 340912 189967 340914
rect 71773 340856 71778 340912
rect 71834 340856 73066 340912
rect 73122 340856 189906 340912
rect 189962 340856 189967 340912
rect 71773 340854 189967 340856
rect 71773 340851 71839 340854
rect 73061 340851 73127 340854
rect 189901 340851 189967 340854
rect 309777 340914 309843 340917
rect 311893 340914 311959 340917
rect 309777 340912 311959 340914
rect 309777 340856 309782 340912
rect 309838 340856 311898 340912
rect 311954 340856 311959 340912
rect 309777 340854 311959 340856
rect 309777 340851 309843 340854
rect 311893 340851 311959 340854
rect 93209 340098 93275 340101
rect 94446 340098 94452 340100
rect 93209 340096 94452 340098
rect 93209 340040 93214 340096
rect 93270 340040 94452 340096
rect 93209 340038 94452 340040
rect 93209 340035 93275 340038
rect 94446 340036 94452 340038
rect 94516 340098 94522 340100
rect 184289 340098 184355 340101
rect 94516 340096 184355 340098
rect 94516 340040 184294 340096
rect 184350 340040 184355 340096
rect 94516 340038 184355 340040
rect 94516 340036 94522 340038
rect 184289 340035 184355 340038
rect 134609 339690 134675 339693
rect 139393 339690 139459 339693
rect 173157 339690 173223 339693
rect 134609 339688 173223 339690
rect 134609 339632 134614 339688
rect 134670 339632 139398 339688
rect 139454 339632 173162 339688
rect 173218 339632 173223 339688
rect 134609 339630 173223 339632
rect 134609 339627 134675 339630
rect 139393 339627 139459 339630
rect 173157 339627 173223 339630
rect 90909 339554 90975 339557
rect 274081 339554 274147 339557
rect 90909 339552 274147 339554
rect 90909 339496 90914 339552
rect 90970 339496 274086 339552
rect 274142 339496 274147 339552
rect 90909 339494 274147 339496
rect 90909 339491 90975 339494
rect 274081 339491 274147 339494
rect 193949 338738 194015 338741
rect 207749 338738 207815 338741
rect 193949 338736 207815 338738
rect 193949 338680 193954 338736
rect 194010 338680 207754 338736
rect 207810 338680 207815 338736
rect 193949 338678 207815 338680
rect 193949 338675 194015 338678
rect 207749 338675 207815 338678
rect 211889 338738 211955 338741
rect 280889 338738 280955 338741
rect 211889 338736 280955 338738
rect 211889 338680 211894 338736
rect 211950 338680 280894 338736
rect 280950 338680 280955 338736
rect 211889 338678 280955 338680
rect 211889 338675 211955 338678
rect 280889 338675 280955 338678
rect 153837 338602 153903 338605
rect 142110 338600 153903 338602
rect 142110 338544 153842 338600
rect 153898 338544 153903 338600
rect 142110 338542 153903 338544
rect 109534 338404 109540 338468
rect 109604 338466 109610 338468
rect 109677 338466 109743 338469
rect 142110 338466 142170 338542
rect 153837 338539 153903 338542
rect 109604 338464 142170 338466
rect 109604 338408 109682 338464
rect 109738 338408 142170 338464
rect 109604 338406 142170 338408
rect 154481 338466 154547 338469
rect 172421 338466 172487 338469
rect 173198 338466 173204 338468
rect 154481 338464 173204 338466
rect 154481 338408 154486 338464
rect 154542 338408 172426 338464
rect 172482 338408 173204 338464
rect 154481 338406 173204 338408
rect 109604 338404 109610 338406
rect 109677 338403 109743 338406
rect 154481 338403 154547 338406
rect 172421 338403 172487 338406
rect 173198 338404 173204 338406
rect 173268 338404 173274 338468
rect 583520 338452 584960 338692
rect 61745 338330 61811 338333
rect 167637 338330 167703 338333
rect 61745 338328 167703 338330
rect 61745 338272 61750 338328
rect 61806 338272 167642 338328
rect 167698 338272 167703 338328
rect 61745 338270 167703 338272
rect 61745 338267 61811 338270
rect 167637 338267 167703 338270
rect 60457 338194 60523 338197
rect 62757 338194 62823 338197
rect 195329 338194 195395 338197
rect 60457 338192 195395 338194
rect 60457 338136 60462 338192
rect 60518 338136 62762 338192
rect 62818 338136 195334 338192
rect 195390 338136 195395 338192
rect 60457 338134 195395 338136
rect 60457 338131 60523 338134
rect 62757 338131 62823 338134
rect 195329 338131 195395 338134
rect 154021 338058 154087 338061
rect 157977 338058 158043 338061
rect 154021 338056 158043 338058
rect 154021 338000 154026 338056
rect 154082 338000 157982 338056
rect 158038 338000 158043 338056
rect 154021 337998 158043 338000
rect 154021 337995 154087 337998
rect 157977 337995 158043 337998
rect 157333 337378 157399 337381
rect 170254 337378 170260 337380
rect 157333 337376 170260 337378
rect 157333 337320 157338 337376
rect 157394 337320 170260 337376
rect 157333 337318 170260 337320
rect 157333 337315 157399 337318
rect 170254 337316 170260 337318
rect 170324 337316 170330 337380
rect 195094 337316 195100 337380
rect 195164 337378 195170 337380
rect 326337 337378 326403 337381
rect 327717 337378 327783 337381
rect 195164 337376 327783 337378
rect 195164 337320 326342 337376
rect 326398 337320 327722 337376
rect 327778 337320 327783 337376
rect 195164 337318 327783 337320
rect 195164 337316 195170 337318
rect 326337 337315 326403 337318
rect 327717 337315 327783 337318
rect 67633 337242 67699 337245
rect 150525 337242 150591 337245
rect 67633 337240 150591 337242
rect 67633 337184 67638 337240
rect 67694 337184 150530 337240
rect 150586 337184 150591 337240
rect 67633 337182 150591 337184
rect 67633 337179 67699 337182
rect 150525 337179 150591 337182
rect 117221 337106 117287 337109
rect 153193 337106 153259 337109
rect 117221 337104 153259 337106
rect 117221 337048 117226 337104
rect 117282 337048 153198 337104
rect 153254 337048 153259 337104
rect 117221 337046 153259 337048
rect 117221 337043 117287 337046
rect 153193 337043 153259 337046
rect 150433 336970 150499 336973
rect 160093 336970 160159 336973
rect 150433 336968 160159 336970
rect 150433 336912 150438 336968
rect 150494 336912 160098 336968
rect 160154 336912 160159 336968
rect 150433 336910 160159 336912
rect 150433 336907 150499 336910
rect 160093 336907 160159 336910
rect 178677 336970 178743 336973
rect 182817 336970 182883 336973
rect 178677 336968 182883 336970
rect 178677 336912 178682 336968
rect 178738 336912 182822 336968
rect 182878 336912 182883 336968
rect 178677 336910 182883 336912
rect 178677 336907 178743 336910
rect 182817 336907 182883 336910
rect 72233 336834 72299 336837
rect 194041 336834 194107 336837
rect 72233 336832 194107 336834
rect 72233 336776 72238 336832
rect 72294 336776 194046 336832
rect 194102 336776 194107 336832
rect 72233 336774 194107 336776
rect 72233 336771 72299 336774
rect 194041 336771 194107 336774
rect 271873 336698 271939 336701
rect 272517 336698 272583 336701
rect 271873 336696 272583 336698
rect 271873 336640 271878 336696
rect 271934 336640 272522 336696
rect 272578 336640 272583 336696
rect 271873 336638 272583 336640
rect 271873 336635 271939 336638
rect 272517 336635 272583 336638
rect 97809 336154 97875 336157
rect 137277 336154 137343 336157
rect 97809 336152 137343 336154
rect 97809 336096 97814 336152
rect 97870 336096 137282 336152
rect 137338 336096 137343 336152
rect 97809 336094 137343 336096
rect 97809 336091 97875 336094
rect 137277 336091 137343 336094
rect 57605 336018 57671 336021
rect 150433 336018 150499 336021
rect 57605 336016 150499 336018
rect 57605 335960 57610 336016
rect 57666 335960 150438 336016
rect 150494 335960 150499 336016
rect 57605 335958 150499 335960
rect 57605 335955 57671 335958
rect 150433 335955 150499 335958
rect 178861 336018 178927 336021
rect 188838 336018 188844 336020
rect 178861 336016 188844 336018
rect 178861 335960 178866 336016
rect 178922 335960 188844 336016
rect 178861 335958 188844 335960
rect 178861 335955 178927 335958
rect 188838 335956 188844 335958
rect 188908 336018 188914 336020
rect 582373 336018 582439 336021
rect 188908 336016 582439 336018
rect 188908 335960 582378 336016
rect 582434 335960 582439 336016
rect 188908 335958 582439 335960
rect 188908 335956 188914 335958
rect 582373 335955 582439 335958
rect 151905 335746 151971 335749
rect 153101 335746 153167 335749
rect 159398 335746 159404 335748
rect 151905 335744 159404 335746
rect 151905 335688 151910 335744
rect 151966 335688 153106 335744
rect 153162 335688 159404 335744
rect 151905 335686 159404 335688
rect 151905 335683 151971 335686
rect 153101 335683 153167 335686
rect 159398 335684 159404 335686
rect 159468 335684 159474 335748
rect 124213 335610 124279 335613
rect 177481 335610 177547 335613
rect 124213 335608 177547 335610
rect 124213 335552 124218 335608
rect 124274 335552 177486 335608
rect 177542 335552 177547 335608
rect 124213 335550 177547 335552
rect 124213 335547 124279 335550
rect 177481 335547 177547 335550
rect 21357 335474 21423 335477
rect 124949 335474 125015 335477
rect 21357 335472 125015 335474
rect 21357 335416 21362 335472
rect 21418 335416 124954 335472
rect 125010 335416 125015 335472
rect 21357 335414 125015 335416
rect 21357 335411 21423 335414
rect 124949 335411 125015 335414
rect 139209 335474 139275 335477
rect 271873 335474 271939 335477
rect 139209 335472 271939 335474
rect 139209 335416 139214 335472
rect 139270 335416 271878 335472
rect 271934 335416 271939 335472
rect 139209 335414 271939 335416
rect 139209 335411 139275 335414
rect 271873 335411 271939 335414
rect 160093 334794 160159 334797
rect 245653 334794 245719 334797
rect 160093 334792 245719 334794
rect 160093 334736 160098 334792
rect 160154 334736 245658 334792
rect 245714 334736 245719 334792
rect 160093 334734 245719 334736
rect 160093 334731 160159 334734
rect 245653 334731 245719 334734
rect 58985 334658 59051 334661
rect 129181 334658 129247 334661
rect 58985 334656 129247 334658
rect 58985 334600 58990 334656
rect 59046 334600 129186 334656
rect 129242 334600 129247 334656
rect 58985 334598 129247 334600
rect 58985 334595 59051 334598
rect 129181 334595 129247 334598
rect 153193 334658 153259 334661
rect 247033 334658 247099 334661
rect 153193 334656 247099 334658
rect 153193 334600 153198 334656
rect 153254 334600 247038 334656
rect 247094 334600 247099 334656
rect 153193 334598 247099 334600
rect 153193 334595 153259 334598
rect 247033 334595 247099 334598
rect 150433 334522 150499 334525
rect 160829 334522 160895 334525
rect 150433 334520 160895 334522
rect 150433 334464 150438 334520
rect 150494 334464 160834 334520
rect 160890 334464 160895 334520
rect 150433 334462 160895 334464
rect 150433 334459 150499 334462
rect 160829 334459 160895 334462
rect 146201 334250 146267 334253
rect 159633 334250 159699 334253
rect 146201 334248 159699 334250
rect 146201 334192 146206 334248
rect 146262 334192 159638 334248
rect 159694 334192 159699 334248
rect 146201 334190 159699 334192
rect 146201 334187 146267 334190
rect 159633 334187 159699 334190
rect 106641 334114 106707 334117
rect 150433 334114 150499 334117
rect 106641 334112 150499 334114
rect 106641 334056 106646 334112
rect 106702 334056 150438 334112
rect 150494 334056 150499 334112
rect 106641 334054 150499 334056
rect 106641 334051 106707 334054
rect 150433 334051 150499 334054
rect 157977 333434 158043 333437
rect 241646 333434 241652 333436
rect 157977 333432 241652 333434
rect 157977 333376 157982 333432
rect 158038 333376 241652 333432
rect 157977 333374 241652 333376
rect 157977 333371 158043 333374
rect 241646 333372 241652 333374
rect 241716 333372 241722 333436
rect 73245 333298 73311 333301
rect 73981 333298 74047 333301
rect 75177 333298 75243 333301
rect 73245 333296 75243 333298
rect 73245 333240 73250 333296
rect 73306 333240 73986 333296
rect 74042 333240 75182 333296
rect 75238 333240 75243 333296
rect 73245 333238 75243 333240
rect 73245 333235 73311 333238
rect 73981 333235 74047 333238
rect 75177 333235 75243 333238
rect 82997 333298 83063 333301
rect 109677 333298 109743 333301
rect 82997 333296 109743 333298
rect 82997 333240 83002 333296
rect 83058 333240 109682 333296
rect 109738 333240 109743 333296
rect 82997 333238 109743 333240
rect 82997 333235 83063 333238
rect 109677 333235 109743 333238
rect 110137 333298 110203 333301
rect 120717 333298 120783 333301
rect 110137 333296 120783 333298
rect 110137 333240 110142 333296
rect 110198 333240 120722 333296
rect 120778 333240 120783 333296
rect 110137 333238 120783 333240
rect 110137 333235 110203 333238
rect 120717 333235 120783 333238
rect 155217 333298 155283 333301
rect 582373 333298 582439 333301
rect 155217 333296 582439 333298
rect 155217 333240 155222 333296
rect 155278 333240 582378 333296
rect 582434 333240 582439 333296
rect 155217 333238 582439 333240
rect 155217 333235 155283 333238
rect 582373 333235 582439 333238
rect 107837 333026 107903 333029
rect 189717 333026 189783 333029
rect 107837 333024 189783 333026
rect 107837 332968 107842 333024
rect 107898 332968 189722 333024
rect 189778 332968 189783 333024
rect 107837 332966 189783 332968
rect 107837 332963 107903 332966
rect 189717 332963 189783 332966
rect 124857 332890 124923 332893
rect 125409 332890 125475 332893
rect 153101 332890 153167 332893
rect 124857 332888 153167 332890
rect 124857 332832 124862 332888
rect 124918 332832 125414 332888
rect 125470 332832 153106 332888
rect 153162 332832 153167 332888
rect 124857 332830 153167 332832
rect 124857 332827 124923 332830
rect 125409 332827 125475 332830
rect 153101 332827 153167 332830
rect 121821 332754 121887 332757
rect 158161 332754 158227 332757
rect 121821 332752 158227 332754
rect 121821 332696 121826 332752
rect 121882 332696 158166 332752
rect 158222 332696 158227 332752
rect 121821 332694 158227 332696
rect 121821 332691 121887 332694
rect 158161 332691 158227 332694
rect 59077 332618 59143 332621
rect 73245 332618 73311 332621
rect 59077 332616 73311 332618
rect 59077 332560 59082 332616
rect 59138 332560 73250 332616
rect 73306 332560 73311 332616
rect 59077 332558 73311 332560
rect 59077 332555 59143 332558
rect 73245 332555 73311 332558
rect 152457 332482 152523 332485
rect 155309 332482 155375 332485
rect 152457 332480 155375 332482
rect -960 332196 480 332436
rect 152457 332424 152462 332480
rect 152518 332424 155314 332480
rect 155370 332424 155375 332480
rect 152457 332422 155375 332424
rect 152457 332419 152523 332422
rect 155309 332419 155375 332422
rect 75177 332346 75243 332349
rect 75821 332346 75887 332349
rect 75177 332344 75887 332346
rect 75177 332288 75182 332344
rect 75238 332288 75826 332344
rect 75882 332288 75887 332344
rect 75177 332286 75887 332288
rect 75177 332283 75243 332286
rect 75821 332283 75887 332286
rect 62021 331938 62087 331941
rect 84101 331938 84167 331941
rect 62021 331936 84167 331938
rect 62021 331880 62026 331936
rect 62082 331880 84106 331936
rect 84162 331880 84167 331936
rect 62021 331878 84167 331880
rect 62021 331875 62087 331878
rect 84101 331875 84167 331878
rect 142061 331938 142127 331941
rect 146201 331938 146267 331941
rect 142061 331936 146267 331938
rect 142061 331880 142066 331936
rect 142122 331880 146206 331936
rect 146262 331880 146267 331936
rect 142061 331878 146267 331880
rect 142061 331875 142127 331878
rect 146201 331875 146267 331878
rect 153101 331938 153167 331941
rect 164785 331938 164851 331941
rect 153101 331936 164851 331938
rect 153101 331880 153106 331936
rect 153162 331880 164790 331936
rect 164846 331880 164851 331936
rect 153101 331878 164851 331880
rect 153101 331875 153167 331878
rect 164785 331875 164851 331878
rect 178534 331876 178540 331940
rect 178604 331938 178610 331940
rect 189809 331938 189875 331941
rect 178604 331936 189875 331938
rect 178604 331880 189814 331936
rect 189870 331880 189875 331936
rect 178604 331878 189875 331880
rect 178604 331876 178610 331878
rect 189809 331875 189875 331878
rect 69841 331802 69907 331805
rect 151905 331802 151971 331805
rect 69841 331800 151971 331802
rect 69841 331744 69846 331800
rect 69902 331744 151910 331800
rect 151966 331744 151971 331800
rect 69841 331742 151971 331744
rect 69841 331739 69907 331742
rect 151905 331739 151971 331742
rect 154849 331802 154915 331805
rect 155769 331802 155835 331805
rect 154849 331800 155835 331802
rect 154849 331744 154854 331800
rect 154910 331744 155774 331800
rect 155830 331744 155835 331800
rect 154849 331742 155835 331744
rect 154849 331739 154915 331742
rect 155769 331739 155835 331742
rect 163589 331802 163655 331805
rect 262305 331802 262371 331805
rect 163589 331800 262371 331802
rect 163589 331744 163594 331800
rect 163650 331744 262310 331800
rect 262366 331744 262371 331800
rect 163589 331742 262371 331744
rect 163589 331739 163655 331742
rect 262305 331739 262371 331742
rect 155769 331394 155835 331397
rect 162158 331394 162164 331396
rect 155769 331392 162164 331394
rect 155769 331336 155774 331392
rect 155830 331336 162164 331392
rect 155769 331334 162164 331336
rect 155769 331331 155835 331334
rect 162158 331332 162164 331334
rect 162228 331332 162234 331396
rect 149697 331258 149763 331261
rect 150249 331258 150315 331261
rect 180425 331258 180491 331261
rect 149697 331256 180491 331258
rect 149697 331200 149702 331256
rect 149758 331200 150254 331256
rect 150310 331200 180430 331256
rect 180486 331200 180491 331256
rect 149697 331198 180491 331200
rect 149697 331195 149763 331198
rect 150249 331195 150315 331198
rect 180425 331195 180491 331198
rect 129733 331122 129799 331125
rect 153193 331122 153259 331125
rect 129733 331120 153259 331122
rect 129733 331064 129738 331120
rect 129794 331064 153198 331120
rect 153254 331064 153259 331120
rect 129733 331062 153259 331064
rect 129733 331059 129799 331062
rect 153193 331059 153259 331062
rect 153837 330578 153903 330581
rect 157926 330578 157932 330580
rect 153837 330576 157932 330578
rect 153837 330520 153842 330576
rect 153898 330520 157932 330576
rect 153837 330518 157932 330520
rect 153837 330515 153903 330518
rect 157926 330516 157932 330518
rect 157996 330516 158002 330580
rect 216029 330578 216095 330581
rect 252502 330578 252508 330580
rect 216029 330576 252508 330578
rect 216029 330520 216034 330576
rect 216090 330520 252508 330576
rect 216029 330518 252508 330520
rect 216029 330515 216095 330518
rect 252502 330516 252508 330518
rect 252572 330516 252578 330580
rect 145281 330442 145347 330445
rect 242249 330442 242315 330445
rect 145281 330440 242315 330442
rect 145281 330384 145286 330440
rect 145342 330384 242254 330440
rect 242310 330384 242315 330440
rect 145281 330382 242315 330384
rect 145281 330379 145347 330382
rect 242249 330379 242315 330382
rect 39297 330034 39363 330037
rect 125409 330034 125475 330037
rect 39297 330032 125475 330034
rect 39297 329976 39302 330032
rect 39358 329976 125414 330032
rect 125470 329976 125475 330032
rect 39297 329974 125475 329976
rect 39297 329971 39363 329974
rect 125409 329971 125475 329974
rect 154113 330034 154179 330037
rect 156822 330034 156828 330036
rect 154113 330032 156828 330034
rect 154113 329976 154118 330032
rect 154174 329976 156828 330032
rect 154113 329974 156828 329976
rect 154113 329971 154179 329974
rect 156822 329972 156828 329974
rect 156892 329972 156898 330036
rect 7557 329898 7623 329901
rect 126237 329898 126303 329901
rect 7557 329896 126303 329898
rect 7557 329840 7562 329896
rect 7618 329840 126242 329896
rect 126298 329840 126303 329896
rect 7557 329838 126303 329840
rect 7557 329835 7623 329838
rect 126237 329835 126303 329838
rect 136449 329898 136515 329901
rect 145373 329898 145439 329901
rect 136449 329896 145439 329898
rect 136449 329840 136454 329896
rect 136510 329840 145378 329896
rect 145434 329840 145439 329896
rect 136449 329838 145439 329840
rect 136449 329835 136515 329838
rect 145373 329835 145439 329838
rect 155953 329898 156019 329901
rect 340137 329898 340203 329901
rect 155953 329896 340203 329898
rect 155953 329840 155958 329896
rect 156014 329840 340142 329896
rect 340198 329840 340203 329896
rect 155953 329838 340203 329840
rect 155953 329835 156019 329838
rect 340137 329835 340203 329838
rect 156873 329762 156939 329765
rect 162117 329762 162183 329765
rect 156873 329760 162183 329762
rect 156873 329704 156878 329760
rect 156934 329704 162122 329760
rect 162178 329704 162183 329760
rect 156873 329702 162183 329704
rect 156873 329699 156939 329702
rect 162117 329699 162183 329702
rect 69422 329564 69428 329628
rect 69492 329626 69498 329628
rect 72918 329626 72924 329628
rect 69492 329566 72924 329626
rect 69492 329564 69498 329566
rect 72918 329564 72924 329566
rect 72988 329564 72994 329628
rect 75177 329490 75243 329493
rect 75678 329490 75684 329492
rect 75177 329488 75684 329490
rect 75177 329432 75182 329488
rect 75238 329432 75684 329488
rect 75177 329430 75684 329432
rect 75177 329427 75243 329430
rect 75678 329428 75684 329430
rect 75748 329428 75754 329492
rect 70025 329354 70091 329357
rect 69430 329352 70091 329354
rect 69430 329296 70030 329352
rect 70086 329296 70091 329352
rect 69430 329294 70091 329296
rect 69430 328916 69490 329294
rect 70025 329291 70091 329294
rect 195237 329082 195303 329085
rect 258717 329082 258783 329085
rect 372705 329082 372771 329085
rect 195237 329080 372771 329082
rect 195237 329024 195242 329080
rect 195298 329024 258722 329080
rect 258778 329024 372710 329080
rect 372766 329024 372771 329080
rect 195237 329022 372771 329024
rect 195237 329019 195303 329022
rect 258717 329019 258783 329022
rect 372705 329019 372771 329022
rect 159725 328674 159791 328677
rect 232681 328674 232747 328677
rect 156676 328672 159791 328674
rect 156676 328616 159730 328672
rect 159786 328616 159791 328672
rect 156676 328614 159791 328616
rect 159725 328611 159791 328614
rect 161430 328672 232747 328674
rect 161430 328616 232686 328672
rect 232742 328616 232747 328672
rect 161430 328614 232747 328616
rect 156873 328538 156939 328541
rect 161430 328538 161490 328614
rect 232681 328611 232747 328614
rect 156873 328536 161490 328538
rect 156873 328480 156878 328536
rect 156934 328480 161490 328536
rect 156873 328478 161490 328480
rect 156873 328475 156939 328478
rect 69422 328340 69428 328404
rect 69492 328340 69498 328404
rect 244273 328402 244339 328405
rect 245009 328402 245075 328405
rect 244273 328400 245075 328402
rect 244273 328344 244278 328400
rect 244334 328344 245014 328400
rect 245070 328344 245075 328400
rect 244273 328342 245075 328344
rect 69430 327828 69490 328340
rect 244273 328339 244339 328342
rect 245009 328339 245075 328342
rect 156822 328204 156828 328268
rect 156892 328266 156898 328268
rect 162945 328266 163011 328269
rect 156892 328264 163011 328266
rect 156892 328208 162950 328264
rect 163006 328208 163011 328264
rect 156892 328206 163011 328208
rect 156892 328204 156898 328206
rect 162945 328203 163011 328206
rect 185669 327858 185735 327861
rect 209129 327858 209195 327861
rect 185669 327856 209195 327858
rect 185669 327800 185674 327856
rect 185730 327800 209134 327856
rect 209190 327800 209195 327856
rect 185669 327798 209195 327800
rect 185669 327795 185735 327798
rect 209129 327795 209195 327798
rect 156873 327722 156939 327725
rect 244273 327722 244339 327725
rect 156873 327720 244339 327722
rect 156873 327664 156878 327720
rect 156934 327664 244278 327720
rect 244334 327664 244339 327720
rect 156873 327662 244339 327664
rect 156873 327659 156939 327662
rect 244273 327659 244339 327662
rect 159541 327586 159607 327589
rect 156676 327584 159607 327586
rect 156676 327528 159546 327584
rect 159602 327528 159607 327584
rect 156676 327526 159607 327528
rect 159541 327523 159607 327526
rect 66253 326770 66319 326773
rect 66253 326768 68908 326770
rect 66253 326712 66258 326768
rect 66314 326712 68908 326768
rect 66253 326710 68908 326712
rect 66253 326707 66319 326710
rect 158713 326498 158779 326501
rect 156676 326496 158779 326498
rect 156676 326440 158718 326496
rect 158774 326440 158779 326496
rect 156676 326438 158779 326440
rect 158713 326435 158779 326438
rect 172053 326362 172119 326365
rect 191598 326362 191604 326364
rect 172053 326360 191604 326362
rect 172053 326304 172058 326360
rect 172114 326304 191604 326360
rect 172053 326302 191604 326304
rect 172053 326299 172119 326302
rect 191598 326300 191604 326302
rect 191668 326362 191674 326364
rect 282177 326362 282243 326365
rect 191668 326360 282243 326362
rect 191668 326304 282182 326360
rect 282238 326304 282243 326360
rect 191668 326302 282243 326304
rect 191668 326300 191674 326302
rect 282177 326299 282243 326302
rect 69430 325548 69490 325652
rect 69422 325484 69428 325548
rect 69492 325484 69498 325548
rect 157742 325410 157748 325412
rect 156676 325350 157748 325410
rect 157742 325348 157748 325350
rect 157812 325348 157818 325412
rect 583017 325274 583083 325277
rect 583520 325274 584960 325364
rect 583017 325272 584960 325274
rect 583017 325216 583022 325272
rect 583078 325216 584960 325272
rect 583017 325214 584960 325216
rect 583017 325211 583083 325214
rect 583520 325124 584960 325214
rect 159633 325002 159699 325005
rect 238109 325002 238175 325005
rect 159633 325000 238175 325002
rect 159633 324944 159638 325000
rect 159694 324944 238114 325000
rect 238170 324944 238175 325000
rect 159633 324942 238175 324944
rect 159633 324939 159699 324942
rect 238109 324939 238175 324942
rect 246297 325002 246363 325005
rect 299473 325002 299539 325005
rect 246297 325000 299539 325002
rect 246297 324944 246302 325000
rect 246358 324944 299478 325000
rect 299534 324944 299539 325000
rect 246297 324942 299539 324944
rect 246297 324939 246363 324942
rect 299473 324939 299539 324942
rect 67265 324594 67331 324597
rect 67265 324592 68908 324594
rect 67265 324536 67270 324592
rect 67326 324536 68908 324592
rect 67265 324534 68908 324536
rect 67265 324531 67331 324534
rect 157742 324396 157748 324460
rect 157812 324458 157818 324460
rect 158897 324458 158963 324461
rect 157812 324456 158963 324458
rect 157812 324400 158902 324456
rect 158958 324400 158963 324456
rect 157812 324398 158963 324400
rect 157812 324396 157818 324398
rect 158897 324395 158963 324398
rect 158713 324322 158779 324325
rect 156676 324320 158779 324322
rect 156676 324264 158718 324320
rect 158774 324264 158779 324320
rect 156676 324262 158779 324264
rect 158713 324259 158779 324262
rect 176101 323778 176167 323781
rect 220854 323778 220860 323780
rect 176101 323776 220860 323778
rect 176101 323720 176106 323776
rect 176162 323720 220860 323776
rect 176101 323718 220860 323720
rect 176101 323715 176167 323718
rect 220854 323716 220860 323718
rect 220924 323716 220930 323780
rect 233877 323778 233943 323781
rect 247718 323778 247724 323780
rect 233877 323776 247724 323778
rect 233877 323720 233882 323776
rect 233938 323720 247724 323776
rect 233877 323718 247724 323720
rect 233877 323715 233943 323718
rect 247718 323716 247724 323718
rect 247788 323716 247794 323780
rect 159725 323642 159791 323645
rect 371325 323642 371391 323645
rect 159725 323640 371391 323642
rect 159725 323584 159730 323640
rect 159786 323584 371330 323640
rect 371386 323584 371391 323640
rect 159725 323582 371391 323584
rect 159725 323579 159791 323582
rect 371325 323579 371391 323582
rect 67817 323506 67883 323509
rect 67817 323504 68908 323506
rect 67817 323448 67822 323504
rect 67878 323448 68908 323504
rect 67817 323446 68908 323448
rect 67817 323443 67883 323446
rect 158805 323234 158871 323237
rect 156676 323232 158871 323234
rect 156676 323176 158810 323232
rect 158866 323176 158871 323232
rect 156676 323174 158871 323176
rect 158805 323171 158871 323174
rect 66529 322418 66595 322421
rect 66529 322416 68908 322418
rect 66529 322360 66534 322416
rect 66590 322360 68908 322416
rect 66529 322358 68908 322360
rect 66529 322355 66595 322358
rect 158713 322146 158779 322149
rect 156676 322144 158779 322146
rect 156676 322088 158718 322144
rect 158774 322088 158779 322144
rect 156676 322086 158779 322088
rect 158713 322083 158779 322086
rect 235993 322146 236059 322149
rect 259453 322146 259519 322149
rect 235993 322144 259519 322146
rect 235993 322088 235998 322144
rect 236054 322088 259458 322144
rect 259514 322088 259519 322144
rect 235993 322086 259519 322088
rect 235993 322083 236059 322086
rect 259453 322083 259519 322086
rect 173709 321602 173775 321605
rect 284937 321602 285003 321605
rect 173709 321600 285003 321602
rect 173709 321544 173714 321600
rect 173770 321544 284942 321600
rect 284998 321544 285003 321600
rect 173709 321542 285003 321544
rect 173709 321539 173775 321542
rect 284937 321539 285003 321542
rect 68878 320650 68938 321300
rect 158713 321058 158779 321061
rect 156676 321056 158779 321058
rect 156676 321000 158718 321056
rect 158774 321000 158779 321056
rect 156676 320998 158779 321000
rect 158713 320995 158779 320998
rect 188337 320922 188403 320925
rect 221457 320922 221523 320925
rect 188337 320920 221523 320922
rect 188337 320864 188342 320920
rect 188398 320864 221462 320920
rect 221518 320864 221523 320920
rect 188337 320862 221523 320864
rect 188337 320859 188403 320862
rect 221457 320859 221523 320862
rect 158897 320786 158963 320789
rect 267733 320786 267799 320789
rect 158897 320784 267799 320786
rect 158897 320728 158902 320784
rect 158958 320728 267738 320784
rect 267794 320728 267799 320784
rect 158897 320726 267799 320728
rect 158897 320723 158963 320726
rect 267733 320723 267799 320726
rect 64830 320590 68938 320650
rect 232221 320650 232287 320653
rect 232681 320650 232747 320653
rect 232221 320648 232747 320650
rect 232221 320592 232226 320648
rect 232282 320592 232686 320648
rect 232742 320592 232747 320648
rect 232221 320590 232747 320592
rect 55070 320180 55076 320244
rect 55140 320242 55146 320244
rect 64830 320242 64890 320590
rect 232221 320587 232287 320590
rect 232681 320587 232747 320590
rect 55140 320182 64890 320242
rect 66805 320242 66871 320245
rect 232681 320242 232747 320245
rect 281574 320242 281580 320244
rect 66805 320240 68908 320242
rect 66805 320184 66810 320240
rect 66866 320184 68908 320240
rect 66805 320182 68908 320184
rect 232681 320240 281580 320242
rect 232681 320184 232686 320240
rect 232742 320184 281580 320240
rect 232681 320182 281580 320184
rect 55140 320180 55146 320182
rect 66805 320179 66871 320182
rect 232681 320179 232747 320182
rect 281574 320180 281580 320182
rect 281644 320180 281650 320244
rect 179413 320106 179479 320109
rect 180241 320106 180307 320109
rect 179413 320104 180307 320106
rect 179413 320048 179418 320104
rect 179474 320048 180246 320104
rect 180302 320048 180307 320104
rect 179413 320046 180307 320048
rect 179413 320043 179479 320046
rect 180241 320043 180307 320046
rect -960 319290 480 319380
rect 4061 319290 4127 319293
rect -960 319288 4127 319290
rect -960 319232 4066 319288
rect 4122 319232 4127 319288
rect -960 319230 4127 319232
rect -960 319140 480 319230
rect 4061 319227 4127 319230
rect 66437 319154 66503 319157
rect 156646 319154 156706 319940
rect 196617 319426 196683 319429
rect 226977 319426 227043 319429
rect 196617 319424 227043 319426
rect 196617 319368 196622 319424
rect 196678 319368 226982 319424
rect 227038 319368 227043 319424
rect 196617 319366 227043 319368
rect 196617 319363 196683 319366
rect 226977 319363 227043 319366
rect 158713 319154 158779 319157
rect 66437 319152 68908 319154
rect 66437 319096 66442 319152
rect 66498 319096 68908 319152
rect 66437 319094 68908 319096
rect 156646 319152 161490 319154
rect 156646 319096 158718 319152
rect 158774 319096 161490 319152
rect 156646 319094 161490 319096
rect 66437 319091 66503 319094
rect 158713 319091 158779 319094
rect 158805 318882 158871 318885
rect 156676 318880 158871 318882
rect 156676 318824 158810 318880
rect 158866 318824 158871 318880
rect 156676 318822 158871 318824
rect 161430 318882 161490 319094
rect 180241 318882 180307 318885
rect 161430 318880 180307 318882
rect 161430 318824 180246 318880
rect 180302 318824 180307 318880
rect 161430 318822 180307 318824
rect 158805 318819 158871 318822
rect 180241 318819 180307 318822
rect 197997 318882 198063 318885
rect 198406 318882 198412 318884
rect 197997 318880 198412 318882
rect 197997 318824 198002 318880
rect 198058 318824 198412 318880
rect 197997 318822 198412 318824
rect 197997 318819 198063 318822
rect 198406 318820 198412 318822
rect 198476 318882 198482 318884
rect 264237 318882 264303 318885
rect 198476 318880 264303 318882
rect 198476 318824 264242 318880
rect 264298 318824 264303 318880
rect 198476 318822 264303 318824
rect 198476 318820 198482 318822
rect 264237 318819 264303 318822
rect 164877 318746 164943 318749
rect 166993 318746 167059 318749
rect 164877 318744 167059 318746
rect 164877 318688 164882 318744
rect 164938 318688 166998 318744
rect 167054 318688 167059 318744
rect 164877 318686 167059 318688
rect 164877 318683 164943 318686
rect 166993 318683 167059 318686
rect 184289 318746 184355 318749
rect 184841 318746 184907 318749
rect 184289 318744 184907 318746
rect 184289 318688 184294 318744
rect 184350 318688 184846 318744
rect 184902 318688 184907 318744
rect 184289 318686 184907 318688
rect 184289 318683 184355 318686
rect 184841 318683 184907 318686
rect 66437 318066 66503 318069
rect 66437 318064 68908 318066
rect 66437 318008 66442 318064
rect 66498 318008 68908 318064
rect 66437 318006 68908 318008
rect 66437 318003 66503 318006
rect 161565 317794 161631 317797
rect 156676 317792 161631 317794
rect 156676 317736 161570 317792
rect 161626 317736 161631 317792
rect 156676 317734 161631 317736
rect 161565 317731 161631 317734
rect 198089 317658 198155 317661
rect 271229 317658 271295 317661
rect 198089 317656 271295 317658
rect 198089 317600 198094 317656
rect 198150 317600 271234 317656
rect 271290 317600 271295 317656
rect 198089 317598 271295 317600
rect 198089 317595 198155 317598
rect 271229 317595 271295 317598
rect 184841 317522 184907 317525
rect 427813 317522 427879 317525
rect 184841 317520 427879 317522
rect 184841 317464 184846 317520
rect 184902 317464 427818 317520
rect 427874 317464 427879 317520
rect 184841 317462 427879 317464
rect 184841 317459 184907 317462
rect 427813 317459 427879 317462
rect 164877 317386 164943 317389
rect 170397 317386 170463 317389
rect 164877 317384 170463 317386
rect 164877 317328 164882 317384
rect 164938 317328 170402 317384
rect 170458 317328 170463 317384
rect 164877 317326 170463 317328
rect 164877 317323 164943 317326
rect 170397 317323 170463 317326
rect 210969 317386 211035 317389
rect 340873 317386 340939 317389
rect 210969 317384 340939 317386
rect 210969 317328 210974 317384
rect 211030 317328 340878 317384
rect 340934 317328 340939 317384
rect 210969 317326 340939 317328
rect 210969 317323 211035 317326
rect 340873 317323 340939 317326
rect 66897 316978 66963 316981
rect 66897 316976 68908 316978
rect 66897 316920 66902 316976
rect 66958 316920 68908 316976
rect 66897 316918 68908 316920
rect 66897 316915 66963 316918
rect 174629 316842 174695 316845
rect 191046 316842 191052 316844
rect 174629 316840 191052 316842
rect 174629 316784 174634 316840
rect 174690 316784 191052 316840
rect 174629 316782 191052 316784
rect 174629 316779 174695 316782
rect 191046 316780 191052 316782
rect 191116 316780 191122 316844
rect 160001 316706 160067 316709
rect 156676 316704 160067 316706
rect 156676 316648 160006 316704
rect 160062 316648 160067 316704
rect 156676 316646 160067 316648
rect 160001 316643 160067 316646
rect 183185 316706 183251 316709
rect 227437 316706 227503 316709
rect 183185 316704 227503 316706
rect 183185 316648 183190 316704
rect 183246 316648 227442 316704
rect 227498 316648 227503 316704
rect 183185 316646 227503 316648
rect 183185 316643 183251 316646
rect 227437 316643 227503 316646
rect 227437 316162 227503 316165
rect 403617 316162 403683 316165
rect 227437 316160 403683 316162
rect 227437 316104 227442 316160
rect 227498 316104 403622 316160
rect 403678 316104 403683 316160
rect 227437 316102 403683 316104
rect 227437 316099 227503 316102
rect 403617 316099 403683 316102
rect 65926 315828 65932 315892
rect 65996 315890 66002 315892
rect 65996 315830 68908 315890
rect 65996 315828 66002 315830
rect 158805 315618 158871 315621
rect 156676 315616 158871 315618
rect 156676 315560 158810 315616
rect 158866 315560 158871 315616
rect 156676 315558 158871 315560
rect 158805 315555 158871 315558
rect 206369 315346 206435 315349
rect 225689 315346 225755 315349
rect 206369 315344 225755 315346
rect 206369 315288 206374 315344
rect 206430 315288 225694 315344
rect 225750 315288 225755 315344
rect 206369 315286 225755 315288
rect 206369 315283 206435 315286
rect 225689 315283 225755 315286
rect 242934 315012 242940 315076
rect 243004 315074 243010 315076
rect 244273 315074 244339 315077
rect 243004 315072 244339 315074
rect 243004 315016 244278 315072
rect 244334 315016 244339 315072
rect 243004 315014 244339 315016
rect 243004 315012 243010 315014
rect 244273 315011 244339 315014
rect 213177 314938 213243 314941
rect 287053 314938 287119 314941
rect 213177 314936 287119 314938
rect 213177 314880 213182 314936
rect 213238 314880 287058 314936
rect 287114 314880 287119 314936
rect 213177 314878 287119 314880
rect 213177 314875 213243 314878
rect 287053 314875 287119 314878
rect 66805 314802 66871 314805
rect 234613 314802 234679 314805
rect 235349 314802 235415 314805
rect 432597 314802 432663 314805
rect 66805 314800 68908 314802
rect 66805 314744 66810 314800
rect 66866 314744 68908 314800
rect 66805 314742 68908 314744
rect 234613 314800 432663 314802
rect 234613 314744 234618 314800
rect 234674 314744 235354 314800
rect 235410 314744 432602 314800
rect 432658 314744 432663 314800
rect 234613 314742 432663 314744
rect 66805 314739 66871 314742
rect 234613 314739 234679 314742
rect 235349 314739 235415 314742
rect 432597 314739 432663 314742
rect 66897 313986 66963 313989
rect 156646 313986 156706 314500
rect 196709 314122 196775 314125
rect 224166 314122 224172 314124
rect 196709 314120 224172 314122
rect 196709 314064 196714 314120
rect 196770 314064 224172 314120
rect 196709 314062 224172 314064
rect 196709 314059 196775 314062
rect 224166 314060 224172 314062
rect 224236 314060 224242 314124
rect 161381 313986 161447 313989
rect 244273 313986 244339 313989
rect 66897 313984 68908 313986
rect 66897 313928 66902 313984
rect 66958 313928 68908 313984
rect 66897 313926 68908 313928
rect 156646 313984 244339 313986
rect 156646 313928 161386 313984
rect 161442 313928 244278 313984
rect 244334 313928 244339 313984
rect 156646 313926 244339 313928
rect 66897 313923 66963 313926
rect 161381 313923 161447 313926
rect 244273 313923 244339 313926
rect 158805 313442 158871 313445
rect 156676 313440 158871 313442
rect 156676 313384 158810 313440
rect 158866 313384 158871 313440
rect 156676 313382 158871 313384
rect 158805 313379 158871 313382
rect 173249 313306 173315 313309
rect 173801 313306 173867 313309
rect 257337 313306 257403 313309
rect 173249 313304 257403 313306
rect 173249 313248 173254 313304
rect 173310 313248 173806 313304
rect 173862 313248 257342 313304
rect 257398 313248 257403 313304
rect 173249 313246 257403 313248
rect 173249 313243 173315 313246
rect 173801 313243 173867 313246
rect 257337 313243 257403 313246
rect 66161 312898 66227 312901
rect 66161 312896 68908 312898
rect 66161 312840 66166 312896
rect 66222 312840 68908 312896
rect 66161 312838 68908 312840
rect 66161 312835 66227 312838
rect 161238 312626 161244 312628
rect 156646 312566 161244 312626
rect 156646 312324 156706 312566
rect 161238 312564 161244 312566
rect 161308 312626 161314 312628
rect 262121 312626 262187 312629
rect 161308 312624 262187 312626
rect 161308 312568 262126 312624
rect 262182 312568 262187 312624
rect 161308 312566 262187 312568
rect 161308 312564 161314 312566
rect 262121 312563 262187 312566
rect 171041 312490 171107 312493
rect 182173 312490 182239 312493
rect 387057 312490 387123 312493
rect 171041 312488 387123 312490
rect 171041 312432 171046 312488
rect 171102 312432 182178 312488
rect 182234 312432 387062 312488
rect 387118 312432 387123 312488
rect 171041 312430 387123 312432
rect 171041 312427 171107 312430
rect 182173 312427 182239 312430
rect 387057 312427 387123 312430
rect 583293 312082 583359 312085
rect 583520 312082 584960 312172
rect 583293 312080 584960 312082
rect 583293 312024 583298 312080
rect 583354 312024 584960 312080
rect 583293 312022 584960 312024
rect 583293 312019 583359 312022
rect 583520 311932 584960 312022
rect 66989 311810 67055 311813
rect 66989 311808 68908 311810
rect 66989 311752 66994 311808
rect 67050 311752 68908 311808
rect 66989 311750 68908 311752
rect 66989 311747 67055 311750
rect 158897 311266 158963 311269
rect 156676 311264 158963 311266
rect 156676 311208 158902 311264
rect 158958 311208 158963 311264
rect 156676 311206 158963 311208
rect 158897 311203 158963 311206
rect 171961 311130 172027 311133
rect 204478 311130 204484 311132
rect 171961 311128 204484 311130
rect 171961 311072 171966 311128
rect 172022 311072 204484 311128
rect 171961 311070 204484 311072
rect 171961 311067 172027 311070
rect 204478 311068 204484 311070
rect 204548 311068 204554 311132
rect 244917 311130 244983 311133
rect 255405 311130 255471 311133
rect 244917 311128 255471 311130
rect 244917 311072 244922 311128
rect 244978 311072 255410 311128
rect 255466 311072 255471 311128
rect 244917 311070 255471 311072
rect 244917 311067 244983 311070
rect 255405 311067 255471 311070
rect 582833 310994 582899 310997
rect 583109 310994 583175 310997
rect 582833 310992 583175 310994
rect 582833 310936 582838 310992
rect 582894 310936 583114 310992
rect 583170 310936 583175 310992
rect 582833 310934 583175 310936
rect 582833 310931 582899 310934
rect 583109 310931 583175 310934
rect 67081 310722 67147 310725
rect 67081 310720 68908 310722
rect 67081 310664 67086 310720
rect 67142 310664 68908 310720
rect 67081 310662 68908 310664
rect 67081 310659 67147 310662
rect 210601 310586 210667 310589
rect 583109 310586 583175 310589
rect 210601 310584 583175 310586
rect 210601 310528 210606 310584
rect 210662 310528 583114 310584
rect 583170 310528 583175 310584
rect 210601 310526 583175 310528
rect 210601 310523 210667 310526
rect 583109 310523 583175 310526
rect 200113 310450 200179 310453
rect 180750 310448 200179 310450
rect 180750 310392 200118 310448
rect 200174 310392 200179 310448
rect 180750 310390 200179 310392
rect 158805 310178 158871 310181
rect 156676 310176 158871 310178
rect 156676 310120 158810 310176
rect 158866 310120 158871 310176
rect 156676 310118 158871 310120
rect 158805 310115 158871 310118
rect 160737 309906 160803 309909
rect 176653 309906 176719 309909
rect 180750 309906 180810 310390
rect 200070 310387 200179 310390
rect 282913 310450 282979 310453
rect 283557 310450 283623 310453
rect 352046 310450 352052 310452
rect 282913 310448 352052 310450
rect 282913 310392 282918 310448
rect 282974 310392 283562 310448
rect 283618 310392 352052 310448
rect 282913 310390 352052 310392
rect 282913 310387 282979 310390
rect 283557 310387 283623 310390
rect 352046 310388 352052 310390
rect 352116 310388 352122 310452
rect 200070 310042 200130 310387
rect 249149 310042 249215 310045
rect 200070 310040 249215 310042
rect 200070 309984 249154 310040
rect 249210 309984 249215 310040
rect 200070 309982 249215 309984
rect 249149 309979 249215 309982
rect 160737 309904 180810 309906
rect 160737 309848 160742 309904
rect 160798 309848 176658 309904
rect 176714 309848 180810 309904
rect 160737 309846 180810 309848
rect 160737 309843 160803 309846
rect 176653 309843 176719 309846
rect 224718 309844 224724 309908
rect 224788 309906 224794 309908
rect 285673 309906 285739 309909
rect 224788 309904 285739 309906
rect 224788 309848 285678 309904
rect 285734 309848 285739 309904
rect 224788 309846 285739 309848
rect 224788 309844 224794 309846
rect 285673 309843 285739 309846
rect 174813 309770 174879 309773
rect 239029 309770 239095 309773
rect 174813 309768 239095 309770
rect 174813 309712 174818 309768
rect 174874 309712 239034 309768
rect 239090 309712 239095 309768
rect 174813 309710 239095 309712
rect 174813 309707 174879 309710
rect 239029 309707 239095 309710
rect 66805 309634 66871 309637
rect 66805 309632 68908 309634
rect 66805 309576 66810 309632
rect 66866 309576 68908 309632
rect 66805 309574 68908 309576
rect 66805 309571 66871 309574
rect 179454 309090 179460 309092
rect 156676 309030 179460 309090
rect 179454 309028 179460 309030
rect 179524 309028 179530 309092
rect 214649 308682 214715 308685
rect 251214 308682 251220 308684
rect 214649 308680 251220 308682
rect 214649 308624 214654 308680
rect 214710 308624 251220 308680
rect 214649 308622 251220 308624
rect 214649 308619 214715 308622
rect 251214 308620 251220 308622
rect 251284 308620 251290 308684
rect 67725 308546 67791 308549
rect 67725 308544 68908 308546
rect 67725 308488 67730 308544
rect 67786 308488 68908 308544
rect 67725 308486 68908 308488
rect 67725 308483 67791 308486
rect 157926 308484 157932 308548
rect 157996 308546 158002 308548
rect 236637 308546 236703 308549
rect 157996 308544 236703 308546
rect 157996 308488 236642 308544
rect 236698 308488 236703 308544
rect 157996 308486 236703 308488
rect 157996 308484 158002 308486
rect 236637 308483 236703 308486
rect 179454 308348 179460 308412
rect 179524 308410 179530 308412
rect 180558 308410 180564 308412
rect 179524 308350 180564 308410
rect 179524 308348 179530 308350
rect 180558 308348 180564 308350
rect 180628 308410 180634 308412
rect 324957 308410 325023 308413
rect 180628 308408 325023 308410
rect 180628 308352 324962 308408
rect 325018 308352 325023 308408
rect 180628 308350 325023 308352
rect 180628 308348 180634 308350
rect 324957 308347 325023 308350
rect 158805 308002 158871 308005
rect 156676 308000 158871 308002
rect 156676 307944 158810 308000
rect 158866 307944 158871 308000
rect 156676 307942 158871 307944
rect 158805 307939 158871 307942
rect 177297 307730 177363 307733
rect 177573 307730 177639 307733
rect 177297 307728 177639 307730
rect 177297 307672 177302 307728
rect 177358 307672 177578 307728
rect 177634 307672 177639 307728
rect 177297 307670 177639 307672
rect 177297 307667 177363 307670
rect 177573 307667 177639 307670
rect 198365 307730 198431 307733
rect 198590 307730 198596 307732
rect 198365 307728 198596 307730
rect 198365 307672 198370 307728
rect 198426 307672 198596 307728
rect 198365 307670 198596 307672
rect 198365 307667 198431 307670
rect 198590 307668 198596 307670
rect 198660 307668 198666 307732
rect 66897 307458 66963 307461
rect 66897 307456 68908 307458
rect 66897 307400 66902 307456
rect 66958 307400 68908 307456
rect 66897 307398 68908 307400
rect 66897 307395 66963 307398
rect 159398 307124 159404 307188
rect 159468 307186 159474 307188
rect 188337 307186 188403 307189
rect 159468 307184 188403 307186
rect 159468 307128 188342 307184
rect 188398 307128 188403 307184
rect 159468 307126 188403 307128
rect 159468 307124 159474 307126
rect 188337 307123 188403 307126
rect 177573 307050 177639 307053
rect 213361 307050 213427 307053
rect 177573 307048 213427 307050
rect 177573 306992 177578 307048
rect 177634 306992 213366 307048
rect 213422 306992 213427 307048
rect 177573 306990 213427 306992
rect 177573 306987 177639 306990
rect 213361 306987 213427 306990
rect 220169 307050 220235 307053
rect 233734 307050 233740 307052
rect 220169 307048 233740 307050
rect 220169 306992 220174 307048
rect 220230 306992 233740 307048
rect 220169 306990 233740 306992
rect 220169 306987 220235 306990
rect 233734 306988 233740 306990
rect 233804 306988 233810 307052
rect 158805 306914 158871 306917
rect 156676 306912 158871 306914
rect 156676 306856 158810 306912
rect 158866 306856 158871 306912
rect 156676 306854 158871 306856
rect 158805 306851 158871 306854
rect 273989 306642 274055 306645
rect 200070 306640 274055 306642
rect 200070 306584 273994 306640
rect 274050 306584 274055 306640
rect 200070 306582 274055 306584
rect 198365 306506 198431 306509
rect 200070 306506 200130 306582
rect 273989 306579 274055 306582
rect 198365 306504 200130 306506
rect 198365 306448 198370 306504
rect 198426 306448 200130 306504
rect 198365 306446 200130 306448
rect 231117 306506 231183 306509
rect 352557 306506 352623 306509
rect 231117 306504 352623 306506
rect 231117 306448 231122 306504
rect 231178 306448 352562 306504
rect 352618 306448 352623 306504
rect 231117 306446 352623 306448
rect 198365 306443 198431 306446
rect 231117 306443 231183 306446
rect 352557 306443 352623 306446
rect 66805 306370 66871 306373
rect 66805 306368 68908 306370
rect -960 306234 480 306324
rect 66805 306312 66810 306368
rect 66866 306312 68908 306368
rect 66805 306310 68908 306312
rect 66805 306307 66871 306310
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 158805 305826 158871 305829
rect 156676 305824 158871 305826
rect 156676 305768 158810 305824
rect 158866 305768 158871 305824
rect 156676 305766 158871 305768
rect 158805 305763 158871 305766
rect 207657 305826 207723 305829
rect 215293 305826 215359 305829
rect 207657 305824 215359 305826
rect 207657 305768 207662 305824
rect 207718 305768 215298 305824
rect 215354 305768 215359 305824
rect 207657 305766 215359 305768
rect 207657 305763 207723 305766
rect 215293 305763 215359 305766
rect 182909 305690 182975 305693
rect 211429 305690 211495 305693
rect 182909 305688 211495 305690
rect 182909 305632 182914 305688
rect 182970 305632 211434 305688
rect 211490 305632 211495 305688
rect 182909 305630 211495 305632
rect 182909 305627 182975 305630
rect 211429 305627 211495 305630
rect 219198 305628 219204 305692
rect 219268 305690 219274 305692
rect 266997 305690 267063 305693
rect 219268 305688 267063 305690
rect 219268 305632 267002 305688
rect 267058 305632 267063 305688
rect 219268 305630 267063 305632
rect 219268 305628 219274 305630
rect 266997 305627 267063 305630
rect 65977 305282 66043 305285
rect 65977 305280 68908 305282
rect 65977 305224 65982 305280
rect 66038 305224 68908 305280
rect 65977 305222 68908 305224
rect 65977 305219 66043 305222
rect 201401 305010 201467 305013
rect 309133 305010 309199 305013
rect 310421 305010 310487 305013
rect 201401 305008 310487 305010
rect 201401 304952 201406 305008
rect 201462 304952 309138 305008
rect 309194 304952 310426 305008
rect 310482 304952 310487 305008
rect 201401 304950 310487 304952
rect 201401 304947 201467 304950
rect 309133 304947 309199 304950
rect 310421 304947 310487 304950
rect 158805 304738 158871 304741
rect 156676 304736 158871 304738
rect 156676 304680 158810 304736
rect 158866 304680 158871 304736
rect 156676 304678 158871 304680
rect 158805 304675 158871 304678
rect 67633 304194 67699 304197
rect 67633 304192 68908 304194
rect 67633 304136 67638 304192
rect 67694 304136 68908 304192
rect 67633 304134 68908 304136
rect 67633 304131 67699 304134
rect 211429 303786 211495 303789
rect 275277 303786 275343 303789
rect 211429 303784 275343 303786
rect 211429 303728 211434 303784
rect 211490 303728 275282 303784
rect 275338 303728 275343 303784
rect 211429 303726 275343 303728
rect 211429 303723 211495 303726
rect 275277 303723 275343 303726
rect 158805 303650 158871 303653
rect 156676 303648 158871 303650
rect 156676 303592 158810 303648
rect 158866 303592 158871 303648
rect 156676 303590 158871 303592
rect 158805 303587 158871 303590
rect 167637 303650 167703 303653
rect 237414 303650 237420 303652
rect 167637 303648 237420 303650
rect 167637 303592 167642 303648
rect 167698 303592 237420 303648
rect 167637 303590 237420 303592
rect 167637 303587 167703 303590
rect 237414 303588 237420 303590
rect 237484 303588 237490 303652
rect 66897 303106 66963 303109
rect 66897 303104 68908 303106
rect 66897 303048 66902 303104
rect 66958 303048 68908 303104
rect 66897 303046 68908 303048
rect 66897 303043 66963 303046
rect 156646 302290 156706 302532
rect 166257 302426 166323 302429
rect 250621 302426 250687 302429
rect 166257 302424 250687 302426
rect 166257 302368 166262 302424
rect 166318 302368 250626 302424
rect 250682 302368 250687 302424
rect 166257 302366 250687 302368
rect 166257 302363 166323 302366
rect 250621 302363 250687 302366
rect 304206 302290 304212 302292
rect 156646 302230 304212 302290
rect 304206 302228 304212 302230
rect 304276 302228 304282 302292
rect 66805 302018 66871 302021
rect 66805 302016 68908 302018
rect 66805 301960 66810 302016
rect 66866 301960 68908 302016
rect 66805 301958 68908 301960
rect 66805 301955 66871 301958
rect 195329 301746 195395 301749
rect 230289 301746 230355 301749
rect 195329 301744 230355 301746
rect 195329 301688 195334 301744
rect 195390 301688 230294 301744
rect 230350 301688 230355 301744
rect 195329 301686 230355 301688
rect 195329 301683 195395 301686
rect 230289 301683 230355 301686
rect 163589 301610 163655 301613
rect 169753 301610 169819 301613
rect 163589 301608 169819 301610
rect 163589 301552 163594 301608
rect 163650 301552 169758 301608
rect 169814 301552 169819 301608
rect 163589 301550 169819 301552
rect 163589 301547 163655 301550
rect 169753 301547 169819 301550
rect 217542 301548 217548 301612
rect 217612 301610 217618 301612
rect 262213 301610 262279 301613
rect 217612 301608 262279 301610
rect 217612 301552 262218 301608
rect 262274 301552 262279 301608
rect 217612 301550 262279 301552
rect 217612 301548 217618 301550
rect 262213 301547 262279 301550
rect 158805 301474 158871 301477
rect 156676 301472 158871 301474
rect 156676 301416 158810 301472
rect 158866 301416 158871 301472
rect 156676 301414 158871 301416
rect 158805 301411 158871 301414
rect 166073 301474 166139 301477
rect 258165 301474 258231 301477
rect 166073 301472 258231 301474
rect 166073 301416 166078 301472
rect 166134 301416 258170 301472
rect 258226 301416 258231 301472
rect 166073 301414 258231 301416
rect 166073 301411 166139 301414
rect 258165 301411 258231 301414
rect 66897 300930 66963 300933
rect 66897 300928 68908 300930
rect 66897 300872 66902 300928
rect 66958 300872 68908 300928
rect 66897 300870 68908 300872
rect 66897 300867 66963 300870
rect 158989 300386 159055 300389
rect 156676 300384 159055 300386
rect 156676 300328 158994 300384
rect 159050 300328 159055 300384
rect 156676 300326 159055 300328
rect 158989 300323 159055 300326
rect 158069 300114 158135 300117
rect 256785 300114 256851 300117
rect 158069 300112 256851 300114
rect 158069 300056 158074 300112
rect 158130 300056 256790 300112
rect 256846 300056 256851 300112
rect 158069 300054 256851 300056
rect 158069 300051 158135 300054
rect 256785 300051 256851 300054
rect 67541 299842 67607 299845
rect 67541 299840 68908 299842
rect 67541 299784 67546 299840
rect 67602 299784 68908 299840
rect 67541 299782 68908 299784
rect 67541 299779 67607 299782
rect 214741 299570 214807 299573
rect 267181 299570 267247 299573
rect 214741 299568 267247 299570
rect 214741 299512 214746 299568
rect 214802 299512 267186 299568
rect 267242 299512 267247 299568
rect 214741 299510 267247 299512
rect 214741 299507 214807 299510
rect 267181 299507 267247 299510
rect 66621 298754 66687 298757
rect 66621 298752 68908 298754
rect 66621 298696 66626 298752
rect 66682 298696 68908 298752
rect 66621 298694 68908 298696
rect 66621 298691 66687 298694
rect 156646 298618 156706 299268
rect 223021 298754 223087 298757
rect 279509 298754 279575 298757
rect 223021 298752 279575 298754
rect 223021 298696 223026 298752
rect 223082 298696 279514 298752
rect 279570 298696 279575 298752
rect 223021 298694 279575 298696
rect 223021 298691 223087 298694
rect 279509 298691 279575 298694
rect 582741 298754 582807 298757
rect 582925 298754 582991 298757
rect 583520 298754 584960 298844
rect 582741 298752 584960 298754
rect 582741 298696 582746 298752
rect 582802 298696 582930 298752
rect 582986 298696 584960 298752
rect 582741 298694 584960 298696
rect 582741 298691 582807 298694
rect 582925 298691 582991 298694
rect 156646 298558 161490 298618
rect 583520 298604 584960 298694
rect 161430 298346 161490 298558
rect 244406 298346 244412 298348
rect 161430 298286 244412 298346
rect 244406 298284 244412 298286
rect 244476 298284 244482 298348
rect 158805 298210 158871 298213
rect 156676 298208 158871 298210
rect 156676 298152 158810 298208
rect 158866 298152 158871 298208
rect 156676 298150 158871 298152
rect 158805 298147 158871 298150
rect 234521 298210 234587 298213
rect 322197 298210 322263 298213
rect 234521 298208 322263 298210
rect 234521 298152 234526 298208
rect 234582 298152 322202 298208
rect 322258 298152 322263 298208
rect 234521 298150 322263 298152
rect 234521 298147 234587 298150
rect 322197 298147 322263 298150
rect 168281 298074 168347 298077
rect 168465 298074 168531 298077
rect 168281 298072 168531 298074
rect 168281 298016 168286 298072
rect 168342 298016 168470 298072
rect 168526 298016 168531 298072
rect 168281 298014 168531 298016
rect 168281 298011 168347 298014
rect 168465 298011 168531 298014
rect 206461 298074 206527 298077
rect 207565 298074 207631 298077
rect 206461 298072 207631 298074
rect 206461 298016 206466 298072
rect 206522 298016 207570 298072
rect 207626 298016 207631 298072
rect 206461 298014 207631 298016
rect 206461 298011 206527 298014
rect 207565 298011 207631 298014
rect 254025 298074 254091 298077
rect 254577 298074 254643 298077
rect 254025 298072 254643 298074
rect 254025 298016 254030 298072
rect 254086 298016 254582 298072
rect 254638 298016 254643 298072
rect 254025 298014 254643 298016
rect 254025 298011 254091 298014
rect 254577 298011 254643 298014
rect 66805 297666 66871 297669
rect 66805 297664 68908 297666
rect 66805 297608 66810 297664
rect 66866 297608 68908 297664
rect 66805 297606 68908 297608
rect 66805 297603 66871 297606
rect 191097 297530 191163 297533
rect 206645 297530 206711 297533
rect 191097 297528 206711 297530
rect 191097 297472 191102 297528
rect 191158 297472 206650 297528
rect 206706 297472 206711 297528
rect 191097 297470 206711 297472
rect 191097 297467 191163 297470
rect 206645 297467 206711 297470
rect 208158 297468 208164 297532
rect 208228 297530 208234 297532
rect 226333 297530 226399 297533
rect 231117 297530 231183 297533
rect 208228 297528 226399 297530
rect 208228 297472 226338 297528
rect 226394 297472 226399 297528
rect 208228 297470 226399 297472
rect 208228 297468 208234 297470
rect 226333 297467 226399 297470
rect 229050 297528 231183 297530
rect 229050 297472 231122 297528
rect 231178 297472 231183 297528
rect 229050 297470 231183 297472
rect 199510 297332 199516 297396
rect 199580 297394 199586 297396
rect 229050 297394 229110 297470
rect 231117 297467 231183 297470
rect 199580 297334 229110 297394
rect 230381 297394 230447 297397
rect 254025 297394 254091 297397
rect 230381 297392 254091 297394
rect 230381 297336 230386 297392
rect 230442 297336 254030 297392
rect 254086 297336 254091 297392
rect 230381 297334 254091 297336
rect 199580 297332 199586 297334
rect 230381 297331 230447 297334
rect 254025 297331 254091 297334
rect 158805 297122 158871 297125
rect 156676 297120 158871 297122
rect 156676 297064 158810 297120
rect 158866 297064 158871 297120
rect 156676 297062 158871 297064
rect 158805 297059 158871 297062
rect 226701 296986 226767 296989
rect 269849 296986 269915 296989
rect 226701 296984 269915 296986
rect 226701 296928 226706 296984
rect 226762 296928 269854 296984
rect 269910 296928 269915 296984
rect 226701 296926 269915 296928
rect 226701 296923 226767 296926
rect 269849 296923 269915 296926
rect 207565 296850 207631 296853
rect 278037 296850 278103 296853
rect 207565 296848 278103 296850
rect 207565 296792 207570 296848
rect 207626 296792 278042 296848
rect 278098 296792 278103 296848
rect 207565 296790 278103 296792
rect 207565 296787 207631 296790
rect 278037 296787 278103 296790
rect 206277 296714 206343 296717
rect 214557 296714 214623 296717
rect 206277 296712 214623 296714
rect 206277 296656 206282 296712
rect 206338 296656 214562 296712
rect 214618 296656 214623 296712
rect 206277 296654 214623 296656
rect 206277 296651 206343 296654
rect 214557 296651 214623 296654
rect 67173 296170 67239 296173
rect 67950 296170 67956 296172
rect 67173 296168 67956 296170
rect 67173 296112 67178 296168
rect 67234 296112 67956 296168
rect 67173 296110 67956 296112
rect 67173 296107 67239 296110
rect 67950 296108 67956 296110
rect 68020 296170 68026 296172
rect 68878 296170 68938 296548
rect 68020 296110 68938 296170
rect 68020 296108 68026 296110
rect 158805 296034 158871 296037
rect 156676 296032 158871 296034
rect 156676 295976 158810 296032
rect 158866 295976 158871 296032
rect 156676 295974 158871 295976
rect 158805 295971 158871 295974
rect 214598 295972 214604 296036
rect 214668 296034 214674 296036
rect 248413 296034 248479 296037
rect 214668 296032 248479 296034
rect 214668 295976 248418 296032
rect 248474 295976 248479 296032
rect 214668 295974 248479 295976
rect 214668 295972 214674 295974
rect 248413 295971 248479 295974
rect 67633 295490 67699 295493
rect 67633 295488 68908 295490
rect 67633 295432 67638 295488
rect 67694 295432 68908 295488
rect 67633 295430 68908 295432
rect 67633 295427 67699 295430
rect 192334 295428 192340 295492
rect 192404 295490 192410 295492
rect 204897 295490 204963 295493
rect 192404 295488 204963 295490
rect 192404 295432 204902 295488
rect 204958 295432 204963 295488
rect 192404 295430 204963 295432
rect 192404 295428 192410 295430
rect 204897 295427 204963 295430
rect 220169 295490 220235 295493
rect 220813 295490 220879 295493
rect 276749 295490 276815 295493
rect 220169 295488 276815 295490
rect 220169 295432 220174 295488
rect 220230 295432 220818 295488
rect 220874 295432 276754 295488
rect 276810 295432 276815 295488
rect 220169 295430 276815 295432
rect 220169 295427 220235 295430
rect 220813 295427 220879 295430
rect 276749 295427 276815 295430
rect 186221 295354 186287 295357
rect 278129 295354 278195 295357
rect 186221 295352 278195 295354
rect 186221 295296 186226 295352
rect 186282 295296 278134 295352
rect 278190 295296 278195 295352
rect 186221 295294 278195 295296
rect 186221 295291 186287 295294
rect 278129 295291 278195 295294
rect 158805 294946 158871 294949
rect 156676 294944 158871 294946
rect 156676 294888 158810 294944
rect 158866 294888 158871 294944
rect 156676 294886 158871 294888
rect 158805 294883 158871 294886
rect 160829 294538 160895 294541
rect 245653 294538 245719 294541
rect 160829 294536 245719 294538
rect 160829 294480 160834 294536
rect 160890 294480 245658 294536
rect 245714 294480 245719 294536
rect 160829 294478 245719 294480
rect 160829 294475 160895 294478
rect 245653 294475 245719 294478
rect 66069 294402 66135 294405
rect 66069 294400 68908 294402
rect 66069 294344 66074 294400
rect 66130 294344 68908 294400
rect 66069 294342 68908 294344
rect 66069 294339 66135 294342
rect 225689 294130 225755 294133
rect 226885 294130 226951 294133
rect 255262 294130 255268 294132
rect 225689 294128 255268 294130
rect 225689 294072 225694 294128
rect 225750 294072 226890 294128
rect 226946 294072 255268 294128
rect 225689 294070 255268 294072
rect 225689 294067 225755 294070
rect 226885 294067 226951 294070
rect 255262 294068 255268 294070
rect 255332 294068 255338 294132
rect 175089 293994 175155 293997
rect 287094 293994 287100 293996
rect 175089 293992 287100 293994
rect 175089 293936 175094 293992
rect 175150 293936 287100 293992
rect 175089 293934 287100 293936
rect 175089 293931 175155 293934
rect 287094 293932 287100 293934
rect 287164 293932 287170 293996
rect 158897 293858 158963 293861
rect 156676 293856 158963 293858
rect 156676 293800 158902 293856
rect 158958 293800 158963 293856
rect 156676 293798 158963 293800
rect 158897 293795 158963 293798
rect 215385 293858 215451 293861
rect 303613 293858 303679 293861
rect 215385 293856 303679 293858
rect 215385 293800 215390 293856
rect 215446 293800 303618 293856
rect 303674 293800 303679 293856
rect 215385 293798 303679 293800
rect 215385 293795 215451 293798
rect 303613 293795 303679 293798
rect 66805 293314 66871 293317
rect 66805 293312 68908 293314
rect -960 293178 480 293268
rect 66805 293256 66810 293312
rect 66866 293256 68908 293312
rect 66805 293254 68908 293256
rect 66805 293251 66871 293254
rect 3601 293178 3667 293181
rect -960 293176 3667 293178
rect -960 293120 3606 293176
rect 3662 293120 3667 293176
rect -960 293118 3667 293120
rect -960 293028 480 293118
rect 3601 293115 3667 293118
rect 193121 293178 193187 293181
rect 203609 293178 203675 293181
rect 193121 293176 203675 293178
rect 193121 293120 193126 293176
rect 193182 293120 203614 293176
rect 203670 293120 203675 293176
rect 193121 293118 203675 293120
rect 193121 293115 193187 293118
rect 203609 293115 203675 293118
rect 158805 293042 158871 293045
rect 156676 293040 158871 293042
rect 156676 292984 158810 293040
rect 158866 292984 158871 293040
rect 156676 292982 158871 292984
rect 158805 292979 158871 292982
rect 212349 292770 212415 292773
rect 215385 292770 215451 292773
rect 212349 292768 215451 292770
rect 212349 292712 212354 292768
rect 212410 292712 215390 292768
rect 215446 292712 215451 292768
rect 212349 292710 215451 292712
rect 212349 292707 212415 292710
rect 215385 292707 215451 292710
rect 221181 292770 221247 292773
rect 262857 292770 262923 292773
rect 221181 292768 262923 292770
rect 221181 292712 221186 292768
rect 221242 292712 262862 292768
rect 262918 292712 262923 292768
rect 221181 292710 262923 292712
rect 221181 292707 221247 292710
rect 262857 292707 262923 292710
rect 169150 292572 169156 292636
rect 169220 292634 169226 292636
rect 232773 292634 232839 292637
rect 169220 292632 232839 292634
rect 169220 292576 232778 292632
rect 232834 292576 232839 292632
rect 169220 292574 232839 292576
rect 169220 292572 169226 292574
rect 232773 292571 232839 292574
rect 303613 292634 303679 292637
rect 304257 292634 304323 292637
rect 303613 292632 304323 292634
rect 303613 292576 303618 292632
rect 303674 292576 304262 292632
rect 304318 292576 304323 292632
rect 303613 292574 304323 292576
rect 303613 292571 303679 292574
rect 304257 292571 304323 292574
rect 160921 292498 160987 292501
rect 227897 292498 227963 292501
rect 160921 292496 227963 292498
rect 160921 292440 160926 292496
rect 160982 292440 227902 292496
rect 227958 292440 227963 292496
rect 160921 292438 227963 292440
rect 160921 292435 160987 292438
rect 227897 292435 227963 292438
rect 66805 292226 66871 292229
rect 66805 292224 68908 292226
rect 66805 292168 66810 292224
rect 66866 292168 68908 292224
rect 66805 292166 68908 292168
rect 66805 292163 66871 292166
rect 227897 292090 227963 292093
rect 228449 292090 228515 292093
rect 227897 292088 228515 292090
rect 227897 292032 227902 292088
rect 227958 292032 228454 292088
rect 228510 292032 228515 292088
rect 227897 292030 228515 292032
rect 227897 292027 227963 292030
rect 228449 292027 228515 292030
rect 158805 291954 158871 291957
rect 156676 291952 158871 291954
rect 156676 291896 158810 291952
rect 158866 291896 158871 291952
rect 156676 291894 158871 291896
rect 158805 291891 158871 291894
rect 200389 291954 200455 291957
rect 202873 291954 202939 291957
rect 200389 291952 202939 291954
rect 200389 291896 200394 291952
rect 200450 291896 202878 291952
rect 202934 291896 202939 291952
rect 200389 291894 202939 291896
rect 200389 291891 200455 291894
rect 202873 291891 202939 291894
rect 246798 291756 246804 291820
rect 246868 291818 246874 291820
rect 365713 291818 365779 291821
rect 246868 291816 365779 291818
rect 246868 291760 365718 291816
rect 365774 291760 365779 291816
rect 246868 291758 365779 291760
rect 246868 291756 246874 291758
rect 365713 291755 365779 291758
rect 202137 291410 202203 291413
rect 260925 291410 260991 291413
rect 202137 291408 260991 291410
rect 202137 291352 202142 291408
rect 202198 291352 260930 291408
rect 260986 291352 260991 291408
rect 202137 291350 260991 291352
rect 202137 291347 202203 291350
rect 260925 291347 260991 291350
rect 226977 291274 227043 291277
rect 227621 291274 227687 291277
rect 304993 291274 305059 291277
rect 226977 291272 305059 291274
rect 226977 291216 226982 291272
rect 227038 291216 227626 291272
rect 227682 291216 304998 291272
rect 305054 291216 305059 291272
rect 226977 291214 305059 291216
rect 226977 291211 227043 291214
rect 227621 291211 227687 291214
rect 304993 291211 305059 291214
rect 67081 291138 67147 291141
rect 67449 291138 67515 291141
rect 67081 291136 68908 291138
rect 67081 291080 67086 291136
rect 67142 291080 67454 291136
rect 67510 291080 68908 291136
rect 67081 291078 68908 291080
rect 67081 291075 67147 291078
rect 67449 291075 67515 291078
rect 198590 291076 198596 291140
rect 198660 291138 198666 291140
rect 198660 291078 200130 291138
rect 198660 291076 198666 291078
rect 200070 291002 200130 291078
rect 200614 291076 200620 291140
rect 200684 291138 200690 291140
rect 207749 291138 207815 291141
rect 226701 291138 226767 291141
rect 200684 291136 207815 291138
rect 200684 291080 207754 291136
rect 207810 291080 207815 291136
rect 200684 291078 207815 291080
rect 200684 291076 200690 291078
rect 207749 291075 207815 291078
rect 209730 291136 226767 291138
rect 209730 291080 226706 291136
rect 226762 291080 226767 291136
rect 209730 291078 226767 291080
rect 200481 291002 200547 291005
rect 209730 291002 209790 291078
rect 226701 291075 226767 291078
rect 200070 291000 209790 291002
rect 200070 290944 200486 291000
rect 200542 290944 209790 291000
rect 200070 290942 209790 290944
rect 220077 291002 220143 291005
rect 234521 291002 234587 291005
rect 220077 291000 234587 291002
rect 220077 290944 220082 291000
rect 220138 290944 234526 291000
rect 234582 290944 234587 291000
rect 220077 290942 234587 290944
rect 200481 290939 200547 290942
rect 220077 290939 220143 290942
rect 234521 290939 234587 290942
rect 158805 290866 158871 290869
rect 156676 290864 158871 290866
rect 156676 290808 158810 290864
rect 158866 290808 158871 290864
rect 156676 290806 158871 290808
rect 158805 290803 158871 290806
rect 233693 290458 233759 290461
rect 240225 290458 240291 290461
rect 265709 290458 265775 290461
rect 233693 290456 265775 290458
rect 233693 290400 233698 290456
rect 233754 290400 240230 290456
rect 240286 290400 265714 290456
rect 265770 290400 265775 290456
rect 233693 290398 265775 290400
rect 233693 290395 233759 290398
rect 240225 290395 240291 290398
rect 265709 290395 265775 290398
rect 66345 290050 66411 290053
rect 246297 290052 246363 290053
rect 246246 290050 246252 290052
rect 66345 290048 68908 290050
rect 66345 289992 66350 290048
rect 66406 289992 68908 290048
rect 66345 289990 68908 289992
rect 246170 289990 246252 290050
rect 246316 290050 246363 290052
rect 295517 290050 295583 290053
rect 295885 290050 295951 290053
rect 246316 290048 295951 290050
rect 246358 289992 295522 290048
rect 295578 289992 295890 290048
rect 295946 289992 295951 290048
rect 66345 289987 66411 289990
rect 246246 289988 246252 289990
rect 246316 289990 295951 289992
rect 246316 289988 246363 289990
rect 246297 289987 246363 289988
rect 295517 289987 295583 289990
rect 295885 289987 295951 289990
rect 191046 289852 191052 289916
rect 191116 289914 191122 289916
rect 223021 289914 223087 289917
rect 191116 289912 223087 289914
rect 191116 289856 223026 289912
rect 223082 289856 223087 289912
rect 191116 289854 223087 289856
rect 191116 289852 191122 289854
rect 223021 289851 223087 289854
rect 224166 289852 224172 289916
rect 224236 289914 224242 289916
rect 297449 289914 297515 289917
rect 224236 289912 297515 289914
rect 224236 289856 297454 289912
rect 297510 289856 297515 289912
rect 224236 289854 297515 289856
rect 224236 289852 224242 289854
rect 297449 289851 297515 289854
rect 158897 289778 158963 289781
rect 187049 289780 187115 289781
rect 156676 289776 158963 289778
rect 156676 289720 158902 289776
rect 158958 289720 158963 289776
rect 156676 289718 158963 289720
rect 158897 289715 158963 289718
rect 186998 289716 187004 289780
rect 187068 289778 187115 289780
rect 203149 289778 203215 289781
rect 204253 289778 204319 289781
rect 187068 289776 187160 289778
rect 187110 289720 187160 289776
rect 187068 289718 187160 289720
rect 203149 289776 204319 289778
rect 203149 289720 203154 289776
rect 203210 289720 204258 289776
rect 204314 289720 204319 289776
rect 203149 289718 204319 289720
rect 187068 289716 187115 289718
rect 187049 289715 187115 289716
rect 203149 289715 203215 289718
rect 204253 289715 204319 289718
rect 211981 289778 212047 289781
rect 213177 289778 213243 289781
rect 211981 289776 213243 289778
rect 211981 289720 211986 289776
rect 212042 289720 213182 289776
rect 213238 289720 213243 289776
rect 211981 289718 213243 289720
rect 211981 289715 212047 289718
rect 213177 289715 213243 289718
rect 160870 289172 160876 289236
rect 160940 289234 160946 289236
rect 168966 289234 168972 289236
rect 160940 289174 168972 289234
rect 160940 289172 160946 289174
rect 168966 289172 168972 289174
rect 169036 289172 169042 289236
rect 204253 289234 204319 289237
rect 238518 289234 238524 289236
rect 204253 289232 238524 289234
rect 204253 289176 204258 289232
rect 204314 289176 238524 289232
rect 204253 289174 238524 289176
rect 204253 289171 204319 289174
rect 238518 289172 238524 289174
rect 238588 289172 238594 289236
rect 162761 289098 162827 289101
rect 186814 289098 186820 289100
rect 162761 289096 186820 289098
rect 162761 289040 162766 289096
rect 162822 289040 186820 289096
rect 162761 289038 186820 289040
rect 162761 289035 162827 289038
rect 186814 289036 186820 289038
rect 186884 289036 186890 289100
rect 187049 289098 187115 289101
rect 209957 289098 210023 289101
rect 210601 289098 210667 289101
rect 187049 289096 210667 289098
rect 187049 289040 187054 289096
rect 187110 289040 209962 289096
rect 210018 289040 210606 289096
rect 210662 289040 210667 289096
rect 187049 289038 210667 289040
rect 187049 289035 187115 289038
rect 209957 289035 210023 289038
rect 210601 289035 210667 289038
rect 218053 289098 218119 289101
rect 232497 289098 232563 289101
rect 359457 289098 359523 289101
rect 218053 289096 359523 289098
rect 218053 289040 218058 289096
rect 218114 289040 232502 289096
rect 232558 289040 359462 289096
rect 359518 289040 359523 289096
rect 218053 289038 359523 289040
rect 218053 289035 218119 289038
rect 232497 289035 232563 289038
rect 359457 289035 359523 289038
rect 66805 288962 66871 288965
rect 66805 288960 68908 288962
rect 66805 288904 66810 288960
rect 66866 288904 68908 288960
rect 66805 288902 68908 288904
rect 66805 288899 66871 288902
rect 158805 288690 158871 288693
rect 156676 288688 158871 288690
rect 156676 288632 158810 288688
rect 158866 288632 158871 288688
rect 156676 288630 158871 288632
rect 158805 288627 158871 288630
rect 241421 288690 241487 288693
rect 258901 288690 258967 288693
rect 241421 288688 258967 288690
rect 241421 288632 241426 288688
rect 241482 288632 258906 288688
rect 258962 288632 258967 288688
rect 241421 288630 258967 288632
rect 241421 288627 241487 288630
rect 258901 288627 258967 288630
rect 195145 288554 195211 288557
rect 211981 288554 212047 288557
rect 195145 288552 212047 288554
rect 195145 288496 195150 288552
rect 195206 288496 211986 288552
rect 212042 288496 212047 288552
rect 195145 288494 212047 288496
rect 195145 288491 195211 288494
rect 211981 288491 212047 288494
rect 220169 288554 220235 288557
rect 226926 288554 226932 288556
rect 220169 288552 226932 288554
rect 220169 288496 220174 288552
rect 220230 288496 226932 288552
rect 220169 288494 226932 288496
rect 220169 288491 220235 288494
rect 226926 288492 226932 288494
rect 226996 288492 227002 288556
rect 232773 288554 232839 288557
rect 253841 288554 253907 288557
rect 232773 288552 253907 288554
rect 232773 288496 232778 288552
rect 232834 288496 253846 288552
rect 253902 288496 253907 288552
rect 232773 288494 253907 288496
rect 232773 288491 232839 288494
rect 253841 288491 253907 288494
rect 215293 288418 215359 288421
rect 216029 288418 216095 288421
rect 215293 288416 216095 288418
rect 215293 288360 215298 288416
rect 215354 288360 216034 288416
rect 216090 288360 216095 288416
rect 215293 288358 216095 288360
rect 215293 288355 215359 288358
rect 216029 288355 216095 288358
rect 225597 288418 225663 288421
rect 332593 288418 332659 288421
rect 225597 288416 332659 288418
rect 225597 288360 225602 288416
rect 225658 288360 332598 288416
rect 332654 288360 332659 288416
rect 225597 288358 332659 288360
rect 225597 288355 225663 288358
rect 332593 288355 332659 288358
rect 67357 287874 67423 287877
rect 67357 287872 68908 287874
rect 67357 287816 67362 287872
rect 67418 287816 68908 287872
rect 67357 287814 68908 287816
rect 67357 287811 67423 287814
rect 216673 287738 216739 287741
rect 254117 287738 254183 287741
rect 216673 287736 254183 287738
rect 216673 287680 216678 287736
rect 216734 287680 254122 287736
rect 254178 287680 254183 287736
rect 216673 287678 254183 287680
rect 216673 287675 216739 287678
rect 254117 287675 254183 287678
rect 158805 287602 158871 287605
rect 156676 287600 158871 287602
rect 156676 287544 158810 287600
rect 158866 287544 158871 287600
rect 156676 287542 158871 287544
rect 158805 287539 158871 287542
rect 215293 287602 215359 287605
rect 215293 287600 219450 287602
rect 215293 287544 215298 287600
rect 215354 287544 219450 287600
rect 215293 287542 219450 287544
rect 215293 287539 215359 287542
rect 194501 287466 194567 287469
rect 215201 287466 215267 287469
rect 194501 287464 215267 287466
rect 194501 287408 194506 287464
rect 194562 287408 215206 287464
rect 215262 287408 215267 287464
rect 194501 287406 215267 287408
rect 219390 287466 219450 287542
rect 232078 287466 232084 287468
rect 219390 287406 232084 287466
rect 194501 287403 194567 287406
rect 215201 287403 215267 287406
rect 232078 287404 232084 287406
rect 232148 287404 232154 287468
rect 196617 287330 196683 287333
rect 217317 287330 217383 287333
rect 196617 287328 217383 287330
rect 196617 287272 196622 287328
rect 196678 287272 217322 287328
rect 217378 287272 217383 287328
rect 196617 287270 217383 287272
rect 196617 287267 196683 287270
rect 217317 287267 217383 287270
rect 183461 287194 183527 287197
rect 217685 287194 217751 287197
rect 183461 287192 217751 287194
rect 183461 287136 183466 287192
rect 183522 287136 217690 287192
rect 217746 287136 217751 287192
rect 183461 287134 217751 287136
rect 183461 287131 183527 287134
rect 217685 287131 217751 287134
rect 234245 287194 234311 287197
rect 243077 287194 243143 287197
rect 234245 287192 243143 287194
rect 234245 287136 234250 287192
rect 234306 287136 243082 287192
rect 243138 287136 243143 287192
rect 234245 287134 243143 287136
rect 234245 287131 234311 287134
rect 243077 287131 243143 287134
rect 66253 286786 66319 286789
rect 66253 286784 68908 286786
rect 66253 286728 66258 286784
rect 66314 286728 68908 286784
rect 66253 286726 68908 286728
rect 66253 286723 66319 286726
rect 156646 285970 156706 286484
rect 253197 286378 253263 286381
rect 283782 286378 283788 286380
rect 253197 286376 283788 286378
rect 253197 286320 253202 286376
rect 253258 286320 283788 286376
rect 253197 286318 283788 286320
rect 253197 286315 253263 286318
rect 283782 286316 283788 286318
rect 283852 286316 283858 286380
rect 238109 286106 238175 286109
rect 243077 286106 243143 286109
rect 238109 286104 243143 286106
rect 238109 286048 238114 286104
rect 238170 286048 243082 286104
rect 243138 286048 243143 286104
rect 238109 286046 243143 286048
rect 238109 286043 238175 286046
rect 243077 286043 243143 286046
rect 237281 285970 237347 285973
rect 156646 285968 237347 285970
rect 156646 285912 237286 285968
rect 237342 285912 237347 285968
rect 156646 285910 237347 285912
rect 237281 285907 237347 285910
rect 237649 285970 237715 285973
rect 243670 285970 243676 285972
rect 237649 285968 243676 285970
rect 237649 285912 237654 285968
rect 237710 285912 243676 285968
rect 237649 285910 243676 285912
rect 237649 285907 237715 285910
rect 243670 285908 243676 285910
rect 243740 285908 243746 285972
rect 212390 285772 212396 285836
rect 212460 285834 212466 285836
rect 217225 285834 217291 285837
rect 212460 285832 217291 285834
rect 212460 285776 217230 285832
rect 217286 285776 217291 285832
rect 212460 285774 217291 285776
rect 212460 285772 212466 285774
rect 217225 285771 217291 285774
rect 222837 285834 222903 285837
rect 225965 285834 226031 285837
rect 222837 285832 226031 285834
rect 222837 285776 222842 285832
rect 222898 285776 225970 285832
rect 226026 285776 226031 285832
rect 222837 285774 226031 285776
rect 222837 285771 222903 285774
rect 225965 285771 226031 285774
rect 236637 285834 236703 285837
rect 250529 285834 250595 285837
rect 236637 285832 250595 285834
rect 236637 285776 236642 285832
rect 236698 285776 250534 285832
rect 250590 285776 250595 285832
rect 236637 285774 250595 285776
rect 236637 285771 236703 285774
rect 250529 285771 250595 285774
rect 66805 285698 66871 285701
rect 195145 285698 195211 285701
rect 66805 285696 68908 285698
rect 66805 285640 66810 285696
rect 66866 285640 68908 285696
rect 66805 285638 68908 285640
rect 195145 285696 202890 285698
rect 195145 285640 195150 285696
rect 195206 285640 202890 285696
rect 195145 285638 202890 285640
rect 66805 285635 66871 285638
rect 195145 285635 195211 285638
rect 202830 285562 202890 285638
rect 204478 285636 204484 285700
rect 204548 285698 204554 285700
rect 205173 285698 205239 285701
rect 204548 285696 205239 285698
rect 204548 285640 205178 285696
rect 205234 285640 205239 285696
rect 204548 285638 205239 285640
rect 204548 285636 204554 285638
rect 205173 285635 205239 285638
rect 215937 285698 216003 285701
rect 218646 285698 218652 285700
rect 215937 285696 218652 285698
rect 215937 285640 215942 285696
rect 215998 285640 218652 285696
rect 215937 285638 218652 285640
rect 215937 285635 216003 285638
rect 218646 285636 218652 285638
rect 218716 285636 218722 285700
rect 223941 285698 224007 285701
rect 224166 285698 224172 285700
rect 223941 285696 224172 285698
rect 223941 285640 223946 285696
rect 224002 285640 224172 285696
rect 223941 285638 224172 285640
rect 223941 285635 224007 285638
rect 224166 285636 224172 285638
rect 224236 285636 224242 285700
rect 225045 285698 225111 285701
rect 228214 285698 228220 285700
rect 225045 285696 228220 285698
rect 225045 285640 225050 285696
rect 225106 285640 228220 285696
rect 225045 285638 228220 285640
rect 225045 285635 225111 285638
rect 228214 285636 228220 285638
rect 228284 285636 228290 285700
rect 235993 285698 236059 285701
rect 236494 285698 236500 285700
rect 235993 285696 236500 285698
rect 235993 285640 235998 285696
rect 236054 285640 236500 285696
rect 235993 285638 236500 285640
rect 235993 285635 236059 285638
rect 236494 285636 236500 285638
rect 236564 285636 236570 285700
rect 242893 285698 242959 285701
rect 243537 285698 243603 285701
rect 338757 285698 338823 285701
rect 242893 285696 338823 285698
rect 242893 285640 242898 285696
rect 242954 285640 243542 285696
rect 243598 285640 338762 285696
rect 338818 285640 338823 285696
rect 242893 285638 338823 285640
rect 242893 285635 242959 285638
rect 243537 285635 243603 285638
rect 338757 285635 338823 285638
rect 237649 285562 237715 285565
rect 202830 285560 237715 285562
rect 202830 285504 237654 285560
rect 237710 285504 237715 285560
rect 202830 285502 237715 285504
rect 237649 285499 237715 285502
rect 158805 285426 158871 285429
rect 156676 285424 158871 285426
rect 156676 285368 158810 285424
rect 158866 285368 158871 285424
rect 156676 285366 158871 285368
rect 158805 285363 158871 285366
rect 583520 285276 584960 285516
rect 188521 285154 188587 285157
rect 247677 285156 247743 285157
rect 192334 285154 192340 285156
rect 188521 285152 192340 285154
rect 188521 285096 188526 285152
rect 188582 285096 192340 285152
rect 188521 285094 192340 285096
rect 188521 285091 188587 285094
rect 192334 285092 192340 285094
rect 192404 285092 192410 285156
rect 247677 285152 247724 285156
rect 247788 285154 247794 285156
rect 247677 285096 247682 285152
rect 247677 285092 247724 285096
rect 247788 285094 247834 285154
rect 247788 285092 247794 285094
rect 247677 285091 247743 285092
rect 181437 285018 181503 285021
rect 204253 285018 204319 285021
rect 181437 285016 204319 285018
rect 181437 284960 181442 285016
rect 181498 284960 204258 285016
rect 204314 284960 204319 285016
rect 181437 284958 204319 284960
rect 181437 284955 181503 284958
rect 204253 284955 204319 284958
rect 237373 285018 237439 285021
rect 253289 285018 253355 285021
rect 237373 285016 253355 285018
rect 237373 284960 237378 285016
rect 237434 284960 253294 285016
rect 253350 284960 253355 285016
rect 237373 284958 253355 284960
rect 237373 284955 237439 284958
rect 253289 284955 253355 284958
rect 158805 284882 158871 284885
rect 202137 284882 202203 284885
rect 158805 284880 202203 284882
rect 158805 284824 158810 284880
rect 158866 284824 202142 284880
rect 202198 284824 202203 284880
rect 158805 284822 202203 284824
rect 158805 284819 158871 284822
rect 202137 284819 202203 284822
rect 204897 284882 204963 284885
rect 243813 284882 243879 284885
rect 204897 284880 243879 284882
rect 204897 284824 204902 284880
rect 204958 284824 243818 284880
rect 243874 284824 243879 284880
rect 204897 284822 243879 284824
rect 204897 284819 204963 284822
rect 243813 284819 243879 284822
rect 66662 284548 66668 284612
rect 66732 284610 66738 284612
rect 66805 284610 66871 284613
rect 66732 284608 68908 284610
rect 66732 284552 66810 284608
rect 66866 284552 68908 284608
rect 66732 284550 68908 284552
rect 66732 284548 66738 284550
rect 66805 284547 66871 284550
rect 218513 284474 218579 284477
rect 244590 284474 244596 284476
rect 218513 284472 244596 284474
rect 218513 284416 218518 284472
rect 218574 284416 244596 284472
rect 218513 284414 244596 284416
rect 218513 284411 218579 284414
rect 244590 284412 244596 284414
rect 244660 284412 244666 284476
rect 160093 284338 160159 284341
rect 156676 284336 160159 284338
rect 156676 284280 160098 284336
rect 160154 284280 160159 284336
rect 156676 284278 160159 284280
rect 160093 284275 160159 284278
rect 198774 284276 198780 284340
rect 198844 284338 198850 284340
rect 206093 284338 206159 284341
rect 198844 284336 206159 284338
rect 198844 284280 206098 284336
rect 206154 284280 206159 284336
rect 198844 284278 206159 284280
rect 198844 284276 198850 284278
rect 206093 284275 206159 284278
rect 243813 284338 243879 284341
rect 332593 284338 332659 284341
rect 243813 284336 332659 284338
rect 243813 284280 243818 284336
rect 243874 284280 332598 284336
rect 332654 284280 332659 284336
rect 243813 284278 332659 284280
rect 243813 284275 243879 284278
rect 332593 284275 332659 284278
rect 243077 284202 243143 284205
rect 268377 284202 268443 284205
rect 243077 284200 268443 284202
rect 243077 284144 243082 284200
rect 243138 284144 268382 284200
rect 268438 284144 268443 284200
rect 243077 284142 268443 284144
rect 243077 284139 243143 284142
rect 268377 284139 268443 284142
rect 192702 284004 192708 284068
rect 192772 284066 192778 284068
rect 200481 284066 200547 284069
rect 192772 284064 200547 284066
rect 192772 284008 200486 284064
rect 200542 284008 200547 284064
rect 192772 284006 200547 284008
rect 192772 284004 192778 284006
rect 200481 284003 200547 284006
rect 242985 284066 243051 284069
rect 280286 284066 280292 284068
rect 242985 284064 280292 284066
rect 242985 284008 242990 284064
rect 243046 284008 280292 284064
rect 242985 284006 280292 284008
rect 242985 284003 243051 284006
rect 280286 284004 280292 284006
rect 280356 284004 280362 284068
rect 205357 283932 205423 283933
rect 214465 283932 214531 283933
rect 216121 283932 216187 283933
rect 205357 283930 205404 283932
rect 205312 283928 205404 283930
rect 205312 283872 205362 283928
rect 205312 283870 205404 283872
rect 205357 283868 205404 283870
rect 205468 283868 205474 283932
rect 214414 283930 214420 283932
rect 214374 283870 214420 283930
rect 214484 283928 214531 283932
rect 216070 283930 216076 283932
rect 214526 283872 214531 283928
rect 214414 283868 214420 283870
rect 214484 283868 214531 283872
rect 216030 283870 216076 283930
rect 216140 283928 216187 283932
rect 216182 283872 216187 283928
rect 216070 283868 216076 283870
rect 216140 283868 216187 283872
rect 205357 283867 205423 283868
rect 214465 283867 214531 283868
rect 216121 283867 216187 283868
rect 220261 283930 220327 283933
rect 222326 283930 222332 283932
rect 220261 283928 222332 283930
rect 220261 283872 220266 283928
rect 220322 283872 222332 283928
rect 220261 283870 222332 283872
rect 220261 283867 220327 283870
rect 222326 283868 222332 283870
rect 222396 283868 222402 283932
rect 223757 283930 223823 283933
rect 226006 283930 226012 283932
rect 223757 283928 226012 283930
rect 223757 283872 223762 283928
rect 223818 283872 226012 283928
rect 223757 283870 226012 283872
rect 223757 283867 223823 283870
rect 226006 283868 226012 283870
rect 226076 283868 226082 283932
rect 229461 283930 229527 283933
rect 229686 283930 229692 283932
rect 229461 283928 229692 283930
rect 229461 283872 229466 283928
rect 229522 283872 229692 283928
rect 229461 283870 229692 283872
rect 229461 283867 229527 283870
rect 229686 283868 229692 283870
rect 229756 283868 229762 283932
rect 230933 283930 230999 283933
rect 231894 283930 231900 283932
rect 230933 283928 231900 283930
rect 230933 283872 230938 283928
rect 230994 283872 231900 283928
rect 230933 283870 231900 283872
rect 230933 283867 230999 283870
rect 231894 283868 231900 283870
rect 231964 283868 231970 283932
rect 236494 283868 236500 283932
rect 236564 283930 236570 283932
rect 236729 283930 236795 283933
rect 236564 283928 236795 283930
rect 236564 283872 236734 283928
rect 236790 283872 236795 283928
rect 236564 283870 236795 283872
rect 236564 283868 236570 283870
rect 236729 283867 236795 283870
rect 246941 283794 247007 283797
rect 244076 283792 247007 283794
rect 66805 283522 66871 283525
rect 200113 283524 200179 283525
rect 66805 283520 68908 283522
rect 66805 283464 66810 283520
rect 66866 283464 68908 283520
rect 66805 283462 68908 283464
rect 66805 283459 66871 283462
rect 200062 283460 200068 283524
rect 200132 283522 200179 283524
rect 200132 283520 200224 283522
rect 200174 283464 200224 283520
rect 200132 283462 200224 283464
rect 200132 283460 200179 283462
rect 200113 283459 200179 283460
rect 184841 283250 184907 283253
rect 200438 283250 200498 283764
rect 244076 283736 246946 283792
rect 247002 283736 247007 283792
rect 244076 283734 247007 283736
rect 246941 283731 247007 283734
rect 244590 283596 244596 283660
rect 244660 283658 244666 283660
rect 257521 283658 257587 283661
rect 244660 283656 257587 283658
rect 244660 283600 257526 283656
rect 257582 283600 257587 283656
rect 244660 283598 257587 283600
rect 244660 283596 244666 283598
rect 257521 283595 257587 283598
rect 297449 283522 297515 283525
rect 334801 283522 334867 283525
rect 297449 283520 334867 283522
rect 297449 283464 297454 283520
rect 297510 283464 334806 283520
rect 334862 283464 334867 283520
rect 297449 283462 334867 283464
rect 297449 283459 297515 283462
rect 334801 283459 334867 283462
rect 246297 283250 246363 283253
rect 184841 283248 200498 283250
rect 156646 282978 156706 283220
rect 184841 283192 184846 283248
rect 184902 283192 200498 283248
rect 184841 283190 200498 283192
rect 244076 283248 246363 283250
rect 244076 283192 246302 283248
rect 246358 283192 246363 283248
rect 244076 283190 246363 283192
rect 184841 283187 184907 283190
rect 246297 283187 246363 283190
rect 183001 283114 183067 283117
rect 184381 283114 184447 283117
rect 183001 283112 184447 283114
rect 183001 283056 183006 283112
rect 183062 283056 184386 283112
rect 184442 283056 184447 283112
rect 183001 283054 184447 283056
rect 183001 283051 183067 283054
rect 184381 283051 184447 283054
rect 183277 282978 183343 282981
rect 156646 282976 183343 282978
rect 156646 282920 183282 282976
rect 183338 282920 183343 282976
rect 156646 282918 183343 282920
rect 183277 282915 183343 282918
rect 198590 282916 198596 282980
rect 198660 282978 198666 282980
rect 198660 282918 200284 282978
rect 198660 282916 198666 282918
rect 188337 282842 188403 282845
rect 191782 282842 191788 282844
rect 188337 282840 191788 282842
rect 188337 282784 188342 282840
rect 188398 282784 191788 282840
rect 188337 282782 191788 282784
rect 188337 282779 188403 282782
rect 191782 282780 191788 282782
rect 191852 282842 191858 282844
rect 192702 282842 192708 282844
rect 191852 282782 192708 282842
rect 191852 282780 191858 282782
rect 192702 282780 192708 282782
rect 192772 282780 192778 282844
rect 251081 282842 251147 282845
rect 263593 282842 263659 282845
rect 251081 282840 263659 282842
rect 251081 282784 251086 282840
rect 251142 282784 263598 282840
rect 263654 282784 263659 282840
rect 251081 282782 263659 282784
rect 251081 282779 251147 282782
rect 263593 282779 263659 282782
rect 67725 282434 67791 282437
rect 197353 282434 197419 282437
rect 247217 282434 247283 282437
rect 67725 282432 68908 282434
rect 67725 282376 67730 282432
rect 67786 282376 68908 282432
rect 67725 282374 68908 282376
rect 197353 282432 200284 282434
rect 197353 282376 197358 282432
rect 197414 282376 200284 282432
rect 197353 282374 200284 282376
rect 244076 282432 247283 282434
rect 244076 282376 247222 282432
rect 247278 282376 247283 282432
rect 244076 282374 247283 282376
rect 67725 282371 67791 282374
rect 197353 282371 197419 282374
rect 247217 282371 247283 282374
rect 158805 282162 158871 282165
rect 185577 282162 185643 282165
rect 156676 282160 158871 282162
rect 156676 282104 158810 282160
rect 158866 282104 158871 282160
rect 156676 282102 158871 282104
rect 158805 282099 158871 282102
rect 161430 282160 185643 282162
rect 161430 282104 185582 282160
rect 185638 282104 185643 282160
rect 161430 282102 185643 282104
rect 158478 281964 158484 282028
rect 158548 282026 158554 282028
rect 161430 282026 161490 282102
rect 185577 282099 185643 282102
rect 253841 282162 253907 282165
rect 366357 282162 366423 282165
rect 253841 282160 366423 282162
rect 253841 282104 253846 282160
rect 253902 282104 366362 282160
rect 366418 282104 366423 282160
rect 253841 282102 366423 282104
rect 253841 282099 253907 282102
rect 366357 282099 366423 282102
rect 158548 281966 161490 282026
rect 158548 281964 158554 281966
rect 195830 281556 195836 281620
rect 195900 281618 195906 281620
rect 198774 281618 198780 281620
rect 195900 281558 198780 281618
rect 195900 281556 195906 281558
rect 198774 281556 198780 281558
rect 198844 281556 198850 281620
rect 199510 281556 199516 281620
rect 199580 281618 199586 281620
rect 245929 281618 245995 281621
rect 199580 281558 200284 281618
rect 244076 281616 245995 281618
rect 244076 281560 245934 281616
rect 245990 281560 245995 281616
rect 244076 281558 245995 281560
rect 199580 281556 199586 281558
rect 245929 281555 245995 281558
rect 67357 281346 67423 281349
rect 67357 281344 68908 281346
rect 67357 281288 67362 281344
rect 67418 281288 68908 281344
rect 67357 281286 68908 281288
rect 67357 281283 67423 281286
rect 199326 281284 199332 281348
rect 199396 281346 199402 281348
rect 200614 281346 200620 281348
rect 199396 281286 200620 281346
rect 199396 281284 199402 281286
rect 200614 281284 200620 281286
rect 200684 281284 200690 281348
rect 243486 281284 243492 281348
rect 243556 281284 243562 281348
rect 158805 281074 158871 281077
rect 156676 281072 158871 281074
rect 156676 281016 158810 281072
rect 158866 281016 158871 281072
rect 243494 281074 243554 281284
rect 246113 281074 246179 281077
rect 243494 281072 246179 281074
rect 243494 281044 246118 281072
rect 156676 281014 158871 281016
rect 243524 281016 246118 281044
rect 246174 281016 246179 281072
rect 243524 281014 246179 281016
rect 158805 281011 158871 281014
rect 246113 281011 246179 281014
rect 69422 280740 69428 280804
rect 69492 280740 69498 280804
rect 197353 280802 197419 280805
rect 308397 280802 308463 280805
rect 370497 280802 370563 280805
rect 197353 280800 200284 280802
rect 197353 280744 197358 280800
rect 197414 280744 200284 280800
rect 197353 280742 200284 280744
rect 308397 280800 370563 280802
rect 308397 280744 308402 280800
rect 308458 280744 370502 280800
rect 370558 280744 370563 280800
rect 308397 280742 370563 280744
rect 67541 280258 67607 280261
rect 69430 280258 69490 280740
rect 197353 280739 197419 280742
rect 308397 280739 308463 280742
rect 370497 280739 370563 280742
rect 67541 280256 69490 280258
rect -960 279972 480 280212
rect 67541 280200 67546 280256
rect 67602 280228 69490 280256
rect 197445 280258 197511 280261
rect 246246 280258 246252 280260
rect 197445 280256 200284 280258
rect 67602 280200 69460 280228
rect 67541 280198 69460 280200
rect 197445 280200 197450 280256
rect 197506 280200 200284 280256
rect 197445 280198 200284 280200
rect 244076 280198 246252 280258
rect 67541 280195 67607 280198
rect 197445 280195 197511 280198
rect 246246 280196 246252 280198
rect 246316 280196 246322 280260
rect 167637 280122 167703 280125
rect 156646 280120 167703 280122
rect 156646 280064 167642 280120
rect 167698 280064 167703 280120
rect 156646 280062 167703 280064
rect 156646 279956 156706 280062
rect 167637 280059 167703 280062
rect 243997 279986 244063 279989
rect 243862 279984 244063 279986
rect 243862 279928 244002 279984
rect 244058 279928 244063 279984
rect 243862 279926 244063 279928
rect 197353 279442 197419 279445
rect 243862 279442 243922 279926
rect 243997 279923 244063 279926
rect 245929 279442 245995 279445
rect 197353 279440 200284 279442
rect 197353 279384 197358 279440
rect 197414 279384 200284 279440
rect 243862 279440 245995 279442
rect 243862 279412 245934 279440
rect 197353 279382 200284 279384
rect 243892 279384 245934 279412
rect 245990 279384 245995 279440
rect 243892 279382 245995 279384
rect 197353 279379 197419 279382
rect 245929 279379 245995 279382
rect 66621 279170 66687 279173
rect 66621 279168 68908 279170
rect 66621 279112 66626 279168
rect 66682 279112 68908 279168
rect 66621 279110 68908 279112
rect 66621 279107 66687 279110
rect 159817 278898 159883 278901
rect 245929 278898 245995 278901
rect 156676 278896 159883 278898
rect 156676 278840 159822 278896
rect 159878 278840 159883 278896
rect 156676 278838 159883 278840
rect 244076 278896 245995 278898
rect 244076 278840 245934 278896
rect 245990 278840 245995 278896
rect 244076 278838 245995 278840
rect 159817 278835 159883 278838
rect 245929 278835 245995 278838
rect 197445 278626 197511 278629
rect 197445 278624 200284 278626
rect 197445 278568 197450 278624
rect 197506 278568 200284 278624
rect 197445 278566 200284 278568
rect 197445 278563 197511 278566
rect 169569 278218 169635 278221
rect 198733 278218 198799 278221
rect 169569 278216 198799 278218
rect 169569 278160 169574 278216
rect 169630 278160 198738 278216
rect 198794 278160 198799 278216
rect 169569 278158 198799 278160
rect 169569 278155 169635 278158
rect 198733 278155 198799 278158
rect 66805 278082 66871 278085
rect 66805 278080 68908 278082
rect 66805 278024 66810 278080
rect 66866 278024 68908 278080
rect 66805 278022 68908 278024
rect 66805 278019 66871 278022
rect 156454 278020 156460 278084
rect 156524 278082 156530 278084
rect 187049 278082 187115 278085
rect 156524 278080 187115 278082
rect 156524 278024 187054 278080
rect 187110 278024 187115 278080
rect 156524 278022 187115 278024
rect 156524 278020 156530 278022
rect 187049 278019 187115 278022
rect 198365 278082 198431 278085
rect 244365 278082 244431 278085
rect 198365 278080 200284 278082
rect 198365 278024 198370 278080
rect 198426 278024 200284 278080
rect 198365 278022 200284 278024
rect 244076 278080 244431 278082
rect 244076 278024 244370 278080
rect 244426 278024 244431 278080
rect 244076 278022 244431 278024
rect 198365 278019 198431 278022
rect 244365 278019 244431 278022
rect 158621 277810 158687 277813
rect 156676 277808 158687 277810
rect 156676 277752 158626 277808
rect 158682 277752 158687 277808
rect 156676 277750 158687 277752
rect 158621 277747 158687 277750
rect 245929 277538 245995 277541
rect 244076 277536 245995 277538
rect 244076 277480 245934 277536
rect 245990 277480 245995 277536
rect 244076 277478 245995 277480
rect 245929 277475 245995 277478
rect 257337 277538 257403 277541
rect 323669 277538 323735 277541
rect 257337 277536 323735 277538
rect 257337 277480 257342 277536
rect 257398 277480 323674 277536
rect 323730 277480 323735 277536
rect 257337 277478 323735 277480
rect 257337 277475 257403 277478
rect 323669 277475 323735 277478
rect 196934 277340 196940 277404
rect 197004 277402 197010 277404
rect 200062 277402 200068 277404
rect 197004 277342 200068 277402
rect 197004 277340 197010 277342
rect 200062 277340 200068 277342
rect 200132 277340 200138 277404
rect 66805 277266 66871 277269
rect 66805 277264 68908 277266
rect 66805 277208 66810 277264
rect 66866 277208 68908 277264
rect 66805 277206 68908 277208
rect 66805 277203 66871 277206
rect 200254 276994 200314 277236
rect 180750 276934 200314 276994
rect 158805 276722 158871 276725
rect 156676 276720 158871 276722
rect 156676 276664 158810 276720
rect 158866 276664 158871 276720
rect 156676 276662 158871 276664
rect 158805 276659 158871 276662
rect 66253 276178 66319 276181
rect 173709 276178 173775 276181
rect 180750 276178 180810 276934
rect 197445 276722 197511 276725
rect 245745 276722 245811 276725
rect 197445 276720 200284 276722
rect 197445 276664 197450 276720
rect 197506 276664 200284 276720
rect 197445 276662 200284 276664
rect 244076 276720 245811 276722
rect 244076 276664 245750 276720
rect 245806 276664 245811 276720
rect 244076 276662 245811 276664
rect 197445 276659 197511 276662
rect 245745 276659 245811 276662
rect 66253 276176 68908 276178
rect 66253 276120 66258 276176
rect 66314 276120 68908 276176
rect 66253 276118 68908 276120
rect 173709 276176 180810 276178
rect 173709 276120 173714 276176
rect 173770 276120 180810 276176
rect 173709 276118 180810 276120
rect 66253 276115 66319 276118
rect 173709 276115 173775 276118
rect 197537 275906 197603 275909
rect 245929 275906 245995 275909
rect 197537 275904 200284 275906
rect 197537 275848 197542 275904
rect 197598 275848 200284 275904
rect 197537 275846 200284 275848
rect 244076 275904 245995 275906
rect 244076 275848 245934 275904
rect 245990 275848 245995 275904
rect 244076 275846 245995 275848
rect 197537 275843 197603 275846
rect 245929 275843 245995 275846
rect 252502 275708 252508 275772
rect 252572 275770 252578 275772
rect 252829 275770 252895 275773
rect 252572 275768 252895 275770
rect 252572 275712 252834 275768
rect 252890 275712 252895 275768
rect 252572 275710 252895 275712
rect 252572 275708 252578 275710
rect 252829 275707 252895 275710
rect 158805 275634 158871 275637
rect 156676 275632 158871 275634
rect 156676 275576 158810 275632
rect 158866 275576 158871 275632
rect 156676 275574 158871 275576
rect 158805 275571 158871 275574
rect 245929 275362 245995 275365
rect 244076 275360 245995 275362
rect 244076 275304 245934 275360
rect 245990 275304 245995 275360
rect 244076 275302 245995 275304
rect 245929 275299 245995 275302
rect 68878 274682 68938 275060
rect 200070 275030 200284 275090
rect 159541 274954 159607 274957
rect 200070 274954 200130 275030
rect 159541 274952 200130 274954
rect 159541 274896 159546 274952
rect 159602 274896 200130 274952
rect 159541 274894 200130 274896
rect 159541 274891 159607 274894
rect 66118 274622 68938 274682
rect 65885 274546 65951 274549
rect 66118 274546 66178 274622
rect 158805 274546 158871 274549
rect 65885 274544 66178 274546
rect 65885 274488 65890 274544
rect 65946 274488 66178 274544
rect 65885 274486 66178 274488
rect 156676 274544 158871 274546
rect 156676 274488 158810 274544
rect 158866 274488 158871 274544
rect 156676 274486 158871 274488
rect 65885 274483 65951 274486
rect 158805 274483 158871 274486
rect 197445 274546 197511 274549
rect 245837 274546 245903 274549
rect 197445 274544 200284 274546
rect 197445 274488 197450 274544
rect 197506 274488 200284 274544
rect 197445 274486 200284 274488
rect 244076 274544 245903 274546
rect 244076 274488 245842 274544
rect 245898 274488 245903 274544
rect 244076 274486 245903 274488
rect 197445 274483 197511 274486
rect 245837 274483 245903 274486
rect 65885 274140 65951 274141
rect 65885 274138 65932 274140
rect 65840 274136 65932 274138
rect 65840 274080 65890 274136
rect 65840 274078 65932 274080
rect 65885 274076 65932 274078
rect 65996 274076 66002 274140
rect 65885 274075 65951 274076
rect 66989 274002 67055 274005
rect 66989 274000 68908 274002
rect 66989 273944 66994 274000
rect 67050 273944 68908 274000
rect 66989 273942 68908 273944
rect 66989 273939 67055 273942
rect 158805 273458 158871 273461
rect 156676 273456 158871 273458
rect 156676 273400 158810 273456
rect 158866 273400 158871 273456
rect 156676 273398 158871 273400
rect 158805 273395 158871 273398
rect 181621 273458 181687 273461
rect 184289 273458 184355 273461
rect 181621 273456 184355 273458
rect 181621 273400 181626 273456
rect 181682 273400 184294 273456
rect 184350 273400 184355 273456
rect 181621 273398 184355 273400
rect 181621 273395 181687 273398
rect 184289 273395 184355 273398
rect 178861 273322 178927 273325
rect 200254 273322 200314 273700
rect 244046 273458 244106 273700
rect 244917 273458 244983 273461
rect 244046 273456 244983 273458
rect 244046 273400 244922 273456
rect 244978 273400 244983 273456
rect 244046 273398 244983 273400
rect 244917 273395 244983 273398
rect 178861 273320 200314 273322
rect 178861 273264 178866 273320
rect 178922 273264 200314 273320
rect 178861 273262 200314 273264
rect 178861 273259 178927 273262
rect 245837 273186 245903 273189
rect 244076 273184 245903 273186
rect 244076 273128 245842 273184
rect 245898 273128 245903 273184
rect 244076 273126 245903 273128
rect 245837 273123 245903 273126
rect 248454 273124 248460 273188
rect 248524 273186 248530 273188
rect 248597 273186 248663 273189
rect 248524 273184 248663 273186
rect 248524 273128 248602 273184
rect 248658 273128 248663 273184
rect 248524 273126 248663 273128
rect 248524 273124 248530 273126
rect 248597 273123 248663 273126
rect 251265 273052 251331 273053
rect 251214 273050 251220 273052
rect 251174 272990 251220 273050
rect 251284 273048 251331 273052
rect 251326 272992 251331 273048
rect 251214 272988 251220 272990
rect 251284 272988 251331 272992
rect 251265 272987 251331 272988
rect 66253 272914 66319 272917
rect 197445 272914 197511 272917
rect 66253 272912 68908 272914
rect 66253 272856 66258 272912
rect 66314 272856 68908 272912
rect 66253 272854 68908 272856
rect 197445 272912 200284 272914
rect 197445 272856 197450 272912
rect 197506 272856 200284 272912
rect 197445 272854 200284 272856
rect 66253 272851 66319 272854
rect 197445 272851 197511 272854
rect 181294 272506 181300 272508
rect 171090 272446 181300 272506
rect 156646 271962 156706 272340
rect 169518 271962 169524 271964
rect 156646 271902 169524 271962
rect 169518 271900 169524 271902
rect 169588 271962 169594 271964
rect 171090 271962 171150 272446
rect 181294 272444 181300 272446
rect 181364 272444 181370 272508
rect 199469 272370 199535 272373
rect 245929 272370 245995 272373
rect 199469 272368 200284 272370
rect 199469 272312 199474 272368
rect 199530 272312 200284 272368
rect 199469 272310 200284 272312
rect 244076 272368 245995 272370
rect 244076 272312 245934 272368
rect 245990 272312 245995 272368
rect 244076 272310 245995 272312
rect 199469 272307 199535 272310
rect 245929 272307 245995 272310
rect 582741 272234 582807 272237
rect 583520 272234 584960 272324
rect 582741 272232 584960 272234
rect 582741 272176 582746 272232
rect 582802 272176 584960 272232
rect 582741 272174 584960 272176
rect 582741 272171 582807 272174
rect 583520 272084 584960 272174
rect 169588 271902 171150 271962
rect 169588 271900 169594 271902
rect 66110 271764 66116 271828
rect 66180 271826 66186 271828
rect 66180 271766 68908 271826
rect 66180 271764 66186 271766
rect 197445 271554 197511 271557
rect 245929 271554 245995 271557
rect 197445 271552 200284 271554
rect 197445 271496 197450 271552
rect 197506 271496 200284 271552
rect 197445 271494 200284 271496
rect 244076 271552 245995 271554
rect 244076 271496 245934 271552
rect 245990 271496 245995 271552
rect 244076 271494 245995 271496
rect 197445 271491 197511 271494
rect 245929 271491 245995 271494
rect 158805 271282 158871 271285
rect 156676 271280 158871 271282
rect 156676 271224 158810 271280
rect 158866 271224 158871 271280
rect 156676 271222 158871 271224
rect 158805 271219 158871 271222
rect 174721 271146 174787 271149
rect 191046 271146 191052 271148
rect 174721 271144 191052 271146
rect 174721 271088 174726 271144
rect 174782 271088 191052 271144
rect 174721 271086 191052 271088
rect 174721 271083 174787 271086
rect 191046 271084 191052 271086
rect 191116 271084 191122 271148
rect 198406 270948 198412 271012
rect 198476 271010 198482 271012
rect 245837 271010 245903 271013
rect 198476 270950 200284 271010
rect 244076 271008 245903 271010
rect 244076 270952 245842 271008
rect 245898 270952 245903 271008
rect 244076 270950 245903 270952
rect 198476 270948 198482 270950
rect 245837 270947 245903 270950
rect 66897 270738 66963 270741
rect 66897 270736 68908 270738
rect 66897 270680 66902 270736
rect 66958 270680 68908 270736
rect 66897 270678 68908 270680
rect 66897 270675 66963 270678
rect 250294 270404 250300 270468
rect 250364 270466 250370 270468
rect 251265 270466 251331 270469
rect 250364 270464 251331 270466
rect 250364 270408 251270 270464
rect 251326 270408 251331 270464
rect 250364 270406 251331 270408
rect 250364 270404 250370 270406
rect 251265 270403 251331 270406
rect 159950 270194 159956 270196
rect 156676 270134 159956 270194
rect 159950 270132 159956 270134
rect 160020 270194 160026 270196
rect 163446 270194 163452 270196
rect 160020 270134 163452 270194
rect 160020 270132 160026 270134
rect 163446 270132 163452 270134
rect 163516 270132 163522 270196
rect 197445 270194 197511 270197
rect 245929 270194 245995 270197
rect 197445 270192 200284 270194
rect 197445 270136 197450 270192
rect 197506 270136 200284 270192
rect 197445 270134 200284 270136
rect 244076 270192 245995 270194
rect 244076 270136 245934 270192
rect 245990 270136 245995 270192
rect 244076 270134 245995 270136
rect 197445 270131 197511 270134
rect 245929 270131 245995 270134
rect 67766 269588 67772 269652
rect 67836 269650 67842 269652
rect 244273 269650 244339 269653
rect 246297 269650 246363 269653
rect 67836 269590 68908 269650
rect 244076 269648 246363 269650
rect 244076 269592 244278 269648
rect 244334 269592 246302 269648
rect 246358 269592 246363 269648
rect 244076 269590 246363 269592
rect 67836 269588 67842 269590
rect 244273 269587 244339 269590
rect 246297 269587 246363 269590
rect 200070 269318 200284 269378
rect 169661 269242 169727 269245
rect 170397 269242 170463 269245
rect 200070 269242 200130 269318
rect 169661 269240 200130 269242
rect 169661 269184 169666 269240
rect 169722 269184 170402 269240
rect 170458 269184 200130 269240
rect 169661 269182 200130 269184
rect 253289 269242 253355 269245
rect 260046 269242 260052 269244
rect 253289 269240 260052 269242
rect 253289 269184 253294 269240
rect 253350 269184 260052 269240
rect 253289 269182 260052 269184
rect 169661 269179 169727 269182
rect 170397 269179 170463 269182
rect 253289 269179 253355 269182
rect 260046 269180 260052 269182
rect 260116 269180 260122 269244
rect 158805 269106 158871 269109
rect 156676 269104 158871 269106
rect 156676 269048 158810 269104
rect 158866 269048 158871 269104
rect 156676 269046 158871 269048
rect 158805 269043 158871 269046
rect 197537 268834 197603 268837
rect 244457 268834 244523 268837
rect 197537 268832 200284 268834
rect 197537 268776 197542 268832
rect 197598 268776 200284 268832
rect 197537 268774 200284 268776
rect 244076 268832 244523 268834
rect 244076 268776 244462 268832
rect 244518 268776 244523 268832
rect 244076 268774 244523 268776
rect 197537 268771 197603 268774
rect 244457 268771 244523 268774
rect 66805 268562 66871 268565
rect 187141 268562 187207 268565
rect 196750 268562 196756 268564
rect 66805 268560 68908 268562
rect 66805 268504 66810 268560
rect 66866 268504 68908 268560
rect 66805 268502 68908 268504
rect 187141 268560 196756 268562
rect 187141 268504 187146 268560
rect 187202 268504 196756 268560
rect 187141 268502 196756 268504
rect 66805 268499 66871 268502
rect 187141 268499 187207 268502
rect 196750 268500 196756 268502
rect 196820 268500 196826 268564
rect 171961 268426 172027 268429
rect 196566 268426 196572 268428
rect 171961 268424 196572 268426
rect 171961 268368 171966 268424
rect 172022 268368 196572 268424
rect 171961 268366 196572 268368
rect 171961 268363 172027 268366
rect 196566 268364 196572 268366
rect 196636 268364 196642 268428
rect 159357 268018 159423 268021
rect 156676 268016 159423 268018
rect 156676 267960 159362 268016
rect 159418 267960 159423 268016
rect 156676 267958 159423 267960
rect 159357 267955 159423 267958
rect 198273 268018 198339 268021
rect 246798 268018 246804 268020
rect 198273 268016 200284 268018
rect 198273 267960 198278 268016
rect 198334 267960 200284 268016
rect 198273 267958 200284 267960
rect 244076 267958 246804 268018
rect 198273 267955 198339 267958
rect 246798 267956 246804 267958
rect 246868 267956 246874 268020
rect 67214 267412 67220 267476
rect 67284 267474 67290 267476
rect 246614 267474 246620 267476
rect 67284 267414 68908 267474
rect 244076 267414 246620 267474
rect 67284 267412 67290 267414
rect 246614 267412 246620 267414
rect 246684 267412 246690 267476
rect -960 267202 480 267292
rect 3141 267202 3207 267205
rect -960 267200 3207 267202
rect -960 267144 3146 267200
rect 3202 267144 3207 267200
rect -960 267142 3207 267144
rect -960 267052 480 267142
rect 3141 267139 3207 267142
rect 197537 267202 197603 267205
rect 197537 267200 200284 267202
rect 197537 267144 197542 267200
rect 197598 267144 200284 267200
rect 197537 267142 200284 267144
rect 197537 267139 197603 267142
rect 170857 267066 170923 267069
rect 184197 267066 184263 267069
rect 170857 267064 184263 267066
rect 170857 267008 170862 267064
rect 170918 267008 184202 267064
rect 184258 267008 184263 267064
rect 170857 267006 184263 267008
rect 170857 267003 170923 267006
rect 184197 267003 184263 267006
rect 246614 267004 246620 267068
rect 246684 267066 246690 267068
rect 277393 267066 277459 267069
rect 246684 267064 277459 267066
rect 246684 267008 277398 267064
rect 277454 267008 277459 267064
rect 246684 267006 277459 267008
rect 246684 267004 246690 267006
rect 277393 267003 277459 267006
rect 67766 266324 67772 266388
rect 67836 266386 67842 266388
rect 156646 266386 156706 266900
rect 197445 266658 197511 266661
rect 245745 266658 245811 266661
rect 197445 266656 200284 266658
rect 197445 266600 197450 266656
rect 197506 266600 200284 266656
rect 197445 266598 200284 266600
rect 244076 266656 245811 266658
rect 244076 266600 245750 266656
rect 245806 266600 245811 266656
rect 244076 266598 245811 266600
rect 197445 266595 197511 266598
rect 245745 266595 245811 266598
rect 170857 266386 170923 266389
rect 67836 266326 68908 266386
rect 156646 266384 170923 266386
rect 156646 266328 170862 266384
rect 170918 266328 170923 266384
rect 156646 266326 170923 266328
rect 67836 266324 67842 266326
rect 170857 266323 170923 266326
rect 261477 266386 261543 266389
rect 272425 266386 272491 266389
rect 261477 266384 272491 266386
rect 261477 266328 261482 266384
rect 261538 266328 272430 266384
rect 272486 266328 272491 266384
rect 261477 266326 272491 266328
rect 261477 266323 261543 266326
rect 272425 266323 272491 266326
rect 397361 266386 397427 266389
rect 583201 266386 583267 266389
rect 397361 266384 583267 266386
rect 397361 266328 397366 266384
rect 397422 266328 583206 266384
rect 583262 266328 583267 266384
rect 397361 266326 583267 266328
rect 397361 266323 397427 266326
rect 583201 266323 583267 266326
rect 158805 265842 158871 265845
rect 245837 265842 245903 265845
rect 156676 265840 158871 265842
rect 156676 265784 158810 265840
rect 158866 265784 158871 265840
rect 244076 265840 245903 265842
rect 156676 265782 158871 265784
rect 158805 265779 158871 265782
rect 195145 265570 195211 265573
rect 200254 265570 200314 265812
rect 244076 265784 245842 265840
rect 245898 265784 245903 265840
rect 244076 265782 245903 265784
rect 245837 265779 245903 265782
rect 195145 265568 200314 265570
rect 195145 265512 195150 265568
rect 195206 265512 200314 265568
rect 195145 265510 200314 265512
rect 195145 265507 195211 265510
rect 66805 265298 66871 265301
rect 246021 265298 246087 265301
rect 66805 265296 68908 265298
rect 66805 265240 66810 265296
rect 66866 265240 68908 265296
rect 66805 265238 68908 265240
rect 200070 265238 200284 265298
rect 244076 265296 246087 265298
rect 244076 265240 246026 265296
rect 246082 265240 246087 265296
rect 244076 265238 246087 265240
rect 66805 265235 66871 265238
rect 188337 265162 188403 265165
rect 200070 265162 200130 265238
rect 246021 265235 246087 265238
rect 188337 265160 200130 265162
rect 188337 265104 188342 265160
rect 188398 265104 200130 265160
rect 188337 265102 200130 265104
rect 188337 265099 188403 265102
rect 171041 265026 171107 265029
rect 195145 265026 195211 265029
rect 171041 265024 195211 265026
rect 171041 264968 171046 265024
rect 171102 264968 195150 265024
rect 195206 264968 195211 265024
rect 171041 264966 195211 264968
rect 171041 264963 171107 264966
rect 195145 264963 195211 264966
rect 257521 264890 257587 264893
rect 258073 264890 258139 264893
rect 257521 264888 258139 264890
rect 257521 264832 257526 264888
rect 257582 264832 258078 264888
rect 258134 264832 258139 264888
rect 257521 264830 258139 264832
rect 257521 264827 257587 264830
rect 258073 264827 258139 264830
rect 158805 264754 158871 264757
rect 258809 264754 258875 264757
rect 259361 264754 259427 264757
rect 156676 264752 158871 264754
rect 156676 264696 158810 264752
rect 158866 264696 158871 264752
rect 156676 264694 158871 264696
rect 158805 264691 158871 264694
rect 248370 264752 259427 264754
rect 248370 264696 258814 264752
rect 258870 264696 259366 264752
rect 259422 264696 259427 264752
rect 248370 264694 259427 264696
rect 197445 264482 197511 264485
rect 244457 264482 244523 264485
rect 197445 264480 200284 264482
rect 197445 264424 197450 264480
rect 197506 264424 200284 264480
rect 197445 264422 200284 264424
rect 244076 264480 244523 264482
rect 244076 264424 244462 264480
rect 244518 264424 244523 264480
rect 244076 264422 244523 264424
rect 197445 264419 197511 264422
rect 244457 264419 244523 264422
rect 66897 264210 66963 264213
rect 187233 264210 187299 264213
rect 197302 264210 197308 264212
rect 66897 264208 68908 264210
rect 66897 264152 66902 264208
rect 66958 264152 68908 264208
rect 66897 264150 68908 264152
rect 187233 264208 197308 264210
rect 187233 264152 187238 264208
rect 187294 264152 197308 264208
rect 187233 264150 197308 264152
rect 66897 264147 66963 264150
rect 187233 264147 187299 264150
rect 197302 264148 197308 264150
rect 197372 264148 197378 264212
rect 248370 264210 248430 264694
rect 258809 264691 258875 264694
rect 259361 264691 259427 264694
rect 244046 264150 248430 264210
rect 244046 263908 244106 264150
rect 186957 263802 187023 263805
rect 156646 263800 187023 263802
rect 156646 263744 186962 263800
rect 187018 263744 187023 263800
rect 156646 263742 187023 263744
rect 156646 263636 156706 263742
rect 186957 263739 187023 263742
rect 197445 263666 197511 263669
rect 197445 263664 200284 263666
rect 197445 263608 197450 263664
rect 197506 263608 200284 263664
rect 197445 263606 200284 263608
rect 197445 263603 197511 263606
rect 246798 263468 246804 263532
rect 246868 263530 246874 263532
rect 261477 263530 261543 263533
rect 246868 263528 261543 263530
rect 246868 263472 261482 263528
rect 261538 263472 261543 263528
rect 246868 263470 261543 263472
rect 246868 263468 246874 263470
rect 261477 263467 261543 263470
rect 66805 263122 66871 263125
rect 66805 263120 68908 263122
rect 66805 263064 66810 263120
rect 66866 263064 68908 263120
rect 66805 263062 68908 263064
rect 66805 263059 66871 263062
rect 197302 263060 197308 263124
rect 197372 263122 197378 263124
rect 197372 263062 200284 263122
rect 197372 263060 197378 263062
rect 167637 262850 167703 262853
rect 193806 262850 193812 262852
rect 167637 262848 193812 262850
rect 167637 262792 167642 262848
rect 167698 262792 193812 262848
rect 167637 262790 193812 262792
rect 167637 262787 167703 262790
rect 193806 262788 193812 262790
rect 193876 262788 193882 262852
rect 158805 262578 158871 262581
rect 156676 262576 158871 262578
rect 156676 262520 158810 262576
rect 158866 262520 158871 262576
rect 156676 262518 158871 262520
rect 244046 262578 244106 263092
rect 272425 262850 272491 262853
rect 396809 262850 396875 262853
rect 397361 262850 397427 262853
rect 272425 262848 397427 262850
rect 272425 262792 272430 262848
rect 272486 262792 396814 262848
rect 396870 262792 397366 262848
rect 397422 262792 397427 262848
rect 272425 262790 397427 262792
rect 272425 262787 272491 262790
rect 396809 262787 396875 262790
rect 397361 262787 397427 262790
rect 244222 262578 244228 262580
rect 244046 262518 244228 262578
rect 158805 262515 158871 262518
rect 244222 262516 244228 262518
rect 244292 262516 244298 262580
rect 198457 262306 198523 262309
rect 245837 262306 245903 262309
rect 198457 262304 200284 262306
rect 198457 262248 198462 262304
rect 198518 262248 200284 262304
rect 198457 262246 200284 262248
rect 244076 262304 245903 262306
rect 244076 262248 245842 262304
rect 245898 262248 245903 262304
rect 244076 262246 245903 262248
rect 198457 262243 198523 262246
rect 245837 262243 245903 262246
rect 66253 262034 66319 262037
rect 66253 262032 68908 262034
rect 66253 261976 66258 262032
rect 66314 261976 68908 262032
rect 66253 261974 68908 261976
rect 66253 261971 66319 261974
rect 156822 261700 156828 261764
rect 156892 261762 156898 261764
rect 167085 261762 167151 261765
rect 244365 261762 244431 261765
rect 156892 261760 167151 261762
rect 156892 261704 167090 261760
rect 167146 261704 167151 261760
rect 156892 261702 167151 261704
rect 244076 261760 244431 261762
rect 244076 261704 244370 261760
rect 244426 261704 244431 261760
rect 244076 261702 244431 261704
rect 156892 261700 156898 261702
rect 167085 261699 167151 261702
rect 244365 261699 244431 261702
rect 158621 261490 158687 261493
rect 156676 261488 158687 261490
rect 156676 261432 158626 261488
rect 158682 261432 158687 261488
rect 156676 261430 158687 261432
rect 158621 261427 158687 261430
rect 197445 261490 197511 261493
rect 197445 261488 200284 261490
rect 197445 261432 197450 261488
rect 197506 261432 200284 261488
rect 197445 261430 200284 261432
rect 197445 261427 197511 261430
rect 66805 260946 66871 260949
rect 198089 260946 198155 260949
rect 247125 260946 247191 260949
rect 249742 260946 249748 260948
rect 66805 260944 68908 260946
rect 66805 260888 66810 260944
rect 66866 260888 68908 260944
rect 66805 260886 68908 260888
rect 198089 260944 200284 260946
rect 198089 260888 198094 260944
rect 198150 260888 200284 260944
rect 198089 260886 200284 260888
rect 244076 260944 249748 260946
rect 244076 260888 247130 260944
rect 247186 260888 249748 260944
rect 244076 260886 249748 260888
rect 66805 260883 66871 260886
rect 198089 260883 198155 260886
rect 247125 260883 247191 260886
rect 249742 260884 249748 260886
rect 249812 260884 249818 260948
rect 158897 260402 158963 260405
rect 159214 260402 159220 260404
rect 156676 260400 159220 260402
rect 156676 260344 158902 260400
rect 158958 260344 159220 260400
rect 156676 260342 159220 260344
rect 158897 260339 158963 260342
rect 159214 260340 159220 260342
rect 159284 260340 159290 260404
rect 197445 260130 197511 260133
rect 246021 260130 246087 260133
rect 197445 260128 200284 260130
rect 197445 260072 197450 260128
rect 197506 260072 200284 260128
rect 197445 260070 200284 260072
rect 244076 260128 246087 260130
rect 244076 260072 246026 260128
rect 246082 260072 246087 260128
rect 244076 260070 246087 260072
rect 197445 260067 197511 260070
rect 246021 260067 246087 260070
rect 65977 259858 66043 259861
rect 65977 259856 68908 259858
rect 65977 259800 65982 259856
rect 66038 259800 68908 259856
rect 65977 259798 68908 259800
rect 65977 259795 66043 259798
rect 244406 259586 244412 259588
rect 244076 259526 244412 259586
rect 244406 259524 244412 259526
rect 244476 259586 244482 259588
rect 245653 259586 245719 259589
rect 244476 259584 245719 259586
rect 244476 259528 245658 259584
rect 245714 259528 245719 259584
rect 244476 259526 245719 259528
rect 244476 259524 244482 259526
rect 245653 259523 245719 259526
rect 195094 259450 195100 259452
rect 156646 259390 195100 259450
rect 156646 259284 156706 259390
rect 195094 259388 195100 259390
rect 195164 259388 195170 259452
rect 197445 259314 197511 259317
rect 243997 259314 244063 259317
rect 197445 259312 200284 259314
rect 197445 259256 197450 259312
rect 197506 259256 200284 259312
rect 197445 259254 200284 259256
rect 243997 259312 244106 259314
rect 243997 259256 244002 259312
rect 244058 259256 244106 259312
rect 197445 259251 197511 259254
rect 243997 259251 244106 259256
rect 66253 258090 66319 258093
rect 66253 258088 66362 258090
rect 66253 258032 66258 258088
rect 66314 258032 66362 258088
rect 66253 258027 66362 258032
rect 66302 257954 66362 258027
rect 68878 257954 68938 258740
rect 191598 258708 191604 258772
rect 191668 258770 191674 258772
rect 244046 258770 244106 259251
rect 582833 258906 582899 258909
rect 583520 258906 584960 258996
rect 582833 258904 584960 258906
rect 582833 258848 582838 258904
rect 582894 258848 584960 258904
rect 582833 258846 584960 258848
rect 582833 258843 582899 258846
rect 245653 258770 245719 258773
rect 191668 258710 200284 258770
rect 244046 258768 245719 258770
rect 244046 258740 245658 258768
rect 244076 258712 245658 258740
rect 245714 258712 245719 258768
rect 583520 258756 584960 258846
rect 244076 258710 245719 258712
rect 191668 258708 191674 258710
rect 245653 258707 245719 258710
rect 158805 258226 158871 258229
rect 245837 258226 245903 258229
rect 156676 258224 158871 258226
rect 156676 258168 158810 258224
rect 158866 258168 158871 258224
rect 156676 258166 158871 258168
rect 244076 258224 245903 258226
rect 244076 258168 245842 258224
rect 245898 258168 245903 258224
rect 244076 258166 245903 258168
rect 158805 258163 158871 258166
rect 245837 258163 245903 258166
rect 66302 257894 68938 257954
rect 197445 257954 197511 257957
rect 197445 257952 200284 257954
rect 197445 257896 197450 257952
rect 197506 257896 200284 257952
rect 197445 257894 200284 257896
rect 197445 257891 197511 257894
rect 66897 257682 66963 257685
rect 66897 257680 68908 257682
rect 66897 257624 66902 257680
rect 66958 257624 68908 257680
rect 66897 257622 68908 257624
rect 66897 257619 66963 257622
rect 197537 257410 197603 257413
rect 245837 257410 245903 257413
rect 197537 257408 200284 257410
rect 197537 257352 197542 257408
rect 197598 257352 200284 257408
rect 197537 257350 200284 257352
rect 244076 257408 245903 257410
rect 244076 257352 245842 257408
rect 245898 257352 245903 257408
rect 244076 257350 245903 257352
rect 197537 257347 197603 257350
rect 245837 257347 245903 257350
rect 159265 257138 159331 257141
rect 156676 257136 159331 257138
rect 156676 257080 159270 257136
rect 159326 257080 159331 257136
rect 156676 257078 159331 257080
rect 159265 257075 159331 257078
rect 197445 256594 197511 256597
rect 245837 256594 245903 256597
rect 197445 256592 200284 256594
rect 69430 256052 69490 256564
rect 197445 256536 197450 256592
rect 197506 256536 200284 256592
rect 197445 256534 200284 256536
rect 244076 256592 245903 256594
rect 244076 256536 245842 256592
rect 245898 256536 245903 256592
rect 244076 256534 245903 256536
rect 197445 256531 197511 256534
rect 245837 256531 245903 256534
rect 158805 256322 158871 256325
rect 156676 256320 158871 256322
rect 156676 256264 158810 256320
rect 158866 256264 158871 256320
rect 156676 256262 158871 256264
rect 158805 256259 158871 256262
rect 69422 255988 69428 256052
rect 69492 255988 69498 256052
rect 245837 256050 245903 256053
rect 244076 256048 245903 256050
rect 244076 255992 245842 256048
rect 245898 255992 245903 256048
rect 244076 255990 245903 255992
rect 245837 255987 245903 255990
rect 191046 255580 191052 255644
rect 191116 255642 191122 255644
rect 196934 255642 196940 255644
rect 191116 255582 196940 255642
rect 191116 255580 191122 255582
rect 196934 255580 196940 255582
rect 197004 255580 197010 255644
rect 66805 255506 66871 255509
rect 170489 255506 170555 255509
rect 200254 255506 200314 255748
rect 66805 255504 68908 255506
rect 66805 255448 66810 255504
rect 66866 255448 68908 255504
rect 66805 255446 68908 255448
rect 170489 255504 200314 255506
rect 170489 255448 170494 255504
rect 170550 255448 200314 255504
rect 170489 255446 200314 255448
rect 66805 255443 66871 255446
rect 170489 255443 170555 255446
rect 170949 255370 171015 255373
rect 193213 255370 193279 255373
rect 194409 255370 194475 255373
rect 170949 255368 194475 255370
rect 170949 255312 170954 255368
rect 171010 255312 193218 255368
rect 193274 255312 194414 255368
rect 194470 255312 194475 255368
rect 170949 255310 194475 255312
rect 170949 255307 171015 255310
rect 193213 255307 193279 255310
rect 194409 255307 194475 255310
rect 158897 255234 158963 255237
rect 156676 255232 158963 255234
rect 156676 255176 158902 255232
rect 158958 255176 158963 255232
rect 156676 255174 158963 255176
rect 158897 255171 158963 255174
rect 197445 255234 197511 255237
rect 245837 255234 245903 255237
rect 197445 255232 200284 255234
rect 197445 255176 197450 255232
rect 197506 255176 200284 255232
rect 197445 255174 200284 255176
rect 244076 255232 245903 255234
rect 244076 255176 245842 255232
rect 245898 255176 245903 255232
rect 244076 255174 245903 255176
rect 197445 255171 197511 255174
rect 245837 255171 245903 255174
rect 157977 254554 158043 254557
rect 167085 254554 167151 254557
rect 157977 254552 167151 254554
rect 157977 254496 157982 254552
rect 158038 254496 167090 254552
rect 167146 254496 167151 254552
rect 157977 254494 167151 254496
rect 157977 254491 158043 254494
rect 167085 254491 167151 254494
rect 66805 254418 66871 254421
rect 196893 254418 196959 254421
rect 246021 254418 246087 254421
rect 66805 254416 68908 254418
rect 66805 254360 66810 254416
rect 66866 254360 68908 254416
rect 66805 254358 68908 254360
rect 196893 254416 200284 254418
rect 196893 254360 196898 254416
rect 196954 254360 200284 254416
rect 196893 254358 200284 254360
rect 244076 254416 246087 254418
rect 244076 254360 246026 254416
rect 246082 254360 246087 254416
rect 244076 254358 246087 254360
rect 66805 254355 66871 254358
rect 196893 254355 196959 254358
rect 246021 254355 246087 254358
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect 158805 254146 158871 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect 156676 254144 158871 254146
rect 156676 254088 158810 254144
rect 158866 254088 158871 254144
rect 156676 254086 158871 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 158805 254083 158871 254086
rect 243486 254084 243492 254148
rect 243556 254084 243562 254148
rect 243494 253874 243554 254084
rect 245653 253874 245719 253877
rect 243494 253872 245719 253874
rect 243494 253844 245658 253872
rect 243524 253816 245658 253844
rect 245714 253816 245719 253872
rect 243524 253814 245719 253816
rect 245653 253811 245719 253814
rect 197905 253602 197971 253605
rect 197905 253600 200284 253602
rect 197905 253544 197910 253600
rect 197966 253544 200284 253600
rect 197905 253542 200284 253544
rect 197905 253539 197971 253542
rect 66805 253330 66871 253333
rect 66805 253328 68908 253330
rect 66805 253272 66810 253328
rect 66866 253272 68908 253328
rect 66805 253270 68908 253272
rect 66805 253267 66871 253270
rect 158805 253058 158871 253061
rect 156676 253056 158871 253058
rect 156676 253000 158810 253056
rect 158866 253000 158871 253056
rect 156676 252998 158871 253000
rect 158805 252995 158871 252998
rect 197445 253058 197511 253061
rect 246021 253058 246087 253061
rect 197445 253056 200284 253058
rect 197445 253000 197450 253056
rect 197506 253000 200284 253056
rect 197445 252998 200284 253000
rect 244076 253056 246087 253058
rect 244076 253000 246026 253056
rect 246082 253000 246087 253056
rect 244076 252998 246087 253000
rect 197445 252995 197511 252998
rect 246021 252995 246087 252998
rect 66662 252180 66668 252244
rect 66732 252242 66738 252244
rect 198641 252242 198707 252245
rect 199510 252242 199516 252244
rect 66732 252182 68908 252242
rect 198641 252240 199516 252242
rect 198641 252184 198646 252240
rect 198702 252184 199516 252240
rect 198641 252182 199516 252184
rect 66732 252180 66738 252182
rect 198641 252179 198707 252182
rect 199510 252180 199516 252182
rect 199580 252242 199586 252244
rect 245837 252242 245903 252245
rect 199580 252182 200284 252242
rect 244076 252240 245903 252242
rect 244076 252184 245842 252240
rect 245898 252184 245903 252240
rect 244076 252182 245903 252184
rect 199580 252180 199586 252182
rect 245837 252179 245903 252182
rect 158897 251970 158963 251973
rect 156676 251968 158963 251970
rect 156676 251912 158902 251968
rect 158958 251912 158963 251968
rect 156676 251910 158963 251912
rect 158897 251907 158963 251910
rect 244038 251908 244044 251972
rect 244108 251970 244114 251972
rect 289905 251970 289971 251973
rect 291101 251970 291167 251973
rect 244108 251968 291167 251970
rect 244108 251912 289910 251968
rect 289966 251912 291106 251968
rect 291162 251912 291167 251968
rect 244108 251910 291167 251912
rect 244108 251908 244114 251910
rect 289905 251907 289971 251910
rect 291101 251907 291167 251910
rect 167637 251834 167703 251837
rect 194777 251834 194843 251837
rect 167637 251832 194843 251834
rect 167637 251776 167642 251832
rect 167698 251776 194782 251832
rect 194838 251776 194843 251832
rect 167637 251774 194843 251776
rect 167637 251771 167703 251774
rect 194777 251771 194843 251774
rect 251081 251834 251147 251837
rect 298829 251834 298895 251837
rect 251081 251832 298895 251834
rect 251081 251776 251086 251832
rect 251142 251776 298834 251832
rect 298890 251776 298895 251832
rect 251081 251774 298895 251776
rect 251081 251771 251147 251774
rect 298829 251771 298895 251774
rect 197077 251698 197143 251701
rect 246021 251698 246087 251701
rect 197077 251696 200284 251698
rect 197077 251640 197082 251696
rect 197138 251640 200284 251696
rect 197077 251638 200284 251640
rect 244076 251696 246087 251698
rect 244076 251640 246026 251696
rect 246082 251640 246087 251696
rect 244076 251638 246087 251640
rect 197077 251635 197143 251638
rect 246021 251635 246087 251638
rect 67541 251154 67607 251157
rect 67541 251152 68908 251154
rect 67541 251096 67546 251152
rect 67602 251096 68908 251152
rect 67541 251094 68908 251096
rect 67541 251091 67607 251094
rect 158805 250882 158871 250885
rect 156676 250880 158871 250882
rect 156676 250824 158810 250880
rect 158866 250824 158871 250880
rect 156676 250822 158871 250824
rect 158805 250819 158871 250822
rect 197445 250882 197511 250885
rect 245653 250882 245719 250885
rect 197445 250880 200284 250882
rect 197445 250824 197450 250880
rect 197506 250824 200284 250880
rect 197445 250822 200284 250824
rect 244076 250880 245719 250882
rect 244076 250824 245658 250880
rect 245714 250824 245719 250880
rect 244076 250822 245719 250824
rect 197445 250819 197511 250822
rect 245653 250819 245719 250822
rect 178769 250474 178835 250477
rect 199469 250474 199535 250477
rect 178769 250472 199535 250474
rect 178769 250416 178774 250472
rect 178830 250416 199474 250472
rect 199530 250416 199535 250472
rect 178769 250414 199535 250416
rect 178769 250411 178835 250414
rect 199469 250411 199535 250414
rect 247309 250338 247375 250341
rect 244076 250336 247375 250338
rect 244076 250280 247314 250336
rect 247370 250280 247375 250336
rect 244076 250278 247375 250280
rect 247309 250275 247375 250278
rect 67817 250066 67883 250069
rect 197261 250066 197327 250069
rect 67817 250064 68908 250066
rect 67817 250008 67822 250064
rect 67878 250008 68908 250064
rect 67817 250006 68908 250008
rect 197261 250064 200284 250066
rect 197261 250008 197266 250064
rect 197322 250008 200284 250064
rect 197261 250006 200284 250008
rect 67817 250003 67883 250006
rect 197261 250003 197327 250006
rect 243486 250004 243492 250068
rect 243556 250066 243562 250068
rect 307753 250066 307819 250069
rect 243556 250064 307819 250066
rect 243556 250008 307758 250064
rect 307814 250008 307819 250064
rect 243556 250006 307819 250008
rect 243556 250004 243562 250006
rect 307753 250003 307819 250006
rect 158805 249794 158871 249797
rect 156676 249792 158871 249794
rect 156676 249736 158810 249792
rect 158866 249736 158871 249792
rect 156676 249734 158871 249736
rect 158805 249731 158871 249734
rect 197445 249522 197511 249525
rect 200021 249522 200087 249525
rect 246021 249522 246087 249525
rect 197445 249520 200284 249522
rect 197445 249464 197450 249520
rect 197506 249464 200026 249520
rect 200082 249464 200284 249520
rect 197445 249462 200284 249464
rect 244076 249520 246087 249522
rect 244076 249464 246026 249520
rect 246082 249464 246087 249520
rect 244076 249462 246087 249464
rect 197445 249459 197511 249462
rect 200021 249459 200087 249462
rect 246021 249459 246087 249462
rect 158897 249250 158963 249253
rect 172462 249250 172468 249252
rect 158897 249248 172468 249250
rect 158897 249192 158902 249248
rect 158958 249192 172468 249248
rect 158897 249190 172468 249192
rect 158897 249187 158963 249190
rect 172462 249188 172468 249190
rect 172532 249188 172538 249252
rect 168189 249114 168255 249117
rect 199326 249114 199332 249116
rect 168189 249112 199332 249114
rect 168189 249056 168194 249112
rect 168250 249056 199332 249112
rect 168189 249054 199332 249056
rect 168189 249051 168255 249054
rect 199326 249052 199332 249054
rect 199396 249052 199402 249116
rect 67173 248978 67239 248981
rect 67173 248976 68908 248978
rect 67173 248920 67178 248976
rect 67234 248920 68908 248976
rect 67173 248918 68908 248920
rect 67173 248915 67239 248918
rect 159449 248706 159515 248709
rect 156676 248704 159515 248706
rect 156676 248648 159454 248704
rect 159510 248648 159515 248704
rect 156676 248646 159515 248648
rect 159449 248643 159515 248646
rect 197445 248706 197511 248709
rect 247125 248706 247191 248709
rect 197445 248704 200284 248706
rect 197445 248648 197450 248704
rect 197506 248648 200284 248704
rect 197445 248646 200284 248648
rect 244076 248704 247191 248706
rect 244076 248648 247130 248704
rect 247186 248648 247191 248704
rect 244076 248646 247191 248648
rect 197445 248643 197511 248646
rect 247125 248643 247191 248646
rect 197721 247890 197787 247893
rect 197721 247888 200284 247890
rect 59118 247012 59124 247076
rect 59188 247074 59194 247076
rect 68878 247074 68938 247860
rect 197721 247832 197726 247888
rect 197782 247832 200284 247888
rect 197721 247830 200284 247832
rect 197721 247827 197787 247830
rect 160001 247618 160067 247621
rect 156676 247616 160067 247618
rect 156676 247560 160006 247616
rect 160062 247560 160067 247616
rect 156676 247558 160067 247560
rect 160001 247555 160067 247558
rect 177481 247618 177547 247621
rect 184841 247618 184907 247621
rect 244046 247618 244106 248132
rect 409873 247618 409939 247621
rect 583017 247618 583083 247621
rect 177481 247616 190470 247618
rect 177481 247560 177486 247616
rect 177542 247560 184846 247616
rect 184902 247560 190470 247616
rect 177481 247558 190470 247560
rect 244046 247558 248430 247618
rect 177481 247555 177547 247558
rect 184841 247555 184907 247558
rect 59188 247014 68938 247074
rect 190410 247074 190470 247558
rect 245837 247346 245903 247349
rect 244076 247344 245903 247346
rect 200254 247074 200314 247316
rect 244076 247288 245842 247344
rect 245898 247288 245903 247344
rect 244076 247286 245903 247288
rect 245837 247283 245903 247286
rect 190410 247014 200314 247074
rect 248370 247074 248430 247558
rect 409873 247616 583083 247618
rect 409873 247560 409878 247616
rect 409934 247560 583022 247616
rect 583078 247560 583083 247616
rect 409873 247558 583083 247560
rect 409873 247555 409939 247558
rect 583017 247555 583083 247558
rect 251817 247074 251883 247077
rect 262765 247074 262831 247077
rect 248370 247072 262831 247074
rect 248370 247016 251822 247072
rect 251878 247016 262770 247072
rect 262826 247016 262831 247072
rect 248370 247014 262831 247016
rect 59188 247012 59194 247014
rect 251817 247011 251883 247014
rect 262765 247011 262831 247014
rect 66805 246802 66871 246805
rect 66805 246800 68908 246802
rect 66805 246744 66810 246800
rect 66866 246744 68908 246800
rect 66805 246742 68908 246744
rect 66805 246739 66871 246742
rect 158805 246530 158871 246533
rect 156676 246528 158871 246530
rect 156676 246472 158810 246528
rect 158866 246472 158871 246528
rect 156676 246470 158871 246472
rect 158805 246467 158871 246470
rect 191649 246530 191715 246533
rect 198641 246530 198707 246533
rect 245694 246530 245700 246532
rect 191649 246528 200284 246530
rect 191649 246472 191654 246528
rect 191710 246472 198646 246528
rect 198702 246472 200284 246528
rect 191649 246470 200284 246472
rect 244076 246470 245700 246530
rect 191649 246467 191715 246470
rect 198641 246467 198707 246470
rect 245694 246468 245700 246470
rect 245764 246468 245770 246532
rect 298001 246394 298067 246397
rect 354029 246394 354095 246397
rect 298001 246392 354095 246394
rect 298001 246336 298006 246392
rect 298062 246336 354034 246392
rect 354090 246336 354095 246392
rect 298001 246334 354095 246336
rect 298001 246331 298067 246334
rect 354029 246331 354095 246334
rect 157926 246196 157932 246260
rect 157996 246258 158002 246260
rect 165061 246258 165127 246261
rect 157996 246256 165127 246258
rect 157996 246200 165066 246256
rect 165122 246200 165127 246256
rect 157996 246198 165127 246200
rect 157996 246196 158002 246198
rect 165061 246195 165127 246198
rect 282177 246258 282243 246261
rect 449157 246258 449223 246261
rect 282177 246256 449223 246258
rect 282177 246200 282182 246256
rect 282238 246200 449162 246256
rect 449218 246200 449223 246256
rect 282177 246198 449223 246200
rect 282177 246195 282243 246198
rect 449157 246195 449223 246198
rect 245653 245986 245719 245989
rect 200070 245926 200284 245986
rect 244076 245984 245719 245986
rect 244076 245928 245658 245984
rect 245714 245928 245719 245984
rect 244076 245926 245719 245928
rect 184289 245850 184355 245853
rect 186221 245850 186287 245853
rect 200070 245850 200130 245926
rect 245653 245923 245719 245926
rect 184289 245848 200130 245850
rect 184289 245792 184294 245848
rect 184350 245792 186226 245848
rect 186282 245792 200130 245848
rect 184289 245790 200130 245792
rect 253105 245850 253171 245853
rect 259729 245850 259795 245853
rect 260741 245850 260807 245853
rect 253105 245848 260807 245850
rect 253105 245792 253110 245848
rect 253166 245792 259734 245848
rect 259790 245792 260746 245848
rect 260802 245792 260807 245848
rect 253105 245790 260807 245792
rect 184289 245787 184355 245790
rect 186221 245787 186287 245790
rect 253105 245787 253171 245790
rect 259729 245787 259795 245790
rect 260741 245787 260807 245790
rect 66805 245714 66871 245717
rect 162301 245714 162367 245717
rect 191649 245714 191715 245717
rect 66805 245712 68908 245714
rect 66805 245656 66810 245712
rect 66866 245656 68908 245712
rect 66805 245654 68908 245656
rect 162301 245712 191715 245714
rect 162301 245656 162306 245712
rect 162362 245656 191654 245712
rect 191710 245656 191715 245712
rect 162301 245654 191715 245656
rect 66805 245651 66871 245654
rect 162301 245651 162367 245654
rect 191649 245651 191715 245654
rect 191782 245652 191788 245716
rect 191852 245714 191858 245716
rect 192201 245714 192267 245717
rect 191852 245712 192267 245714
rect 191852 245656 192206 245712
rect 192262 245656 192267 245712
rect 191852 245654 192267 245656
rect 191852 245652 191858 245654
rect 192201 245651 192267 245654
rect 245694 245652 245700 245716
rect 245764 245714 245770 245716
rect 298001 245714 298067 245717
rect 245764 245712 298067 245714
rect 245764 245656 298006 245712
rect 298062 245656 298067 245712
rect 245764 245654 298067 245656
rect 245764 245652 245770 245654
rect 298001 245651 298067 245654
rect 583017 245578 583083 245581
rect 583520 245578 584960 245668
rect 583017 245576 584960 245578
rect 583017 245520 583022 245576
rect 583078 245520 584960 245576
rect 583017 245518 584960 245520
rect 583017 245515 583083 245518
rect 158805 245442 158871 245445
rect 156676 245440 158871 245442
rect 156676 245384 158810 245440
rect 158866 245384 158871 245440
rect 583520 245428 584960 245518
rect 156676 245382 158871 245384
rect 158805 245379 158871 245382
rect 197353 245170 197419 245173
rect 246021 245170 246087 245173
rect 197353 245168 200284 245170
rect 197353 245112 197358 245168
rect 197414 245112 200284 245168
rect 197353 245110 200284 245112
rect 244076 245168 246087 245170
rect 244076 245112 246026 245168
rect 246082 245112 246087 245168
rect 244076 245110 246087 245112
rect 197353 245107 197419 245110
rect 246021 245107 246087 245110
rect 189717 244898 189783 244901
rect 199326 244898 199332 244900
rect 189717 244896 199332 244898
rect 189717 244840 189722 244896
rect 189778 244840 199332 244896
rect 189717 244838 199332 244840
rect 189717 244835 189783 244838
rect 199326 244836 199332 244838
rect 199396 244836 199402 244900
rect 66897 244626 66963 244629
rect 66897 244624 68908 244626
rect 66897 244568 66902 244624
rect 66958 244568 68908 244624
rect 66897 244566 68908 244568
rect 66897 244563 66963 244566
rect 156822 244564 156828 244628
rect 156892 244626 156898 244628
rect 191046 244626 191052 244628
rect 156892 244566 191052 244626
rect 156892 244564 156898 244566
rect 191046 244564 191052 244566
rect 191116 244626 191122 244628
rect 191782 244626 191788 244628
rect 191116 244566 191788 244626
rect 191116 244564 191122 244566
rect 191782 244564 191788 244566
rect 191852 244564 191858 244628
rect 158805 244354 158871 244357
rect 156676 244352 158871 244354
rect 156676 244296 158810 244352
rect 158866 244296 158871 244352
rect 156676 244294 158871 244296
rect 158805 244291 158871 244294
rect 198549 244354 198615 244357
rect 198549 244352 200652 244354
rect 198549 244296 198554 244352
rect 198610 244324 200652 244352
rect 198610 244296 200682 244324
rect 198549 244294 200682 244296
rect 198549 244291 198615 244294
rect 200622 244084 200682 244294
rect 244046 244221 244106 244596
rect 243997 244216 244106 244221
rect 243997 244160 244002 244216
rect 244058 244160 244106 244216
rect 243997 244158 244106 244160
rect 243997 244155 244063 244158
rect 200614 244020 200620 244084
rect 200684 244020 200690 244084
rect 197353 243810 197419 243813
rect 245745 243810 245811 243813
rect 197353 243808 200284 243810
rect 197353 243752 197358 243808
rect 197414 243752 200284 243808
rect 197353 243750 200284 243752
rect 244076 243808 245811 243810
rect 244076 243752 245750 243808
rect 245806 243752 245811 243808
rect 244076 243750 245811 243752
rect 197353 243747 197419 243750
rect 245745 243747 245811 243750
rect 67265 243540 67331 243541
rect 67214 243538 67220 243540
rect 67174 243478 67220 243538
rect 67284 243536 67331 243540
rect 67326 243480 67331 243536
rect 67214 243476 67220 243478
rect 67284 243476 67331 243480
rect 67265 243475 67331 243476
rect 67449 243538 67515 243541
rect 258717 243538 258783 243541
rect 319437 243538 319503 243541
rect 67449 243536 68908 243538
rect 67449 243480 67454 243536
rect 67510 243480 68908 243536
rect 67449 243478 68908 243480
rect 258030 243536 319503 243538
rect 258030 243480 258722 243536
rect 258778 243480 319442 243536
rect 319498 243480 319503 243536
rect 258030 243478 319503 243480
rect 67449 243475 67515 243478
rect 67541 243402 67607 243405
rect 69422 243402 69428 243404
rect 67541 243400 69428 243402
rect 67541 243344 67546 243400
rect 67602 243344 69428 243400
rect 67541 243342 69428 243344
rect 67541 243339 67607 243342
rect 69422 243340 69428 243342
rect 69492 243340 69498 243404
rect 158805 243266 158871 243269
rect 156676 243264 158871 243266
rect 156676 243208 158810 243264
rect 158866 243208 158871 243264
rect 156676 243206 158871 243208
rect 158805 243203 158871 243206
rect 165521 242994 165587 242997
rect 258030 242994 258090 243478
rect 258717 243475 258783 243478
rect 319437 243475 319503 243478
rect 165521 242992 200284 242994
rect 165521 242936 165526 242992
rect 165582 242936 200284 242992
rect 165521 242934 200284 242936
rect 244076 242934 258090 242994
rect 165521 242931 165587 242934
rect 156689 242858 156755 242861
rect 168189 242858 168255 242861
rect 156689 242856 168255 242858
rect 156689 242800 156694 242856
rect 156750 242800 168194 242856
rect 168250 242800 168255 242856
rect 156689 242798 168255 242800
rect 156689 242795 156755 242798
rect 168189 242795 168255 242798
rect 246113 242450 246179 242453
rect 244076 242448 246179 242450
rect 63125 242042 63191 242045
rect 63125 242040 64890 242042
rect 63125 241984 63130 242040
rect 63186 241984 64890 242040
rect 63125 241982 64890 241984
rect 63125 241979 63191 241982
rect 64830 241770 64890 241982
rect 69430 241906 69490 242420
rect 244076 242392 246118 242448
rect 246174 242392 246179 242448
rect 244076 242390 246179 242392
rect 246113 242387 246179 242390
rect 189073 242314 189139 242317
rect 199929 242314 199995 242317
rect 189073 242312 199995 242314
rect 189073 242256 189078 242312
rect 189134 242256 199934 242312
rect 199990 242256 199995 242312
rect 189073 242254 199995 242256
rect 189073 242251 189139 242254
rect 199929 242251 199995 242254
rect 158069 242178 158135 242181
rect 156676 242176 158135 242178
rect 156676 242120 158074 242176
rect 158130 242120 158135 242176
rect 156676 242118 158135 242120
rect 158069 242115 158135 242118
rect 165245 242178 165311 242181
rect 168373 242178 168439 242181
rect 192334 242178 192340 242180
rect 165245 242176 192340 242178
rect 165245 242120 165250 242176
rect 165306 242120 168378 242176
rect 168434 242120 192340 242176
rect 165245 242118 192340 242120
rect 165245 242115 165311 242118
rect 168373 242115 168439 242118
rect 192334 242116 192340 242118
rect 192404 242116 192410 242180
rect 198457 242178 198523 242181
rect 198457 242176 200284 242178
rect 198457 242120 198462 242176
rect 198518 242120 200284 242176
rect 198457 242118 200284 242120
rect 198457 242115 198523 242118
rect 80973 242044 81039 242045
rect 154665 242044 154731 242045
rect 80973 242042 81020 242044
rect 80928 242040 81020 242042
rect 80928 241984 80978 242040
rect 80928 241982 81020 241984
rect 80973 241980 81020 241982
rect 81084 241980 81090 242044
rect 154614 241980 154620 242044
rect 154684 242042 154731 242044
rect 154684 242040 154776 242042
rect 154726 241984 154776 242040
rect 154684 241982 154776 241984
rect 154684 241980 154731 241982
rect 80973 241979 81039 241980
rect 154665 241979 154731 241980
rect 69749 241906 69815 241909
rect 69430 241904 69815 241906
rect 69430 241848 69754 241904
rect 69810 241848 69815 241904
rect 69430 241846 69815 241848
rect 69749 241843 69815 241846
rect 69933 241770 69999 241773
rect 64830 241768 69999 241770
rect 64830 241712 69938 241768
rect 69994 241712 69999 241768
rect 64830 241710 69999 241712
rect 69933 241707 69999 241710
rect 191782 241572 191788 241636
rect 191852 241634 191858 241636
rect 245653 241634 245719 241637
rect 191852 241574 200284 241634
rect 244076 241632 245719 241634
rect 244076 241576 245658 241632
rect 245714 241576 245719 241632
rect 244076 241574 245719 241576
rect 191852 241572 191858 241574
rect 245653 241571 245719 241574
rect 18597 241498 18663 241501
rect 53649 241498 53715 241501
rect 138887 241498 138953 241501
rect 18597 241496 138953 241498
rect 18597 241440 18602 241496
rect 18658 241440 53654 241496
rect 53710 241440 138892 241496
rect 138948 241440 138953 241496
rect 18597 241438 138953 241440
rect 18597 241435 18663 241438
rect 53649 241435 53715 241438
rect 138887 241435 138953 241438
rect 156367 241498 156433 241501
rect 174629 241498 174695 241501
rect 156367 241496 174695 241498
rect 156367 241440 156372 241496
rect 156428 241440 174634 241496
rect 174690 241440 174695 241496
rect 156367 241438 174695 241440
rect 156367 241435 156433 241438
rect 174629 241435 174695 241438
rect 193857 241498 193923 241501
rect 195789 241498 195855 241501
rect 193857 241496 195855 241498
rect 193857 241440 193862 241496
rect 193918 241440 195794 241496
rect 195850 241440 195855 241496
rect 193857 241438 195855 241440
rect 193857 241435 193923 241438
rect 195789 241435 195855 241438
rect 83958 241300 83964 241364
rect 84028 241362 84034 241364
rect 93853 241362 93919 241365
rect 94911 241362 94977 241365
rect 84028 241360 94977 241362
rect 84028 241304 93858 241360
rect 93914 241304 94916 241360
rect 94972 241304 94977 241360
rect 84028 241302 94977 241304
rect 84028 241300 84034 241302
rect 93853 241299 93919 241302
rect 94911 241299 94977 241302
rect 108159 241362 108225 241365
rect 153101 241362 153167 241365
rect 108159 241360 153167 241362
rect 108159 241304 108164 241360
rect 108220 241304 153106 241360
rect 153162 241304 153167 241360
rect 108159 241302 153167 241304
rect 108159 241299 108225 241302
rect 153101 241299 153167 241302
rect 179413 241362 179479 241365
rect 180517 241362 180583 241365
rect 186313 241362 186379 241365
rect 179413 241360 186379 241362
rect 179413 241304 179418 241360
rect 179474 241304 180522 241360
rect 180578 241304 186318 241360
rect 186374 241304 186379 241360
rect 179413 241302 186379 241304
rect 179413 241299 179479 241302
rect 180517 241299 180583 241302
rect 186313 241299 186379 241302
rect 153009 241226 153075 241229
rect 156454 241226 156460 241228
rect 153009 241224 156460 241226
rect -960 241090 480 241180
rect 153009 241168 153014 241224
rect 153070 241168 156460 241224
rect 153009 241166 156460 241168
rect 153009 241163 153075 241166
rect 156454 241164 156460 241166
rect 156524 241164 156530 241228
rect 3325 241090 3391 241093
rect -960 241088 3391 241090
rect -960 241032 3330 241088
rect 3386 241032 3391 241088
rect -960 241030 3391 241032
rect -960 240940 480 241030
rect 3325 241027 3391 241030
rect 143441 241090 143507 241093
rect 156822 241090 156828 241092
rect 143441 241088 156828 241090
rect 143441 241032 143446 241088
rect 143502 241032 156828 241088
rect 143441 241030 156828 241032
rect 143441 241027 143507 241030
rect 156822 241028 156828 241030
rect 156892 241028 156898 241092
rect 69606 240756 69612 240820
rect 69676 240818 69682 240820
rect 77937 240818 78003 240821
rect 69676 240816 78003 240818
rect 69676 240760 77942 240816
rect 77998 240760 78003 240816
rect 69676 240758 78003 240760
rect 69676 240756 69682 240758
rect 77937 240755 78003 240758
rect 155677 240818 155743 240821
rect 164969 240818 165035 240821
rect 155677 240816 165035 240818
rect 155677 240760 155682 240816
rect 155738 240760 164974 240816
rect 165030 240760 165035 240816
rect 155677 240758 165035 240760
rect 155677 240755 155743 240758
rect 164969 240755 165035 240758
rect 197905 240818 197971 240821
rect 245837 240818 245903 240821
rect 302734 240818 302740 240820
rect 197905 240816 200284 240818
rect 197905 240760 197910 240816
rect 197966 240760 200284 240816
rect 197905 240758 200284 240760
rect 244076 240816 245903 240818
rect 244076 240760 245842 240816
rect 245898 240760 245903 240816
rect 244076 240758 245903 240760
rect 197905 240755 197971 240758
rect 245837 240755 245903 240758
rect 258030 240758 302740 240818
rect 173433 240546 173499 240549
rect 200113 240546 200179 240549
rect 173433 240544 200179 240546
rect 173433 240488 173438 240544
rect 173494 240488 200118 240544
rect 200174 240488 200179 240544
rect 173433 240486 200179 240488
rect 173433 240483 173499 240486
rect 200113 240483 200179 240486
rect 150801 240274 150867 240277
rect 153377 240274 153443 240277
rect 150801 240272 153443 240274
rect 150801 240216 150806 240272
rect 150862 240216 153382 240272
rect 153438 240216 153443 240272
rect 150801 240214 153443 240216
rect 150801 240211 150867 240214
rect 153377 240211 153443 240214
rect 192201 240274 192267 240277
rect 199837 240274 199903 240277
rect 255405 240274 255471 240277
rect 258030 240274 258090 240758
rect 302734 240756 302740 240758
rect 302804 240756 302810 240820
rect 192201 240272 199903 240274
rect 192201 240216 192206 240272
rect 192262 240216 199842 240272
rect 199898 240216 199903 240272
rect 192201 240214 199903 240216
rect 244076 240272 258090 240274
rect 244076 240216 255410 240272
rect 255466 240216 258090 240272
rect 244076 240214 258090 240216
rect 192201 240211 192267 240214
rect 199837 240211 199903 240214
rect 255405 240211 255471 240214
rect 49601 240138 49667 240141
rect 72417 240138 72483 240141
rect 72693 240138 72759 240141
rect 49601 240136 72759 240138
rect 49601 240080 49606 240136
rect 49662 240080 72422 240136
rect 72478 240080 72698 240136
rect 72754 240080 72759 240136
rect 49601 240078 72759 240080
rect 49601 240075 49667 240078
rect 72417 240075 72483 240078
rect 72693 240075 72759 240078
rect 157333 240138 157399 240141
rect 158478 240138 158484 240140
rect 157333 240136 158484 240138
rect 157333 240080 157338 240136
rect 157394 240080 158484 240136
rect 157333 240078 158484 240080
rect 157333 240075 157399 240078
rect 158478 240076 158484 240078
rect 158548 240076 158554 240140
rect 199929 240138 199995 240141
rect 200113 240138 200179 240141
rect 199929 240136 200179 240138
rect 199929 240080 199934 240136
rect 199990 240080 200118 240136
rect 200174 240080 200179 240136
rect 199929 240078 200179 240080
rect 199929 240075 199995 240078
rect 200113 240075 200179 240078
rect 207933 240138 207999 240141
rect 208158 240138 208164 240140
rect 207933 240136 208164 240138
rect 207933 240080 207938 240136
rect 207994 240080 208164 240136
rect 207933 240078 208164 240080
rect 207933 240075 207999 240078
rect 208158 240076 208164 240078
rect 208228 240076 208234 240140
rect 208301 240138 208367 240141
rect 210693 240140 210759 240141
rect 209630 240138 209636 240140
rect 208301 240136 209636 240138
rect 208301 240080 208306 240136
rect 208362 240080 209636 240136
rect 208301 240078 209636 240080
rect 208301 240075 208367 240078
rect 209630 240076 209636 240078
rect 209700 240076 209706 240140
rect 210693 240138 210740 240140
rect 210648 240136 210740 240138
rect 210648 240080 210698 240136
rect 210648 240078 210740 240080
rect 210693 240076 210740 240078
rect 210804 240076 210810 240140
rect 213085 240138 213151 240141
rect 213678 240138 213684 240140
rect 213085 240136 213684 240138
rect 213085 240080 213090 240136
rect 213146 240080 213684 240136
rect 213085 240078 213684 240080
rect 210693 240075 210759 240076
rect 213085 240075 213151 240078
rect 213678 240076 213684 240078
rect 213748 240076 213754 240140
rect 214189 240138 214255 240141
rect 217501 240140 217567 240141
rect 214598 240138 214604 240140
rect 214189 240136 214604 240138
rect 214189 240080 214194 240136
rect 214250 240080 214604 240136
rect 214189 240078 214604 240080
rect 214189 240075 214255 240078
rect 214598 240076 214604 240078
rect 214668 240076 214674 240140
rect 217501 240138 217548 240140
rect 217456 240136 217548 240138
rect 217456 240080 217506 240136
rect 217456 240078 217548 240080
rect 217501 240076 217548 240078
rect 217612 240076 217618 240140
rect 218973 240138 219039 240141
rect 220905 240140 220971 240141
rect 219198 240138 219204 240140
rect 218973 240136 219204 240138
rect 218973 240080 218978 240136
rect 219034 240080 219204 240136
rect 218973 240078 219204 240080
rect 217501 240075 217567 240076
rect 218973 240075 219039 240078
rect 219198 240076 219204 240078
rect 219268 240076 219274 240140
rect 220854 240076 220860 240140
rect 220924 240138 220971 240140
rect 224309 240138 224375 240141
rect 224718 240138 224724 240140
rect 220924 240136 221016 240138
rect 220966 240080 221016 240136
rect 220924 240078 221016 240080
rect 224309 240136 224724 240138
rect 224309 240080 224314 240136
rect 224370 240080 224724 240136
rect 224309 240078 224724 240080
rect 220924 240076 220971 240078
rect 220905 240075 220971 240076
rect 224309 240075 224375 240078
rect 224718 240076 224724 240078
rect 224788 240076 224794 240140
rect 226006 240076 226012 240140
rect 226076 240138 226082 240140
rect 228357 240138 228423 240141
rect 226076 240136 228423 240138
rect 226076 240080 228362 240136
rect 228418 240080 228423 240136
rect 226076 240078 228423 240080
rect 226076 240076 226082 240078
rect 228357 240075 228423 240078
rect 230422 240076 230428 240140
rect 230492 240138 230498 240140
rect 230565 240138 230631 240141
rect 230492 240136 230631 240138
rect 230492 240080 230570 240136
rect 230626 240080 230631 240136
rect 230492 240078 230631 240080
rect 230492 240076 230498 240078
rect 230565 240075 230631 240078
rect 232078 240076 232084 240140
rect 232148 240138 232154 240140
rect 232497 240138 232563 240141
rect 237465 240140 237531 240141
rect 232148 240136 232563 240138
rect 232148 240080 232502 240136
rect 232558 240080 232563 240136
rect 232148 240078 232563 240080
rect 232148 240076 232154 240078
rect 232497 240075 232563 240078
rect 237414 240076 237420 240140
rect 237484 240138 237531 240140
rect 237484 240136 237576 240138
rect 237526 240080 237576 240136
rect 237484 240078 237576 240080
rect 237484 240076 237531 240078
rect 241646 240076 241652 240140
rect 241716 240138 241722 240140
rect 242157 240138 242223 240141
rect 241716 240136 242223 240138
rect 241716 240080 242162 240136
rect 242218 240080 242223 240136
rect 241716 240078 242223 240080
rect 241716 240076 241722 240078
rect 237465 240075 237531 240076
rect 242157 240075 242223 240078
rect 65793 240002 65859 240005
rect 71037 240002 71103 240005
rect 65793 240000 71103 240002
rect 65793 239944 65798 240000
rect 65854 239944 71042 240000
rect 71098 239944 71103 240000
rect 65793 239942 71103 239944
rect 65793 239939 65859 239942
rect 71037 239939 71103 239942
rect 75545 240002 75611 240005
rect 98361 240002 98427 240005
rect 75545 240000 98427 240002
rect 75545 239944 75550 240000
rect 75606 239944 98366 240000
rect 98422 239944 98427 240000
rect 75545 239942 98427 239944
rect 75545 239939 75611 239942
rect 98361 239939 98427 239942
rect 152273 240002 152339 240005
rect 153101 240002 153167 240005
rect 158161 240002 158227 240005
rect 152273 240000 158227 240002
rect 152273 239944 152278 240000
rect 152334 239944 153106 240000
rect 153162 239944 158166 240000
rect 158222 239944 158227 240000
rect 152273 239942 158227 239944
rect 152273 239939 152339 239942
rect 153101 239939 153167 239942
rect 158161 239939 158227 239942
rect 236361 240002 236427 240005
rect 243302 240002 243308 240004
rect 236361 240000 243308 240002
rect 236361 239944 236366 240000
rect 236422 239944 243308 240000
rect 236361 239942 243308 239944
rect 236361 239939 236427 239942
rect 243302 239940 243308 239942
rect 243372 240002 243378 240004
rect 243629 240002 243695 240005
rect 243372 240000 243695 240002
rect 243372 239944 243634 240000
rect 243690 239944 243695 240000
rect 243372 239942 243695 239944
rect 243372 239940 243378 239942
rect 243629 239939 243695 239942
rect 220721 239866 220787 239869
rect 247309 239866 247375 239869
rect 220721 239864 247375 239866
rect 220721 239808 220726 239864
rect 220782 239808 247314 239864
rect 247370 239808 247375 239864
rect 220721 239806 247375 239808
rect 220721 239803 220787 239806
rect 247309 239803 247375 239806
rect 74073 239730 74139 239733
rect 121637 239730 121703 239733
rect 74073 239728 121703 239730
rect 74073 239672 74078 239728
rect 74134 239672 121642 239728
rect 121698 239672 121703 239728
rect 74073 239670 121703 239672
rect 74073 239667 74139 239670
rect 121637 239667 121703 239670
rect 184749 239730 184815 239733
rect 200573 239730 200639 239733
rect 184749 239728 200639 239730
rect 184749 239672 184754 239728
rect 184810 239672 200578 239728
rect 200634 239672 200639 239728
rect 184749 239670 200639 239672
rect 184749 239667 184815 239670
rect 200573 239667 200639 239670
rect 122281 239594 122347 239597
rect 213821 239594 213887 239597
rect 122281 239592 213887 239594
rect 122281 239536 122286 239592
rect 122342 239536 213826 239592
rect 213882 239536 213887 239592
rect 122281 239534 213887 239536
rect 122281 239531 122347 239534
rect 213821 239531 213887 239534
rect 71681 239458 71747 239461
rect 83549 239458 83615 239461
rect 71681 239456 83615 239458
rect 71681 239400 71686 239456
rect 71742 239400 83554 239456
rect 83610 239400 83615 239456
rect 71681 239398 83615 239400
rect 71681 239395 71747 239398
rect 83549 239395 83615 239398
rect 97441 239458 97507 239461
rect 209865 239458 209931 239461
rect 97441 239456 209931 239458
rect 97441 239400 97446 239456
rect 97502 239400 209870 239456
rect 209926 239400 209931 239456
rect 97441 239398 209931 239400
rect 97441 239395 97507 239398
rect 209865 239395 209931 239398
rect 322289 239458 322355 239461
rect 342989 239458 343055 239461
rect 322289 239456 343055 239458
rect 322289 239400 322294 239456
rect 322350 239400 342994 239456
rect 343050 239400 343055 239456
rect 322289 239398 343055 239400
rect 322289 239395 322355 239398
rect 342989 239395 343055 239398
rect 209630 238716 209636 238780
rect 209700 238778 209706 238780
rect 224769 238778 224835 238781
rect 209700 238776 224835 238778
rect 209700 238720 224774 238776
rect 224830 238720 224835 238776
rect 209700 238718 224835 238720
rect 209700 238716 209706 238718
rect 224769 238715 224835 238718
rect 234061 238778 234127 238781
rect 305085 238778 305151 238781
rect 234061 238776 305151 238778
rect 234061 238720 234066 238776
rect 234122 238720 305090 238776
rect 305146 238720 305151 238776
rect 234061 238718 305151 238720
rect 234061 238715 234127 238718
rect 305085 238715 305151 238718
rect 153377 238642 153443 238645
rect 161013 238642 161079 238645
rect 153377 238640 161079 238642
rect 153377 238584 153382 238640
rect 153438 238584 161018 238640
rect 161074 238584 161079 238640
rect 153377 238582 161079 238584
rect 153377 238579 153443 238582
rect 161013 238579 161079 238582
rect 205817 238642 205883 238645
rect 206870 238642 206876 238644
rect 205817 238640 206876 238642
rect 205817 238584 205822 238640
rect 205878 238584 206876 238640
rect 205817 238582 206876 238584
rect 205817 238579 205883 238582
rect 206870 238580 206876 238582
rect 206940 238580 206946 238644
rect 211245 238642 211311 238645
rect 212390 238642 212396 238644
rect 211245 238640 212396 238642
rect 211245 238584 211250 238640
rect 211306 238584 212396 238640
rect 211245 238582 212396 238584
rect 211245 238579 211311 238582
rect 212390 238580 212396 238582
rect 212460 238580 212466 238644
rect 183369 238506 183435 238509
rect 202137 238506 202203 238509
rect 183369 238504 202203 238506
rect 183369 238448 183374 238504
rect 183430 238448 202142 238504
rect 202198 238448 202203 238504
rect 183369 238446 202203 238448
rect 183369 238443 183435 238446
rect 202137 238443 202203 238446
rect 213821 238506 213887 238509
rect 226701 238506 226767 238509
rect 213821 238504 226767 238506
rect 213821 238448 213826 238504
rect 213882 238448 226706 238504
rect 226762 238448 226767 238504
rect 213821 238446 226767 238448
rect 213821 238443 213887 238446
rect 226701 238443 226767 238446
rect 69013 238370 69079 238373
rect 184749 238370 184815 238373
rect 69013 238368 184815 238370
rect 69013 238312 69018 238368
rect 69074 238312 184754 238368
rect 184810 238312 184815 238368
rect 69013 238310 184815 238312
rect 69013 238307 69079 238310
rect 184749 238307 184815 238310
rect 190269 238370 190335 238373
rect 201585 238370 201651 238373
rect 190269 238368 201651 238370
rect 190269 238312 190274 238368
rect 190330 238312 201590 238368
rect 201646 238312 201651 238368
rect 190269 238310 201651 238312
rect 190269 238307 190335 238310
rect 201585 238307 201651 238310
rect 209865 238370 209931 238373
rect 214189 238370 214255 238373
rect 209865 238368 214255 238370
rect 209865 238312 209870 238368
rect 209926 238312 214194 238368
rect 214250 238312 214255 238368
rect 209865 238310 214255 238312
rect 209865 238307 209931 238310
rect 214189 238307 214255 238310
rect 84193 238234 84259 238237
rect 208301 238234 208367 238237
rect 84193 238232 208367 238234
rect 84193 238176 84198 238232
rect 84254 238176 208306 238232
rect 208362 238176 208367 238232
rect 84193 238174 208367 238176
rect 84193 238171 84259 238174
rect 208301 238171 208367 238174
rect 229093 238098 229159 238101
rect 230473 238098 230539 238101
rect 244038 238098 244044 238100
rect 229093 238096 244044 238098
rect 229093 238040 229098 238096
rect 229154 238040 230478 238096
rect 230534 238040 244044 238096
rect 229093 238038 244044 238040
rect 229093 238035 229159 238038
rect 230473 238035 230539 238038
rect 244038 238036 244044 238038
rect 244108 238036 244114 238100
rect 64689 237962 64755 237965
rect 82813 237962 82879 237965
rect 64689 237960 82879 237962
rect 64689 237904 64694 237960
rect 64750 237904 82818 237960
rect 82874 237904 82879 237960
rect 64689 237902 82879 237904
rect 64689 237899 64755 237902
rect 82813 237899 82879 237902
rect 226701 237962 226767 237965
rect 259361 237962 259427 237965
rect 226701 237960 259427 237962
rect 226701 237904 226706 237960
rect 226762 237904 259366 237960
rect 259422 237904 259427 237960
rect 226701 237902 259427 237904
rect 226701 237899 226767 237902
rect 259361 237899 259427 237902
rect 261569 237962 261635 237965
rect 282177 237962 282243 237965
rect 261569 237960 282243 237962
rect 261569 237904 261574 237960
rect 261630 237904 282182 237960
rect 282238 237904 282243 237960
rect 261569 237902 282243 237904
rect 261569 237899 261635 237902
rect 282177 237899 282243 237902
rect 153009 237418 153075 237421
rect 154062 237418 154068 237420
rect 153009 237416 154068 237418
rect 153009 237360 153014 237416
rect 153070 237360 154068 237416
rect 153009 237358 154068 237360
rect 153009 237355 153075 237358
rect 154062 237356 154068 237358
rect 154132 237356 154138 237420
rect 198733 237418 198799 237421
rect 199510 237418 199516 237420
rect 198733 237416 199516 237418
rect 198733 237360 198738 237416
rect 198794 237360 199516 237416
rect 198733 237358 199516 237360
rect 198733 237355 198799 237358
rect 199510 237356 199516 237358
rect 199580 237356 199586 237420
rect 209957 237418 210023 237421
rect 210693 237418 210759 237421
rect 211245 237418 211311 237421
rect 209957 237416 210759 237418
rect 209957 237360 209962 237416
rect 210018 237360 210698 237416
rect 210754 237360 210759 237416
rect 209957 237358 210759 237360
rect 209957 237355 210023 237358
rect 210693 237355 210759 237358
rect 211110 237416 211311 237418
rect 211110 237360 211250 237416
rect 211306 237360 211311 237416
rect 211110 237358 211311 237360
rect 76414 237220 76420 237284
rect 76484 237282 76490 237284
rect 102409 237282 102475 237285
rect 153285 237282 153351 237285
rect 155953 237282 156019 237285
rect 76484 237280 103530 237282
rect 76484 237224 102414 237280
rect 102470 237224 103530 237280
rect 76484 237222 103530 237224
rect 76484 237220 76490 237222
rect 102409 237219 102475 237222
rect 103470 236874 103530 237222
rect 153285 237280 156019 237282
rect 153285 237224 153290 237280
rect 153346 237224 155958 237280
rect 156014 237224 156019 237280
rect 153285 237222 156019 237224
rect 153285 237219 153351 237222
rect 155953 237219 156019 237222
rect 200113 237282 200179 237285
rect 205357 237282 205423 237285
rect 200113 237280 205423 237282
rect 200113 237224 200118 237280
rect 200174 237224 205362 237280
rect 205418 237224 205423 237280
rect 200113 237222 205423 237224
rect 200113 237219 200179 237222
rect 205357 237219 205423 237222
rect 209037 237282 209103 237285
rect 211110 237282 211170 237358
rect 211245 237355 211311 237358
rect 216438 237356 216444 237420
rect 216508 237418 216514 237420
rect 216581 237418 216647 237421
rect 216508 237416 216647 237418
rect 216508 237360 216586 237416
rect 216642 237360 216647 237416
rect 216508 237358 216647 237360
rect 216508 237356 216514 237358
rect 216581 237355 216647 237358
rect 216765 237418 216831 237421
rect 217501 237418 217567 237421
rect 216765 237416 217567 237418
rect 216765 237360 216770 237416
rect 216826 237360 217506 237416
rect 217562 237360 217567 237416
rect 216765 237358 217567 237360
rect 216765 237355 216831 237358
rect 217501 237355 217567 237358
rect 223614 237356 223620 237420
rect 223684 237418 223690 237420
rect 224309 237418 224375 237421
rect 223684 237416 224375 237418
rect 223684 237360 224314 237416
rect 224370 237360 224375 237416
rect 223684 237358 224375 237360
rect 223684 237356 223690 237358
rect 224309 237355 224375 237358
rect 230565 237418 230631 237421
rect 231761 237418 231827 237421
rect 230565 237416 231827 237418
rect 230565 237360 230570 237416
rect 230626 237360 231766 237416
rect 231822 237360 231827 237416
rect 230565 237358 231827 237360
rect 230565 237355 230631 237358
rect 231761 237355 231827 237358
rect 241789 237418 241855 237421
rect 242014 237418 242020 237420
rect 241789 237416 242020 237418
rect 241789 237360 241794 237416
rect 241850 237360 242020 237416
rect 241789 237358 242020 237360
rect 241789 237355 241855 237358
rect 242014 237356 242020 237358
rect 242084 237356 242090 237420
rect 242801 237418 242867 237421
rect 322289 237418 322355 237421
rect 242801 237416 322355 237418
rect 242801 237360 242806 237416
rect 242862 237360 322294 237416
rect 322350 237360 322355 237416
rect 242801 237358 322355 237360
rect 242801 237355 242867 237358
rect 322289 237355 322355 237358
rect 209037 237280 211170 237282
rect 209037 237224 209042 237280
rect 209098 237224 211170 237280
rect 209037 237222 211170 237224
rect 209037 237219 209103 237222
rect 218646 237220 218652 237284
rect 218716 237282 218722 237284
rect 221457 237282 221523 237285
rect 218716 237280 221523 237282
rect 218716 237224 221462 237280
rect 221518 237224 221523 237280
rect 218716 237222 221523 237224
rect 218716 237220 218722 237222
rect 221457 237219 221523 237222
rect 240685 237282 240751 237285
rect 342897 237282 342963 237285
rect 240685 237280 342963 237282
rect 240685 237224 240690 237280
rect 240746 237224 342902 237280
rect 342958 237224 342963 237280
rect 240685 237222 342963 237224
rect 240685 237219 240751 237222
rect 342897 237219 342963 237222
rect 136817 237146 136883 237149
rect 165245 237146 165311 237149
rect 136817 237144 165311 237146
rect 136817 237088 136822 237144
rect 136878 237088 165250 237144
rect 165306 237088 165311 237144
rect 136817 237086 165311 237088
rect 136817 237083 136883 237086
rect 165245 237083 165311 237086
rect 193806 237084 193812 237148
rect 193876 237146 193882 237148
rect 201309 237146 201375 237149
rect 193876 237144 201375 237146
rect 193876 237088 201314 237144
rect 201370 237088 201375 237144
rect 193876 237086 201375 237088
rect 193876 237084 193882 237086
rect 201309 237083 201375 237086
rect 242709 237146 242775 237149
rect 269941 237146 270007 237149
rect 242709 237144 270007 237146
rect 242709 237088 242714 237144
rect 242770 237088 269946 237144
rect 270002 237088 270007 237144
rect 242709 237086 270007 237088
rect 242709 237083 242775 237086
rect 269941 237083 270007 237086
rect 154665 237010 154731 237013
rect 238293 237010 238359 237013
rect 154665 237008 238359 237010
rect 154665 236952 154670 237008
rect 154726 236952 238298 237008
rect 238354 236952 238359 237008
rect 154665 236950 238359 236952
rect 154665 236947 154731 236950
rect 238293 236947 238359 236950
rect 122097 236874 122163 236877
rect 103470 236872 122163 236874
rect 103470 236816 122102 236872
rect 122158 236816 122163 236872
rect 103470 236814 122163 236816
rect 122097 236811 122163 236814
rect 192334 236812 192340 236876
rect 192404 236874 192410 236876
rect 242617 236874 242683 236877
rect 192404 236872 242683 236874
rect 192404 236816 242622 236872
rect 242678 236816 242683 236872
rect 192404 236814 242683 236816
rect 192404 236812 192410 236814
rect 242617 236811 242683 236814
rect 109033 236738 109099 236741
rect 137277 236738 137343 236741
rect 109033 236736 137343 236738
rect 109033 236680 109038 236736
rect 109094 236680 137282 236736
rect 137338 236680 137343 236736
rect 109033 236678 137343 236680
rect 109033 236675 109099 236678
rect 137277 236675 137343 236678
rect 69933 236602 69999 236605
rect 149053 236602 149119 236605
rect 69933 236600 149119 236602
rect 69933 236544 69938 236600
rect 69994 236544 149058 236600
rect 149114 236544 149119 236600
rect 69933 236542 149119 236544
rect 69933 236539 69999 236542
rect 149053 236539 149119 236542
rect 149329 236058 149395 236061
rect 178769 236058 178835 236061
rect 178953 236058 179019 236061
rect 149329 236056 154682 236058
rect 149329 236000 149334 236056
rect 149390 236000 154682 236056
rect 149329 235998 154682 236000
rect 149329 235995 149395 235998
rect 82670 235860 82676 235924
rect 82740 235922 82746 235924
rect 89805 235922 89871 235925
rect 82740 235920 89871 235922
rect 82740 235864 89810 235920
rect 89866 235864 89871 235920
rect 82740 235862 89871 235864
rect 154622 235922 154682 235998
rect 155910 236056 179019 236058
rect 155910 236000 178774 236056
rect 178830 236000 178958 236056
rect 179014 236000 179019 236056
rect 155910 235998 179019 236000
rect 155910 235922 155970 235998
rect 178769 235995 178835 235998
rect 178953 235995 179019 235998
rect 154622 235862 155970 235922
rect 196801 235922 196867 235925
rect 204069 235922 204135 235925
rect 269757 235922 269823 235925
rect 270401 235922 270467 235925
rect 196801 235920 204135 235922
rect 196801 235864 196806 235920
rect 196862 235864 204074 235920
rect 204130 235864 204135 235920
rect 196801 235862 204135 235864
rect 82740 235860 82746 235862
rect 89805 235859 89871 235862
rect 196801 235859 196867 235862
rect 204069 235859 204135 235862
rect 238710 235920 270467 235922
rect 238710 235864 269762 235920
rect 269818 235864 270406 235920
rect 270462 235864 270467 235920
rect 238710 235862 270467 235864
rect 135345 235786 135411 235789
rect 163589 235786 163655 235789
rect 164141 235786 164207 235789
rect 135345 235784 164207 235786
rect 135345 235728 135350 235784
rect 135406 235728 163594 235784
rect 163650 235728 164146 235784
rect 164202 235728 164207 235784
rect 135345 235726 164207 235728
rect 135345 235723 135411 235726
rect 163589 235723 163655 235726
rect 164141 235723 164207 235726
rect 168281 235786 168347 235789
rect 195973 235786 196039 235789
rect 168281 235784 196039 235786
rect 168281 235728 168286 235784
rect 168342 235728 195978 235784
rect 196034 235728 196039 235784
rect 168281 235726 196039 235728
rect 168281 235723 168347 235726
rect 195973 235723 196039 235726
rect 201309 235786 201375 235789
rect 208853 235786 208919 235789
rect 201309 235784 208919 235786
rect 201309 235728 201314 235784
rect 201370 235728 208858 235784
rect 208914 235728 208919 235784
rect 201309 235726 208919 235728
rect 201309 235723 201375 235726
rect 208853 235723 208919 235726
rect 236545 235786 236611 235789
rect 238710 235786 238770 235862
rect 269757 235859 269823 235862
rect 270401 235859 270467 235862
rect 236545 235784 238770 235786
rect 236545 235728 236550 235784
rect 236606 235728 238770 235784
rect 236545 235726 238770 235728
rect 236545 235723 236611 235726
rect 137277 235650 137343 235653
rect 155677 235650 155743 235653
rect 137277 235648 155743 235650
rect 137277 235592 137282 235648
rect 137338 235592 155682 235648
rect 155738 235592 155743 235648
rect 137277 235590 155743 235592
rect 137277 235587 137343 235590
rect 155677 235587 155743 235590
rect 187141 235650 187207 235653
rect 236453 235650 236519 235653
rect 187141 235648 236519 235650
rect 187141 235592 187146 235648
rect 187202 235592 236458 235648
rect 236514 235592 236519 235648
rect 187141 235590 236519 235592
rect 187141 235587 187207 235590
rect 236453 235587 236519 235590
rect 104709 235514 104775 235517
rect 159541 235514 159607 235517
rect 104709 235512 159607 235514
rect 104709 235456 104714 235512
rect 104770 235456 159546 235512
rect 159602 235456 159607 235512
rect 104709 235454 159607 235456
rect 104709 235451 104775 235454
rect 159541 235451 159607 235454
rect 233734 235452 233740 235516
rect 233804 235514 233810 235516
rect 237373 235514 237439 235517
rect 237925 235514 237991 235517
rect 233804 235512 237991 235514
rect 233804 235456 237378 235512
rect 237434 235456 237930 235512
rect 237986 235456 237991 235512
rect 233804 235454 237991 235456
rect 233804 235452 233810 235454
rect 237373 235451 237439 235454
rect 237925 235451 237991 235454
rect 168281 235242 168347 235245
rect 184933 235242 184999 235245
rect 168281 235240 184999 235242
rect 168281 235184 168286 235240
rect 168342 235184 184938 235240
rect 184994 235184 184999 235240
rect 168281 235182 184999 235184
rect 168281 235179 168347 235182
rect 184933 235179 184999 235182
rect 191189 235242 191255 235245
rect 201309 235242 201375 235245
rect 191189 235240 201375 235242
rect 191189 235184 191194 235240
rect 191250 235184 201314 235240
rect 201370 235184 201375 235240
rect 191189 235182 201375 235184
rect 191189 235179 191255 235182
rect 201309 235179 201375 235182
rect 208853 234970 208919 234973
rect 209221 234970 209287 234973
rect 208853 234968 209287 234970
rect 208853 234912 208858 234968
rect 208914 234912 209226 234968
rect 209282 234912 209287 234968
rect 208853 234910 209287 234912
rect 208853 234907 208919 234910
rect 209221 234907 209287 234910
rect 89805 234698 89871 234701
rect 90357 234698 90423 234701
rect 89805 234696 90423 234698
rect 89805 234640 89810 234696
rect 89866 234640 90362 234696
rect 90418 234640 90423 234696
rect 89805 234638 90423 234640
rect 89805 234635 89871 234638
rect 90357 234635 90423 234638
rect 158621 234698 158687 234701
rect 159357 234698 159423 234701
rect 158621 234696 159423 234698
rect 158621 234640 158626 234696
rect 158682 234640 159362 234696
rect 159418 234640 159423 234696
rect 158621 234638 159423 234640
rect 158621 234635 158687 234638
rect 159357 234635 159423 234638
rect 205582 234636 205588 234700
rect 205652 234698 205658 234700
rect 218145 234698 218211 234701
rect 226149 234698 226215 234701
rect 205652 234638 215402 234698
rect 205652 234636 205658 234638
rect 82813 234562 82879 234565
rect 188337 234562 188403 234565
rect 82813 234560 188403 234562
rect 82813 234504 82818 234560
rect 82874 234504 188342 234560
rect 188398 234504 188403 234560
rect 82813 234502 188403 234504
rect 82813 234499 82879 234502
rect 188337 234499 188403 234502
rect 196750 234500 196756 234564
rect 196820 234562 196826 234564
rect 210417 234562 210483 234565
rect 196820 234560 210483 234562
rect 196820 234504 210422 234560
rect 210478 234504 210483 234560
rect 196820 234502 210483 234504
rect 215342 234562 215402 234638
rect 218145 234696 226215 234698
rect 218145 234640 218150 234696
rect 218206 234640 226154 234696
rect 226210 234640 226215 234696
rect 218145 234638 226215 234640
rect 218145 234635 218211 234638
rect 226149 234635 226215 234638
rect 233509 234698 233575 234701
rect 341609 234698 341675 234701
rect 233509 234696 341675 234698
rect 233509 234640 233514 234696
rect 233570 234640 341614 234696
rect 341670 234640 341675 234696
rect 233509 234638 341675 234640
rect 233509 234635 233575 234638
rect 341609 234635 341675 234638
rect 231485 234562 231551 234565
rect 324313 234562 324379 234565
rect 215342 234502 219450 234562
rect 196820 234500 196826 234502
rect 210417 234499 210483 234502
rect 106273 234426 106339 234429
rect 175917 234426 175983 234429
rect 106273 234424 175983 234426
rect 106273 234368 106278 234424
rect 106334 234368 175922 234424
rect 175978 234368 175983 234424
rect 106273 234366 175983 234368
rect 106273 234363 106339 234366
rect 175917 234363 175983 234366
rect 188838 234364 188844 234428
rect 188908 234426 188914 234428
rect 202045 234426 202111 234429
rect 202505 234426 202571 234429
rect 188908 234424 202571 234426
rect 188908 234368 202050 234424
rect 202106 234368 202510 234424
rect 202566 234368 202571 234424
rect 188908 234366 202571 234368
rect 219390 234426 219450 234502
rect 231485 234560 324379 234562
rect 231485 234504 231490 234560
rect 231546 234504 324318 234560
rect 324374 234504 324379 234560
rect 231485 234502 324379 234504
rect 231485 234499 231551 234502
rect 324313 234499 324379 234502
rect 258809 234426 258875 234429
rect 219390 234424 258875 234426
rect 219390 234368 258814 234424
rect 258870 234368 258875 234424
rect 219390 234366 258875 234368
rect 188908 234364 188914 234366
rect 202045 234363 202111 234366
rect 202505 234363 202571 234366
rect 258809 234363 258875 234366
rect 231853 234156 231919 234157
rect 231853 234154 231900 234156
rect 231772 234152 231900 234154
rect 231964 234154 231970 234156
rect 232998 234154 233004 234156
rect 231772 234096 231858 234152
rect 231772 234094 231900 234096
rect 231853 234092 231900 234094
rect 231964 234094 233004 234154
rect 231964 234092 231970 234094
rect 232998 234092 233004 234094
rect 233068 234092 233074 234156
rect 231853 234091 231919 234092
rect 43437 233882 43503 233885
rect 158713 233882 158779 233885
rect 43437 233880 158779 233882
rect 43437 233824 43442 233880
rect 43498 233824 158718 233880
rect 158774 233824 158779 233880
rect 43437 233822 158779 233824
rect 43437 233819 43503 233822
rect 158713 233819 158779 233822
rect 191598 233820 191604 233884
rect 191668 233882 191674 233884
rect 192661 233882 192727 233885
rect 191668 233880 192727 233882
rect 191668 233824 192666 233880
rect 192722 233824 192727 233880
rect 191668 233822 192727 233824
rect 191668 233820 191674 233822
rect 192661 233819 192727 233822
rect 192937 233882 193003 233885
rect 240041 233882 240107 233885
rect 241237 233882 241303 233885
rect 192937 233880 241303 233882
rect 192937 233824 192942 233880
rect 192998 233824 240046 233880
rect 240102 233824 241242 233880
rect 241298 233824 241303 233880
rect 192937 233822 241303 233824
rect 192937 233819 193003 233822
rect 240041 233819 240107 233822
rect 241237 233819 241303 233822
rect 162117 233338 162183 233341
rect 196065 233338 196131 233341
rect 162117 233336 196131 233338
rect 162117 233280 162122 233336
rect 162178 233280 196070 233336
rect 196126 233280 196131 233336
rect 162117 233278 196131 233280
rect 162117 233275 162183 233278
rect 196065 233275 196131 233278
rect 114645 233202 114711 233205
rect 220997 233202 221063 233205
rect 221641 233202 221707 233205
rect 114645 233200 221707 233202
rect 114645 233144 114650 233200
rect 114706 233144 221002 233200
rect 221058 233144 221646 233200
rect 221702 233144 221707 233200
rect 114645 233142 221707 233144
rect 114645 233139 114711 233142
rect 220997 233139 221063 233142
rect 221641 233139 221707 233142
rect 223389 233202 223455 233205
rect 230422 233202 230428 233204
rect 223389 233200 230428 233202
rect 223389 233144 223394 233200
rect 223450 233144 230428 233200
rect 223389 233142 230428 233144
rect 223389 233139 223455 233142
rect 230422 233140 230428 233142
rect 230492 233140 230498 233204
rect 52177 232658 52243 232661
rect 114277 232658 114343 232661
rect 52177 232656 114343 232658
rect 52177 232600 52182 232656
rect 52238 232600 114282 232656
rect 114338 232600 114343 232656
rect 52177 232598 114343 232600
rect 52177 232595 52243 232598
rect 114277 232595 114343 232598
rect 138013 232658 138079 232661
rect 149329 232658 149395 232661
rect 138013 232656 149395 232658
rect 138013 232600 138018 232656
rect 138074 232600 149334 232656
rect 149390 232600 149395 232656
rect 138013 232598 149395 232600
rect 138013 232595 138079 232598
rect 149329 232595 149395 232598
rect 193806 232596 193812 232660
rect 193876 232658 193882 232660
rect 249885 232658 249951 232661
rect 193876 232656 249951 232658
rect 193876 232600 249890 232656
rect 249946 232600 249951 232656
rect 193876 232598 249951 232600
rect 193876 232596 193882 232598
rect 249885 232595 249951 232598
rect 65977 232522 66043 232525
rect 155769 232522 155835 232525
rect 65977 232520 155835 232522
rect 65977 232464 65982 232520
rect 66038 232464 155774 232520
rect 155830 232464 155835 232520
rect 65977 232462 155835 232464
rect 65977 232459 66043 232462
rect 155769 232459 155835 232462
rect 196065 232522 196131 232525
rect 196893 232522 196959 232525
rect 352649 232522 352715 232525
rect 196065 232520 352715 232522
rect 196065 232464 196070 232520
rect 196126 232464 196898 232520
rect 196954 232464 352654 232520
rect 352710 232464 352715 232520
rect 196065 232462 352715 232464
rect 196065 232459 196131 232462
rect 196893 232459 196959 232462
rect 352649 232459 352715 232462
rect 583201 232386 583267 232389
rect 583520 232386 584960 232476
rect 583201 232384 584960 232386
rect 583201 232328 583206 232384
rect 583262 232328 584960 232384
rect 583201 232326 584960 232328
rect 583201 232323 583267 232326
rect 583520 232236 584960 232326
rect 152733 231978 152799 231981
rect 195237 231978 195303 231981
rect 152733 231976 195303 231978
rect 152733 231920 152738 231976
rect 152794 231920 195242 231976
rect 195298 231920 195303 231976
rect 152733 231918 195303 231920
rect 152733 231915 152799 231918
rect 195237 231915 195303 231918
rect 63217 231842 63283 231845
rect 180057 231842 180123 231845
rect 180609 231842 180675 231845
rect 63217 231840 180675 231842
rect 63217 231784 63222 231840
rect 63278 231784 180062 231840
rect 180118 231784 180614 231840
rect 180670 231784 180675 231840
rect 63217 231782 180675 231784
rect 63217 231779 63283 231782
rect 180057 231779 180123 231782
rect 180609 231779 180675 231782
rect 183277 231842 183343 231845
rect 242801 231842 242867 231845
rect 183277 231840 242867 231842
rect 183277 231784 183282 231840
rect 183338 231784 242806 231840
rect 242862 231784 242867 231840
rect 183277 231782 242867 231784
rect 183277 231779 183343 231782
rect 242801 231779 242867 231782
rect 163773 231706 163839 231709
rect 166206 231706 166212 231708
rect 163773 231704 166212 231706
rect 163773 231648 163778 231704
rect 163834 231648 166212 231704
rect 163773 231646 166212 231648
rect 163773 231643 163839 231646
rect 166206 231644 166212 231646
rect 166276 231644 166282 231708
rect 173157 231706 173223 231709
rect 219525 231706 219591 231709
rect 220353 231706 220419 231709
rect 173157 231704 220419 231706
rect 173157 231648 173162 231704
rect 173218 231648 219530 231704
rect 219586 231648 220358 231704
rect 220414 231648 220419 231704
rect 173157 231646 220419 231648
rect 173157 231643 173223 231646
rect 219525 231643 219591 231646
rect 220353 231643 220419 231646
rect 234981 231706 235047 231709
rect 234981 231704 258090 231706
rect 234981 231648 234986 231704
rect 235042 231648 258090 231704
rect 234981 231646 258090 231648
rect 234981 231643 235047 231646
rect 195237 231570 195303 231573
rect 205582 231570 205588 231572
rect 195237 231568 205588 231570
rect 195237 231512 195242 231568
rect 195298 231512 205588 231568
rect 195237 231510 205588 231512
rect 195237 231507 195303 231510
rect 205582 231508 205588 231510
rect 205652 231508 205658 231572
rect 155769 231298 155835 231301
rect 190453 231298 190519 231301
rect 155769 231296 190519 231298
rect 155769 231240 155774 231296
rect 155830 231240 190458 231296
rect 190514 231240 190519 231296
rect 155769 231238 190519 231240
rect 155769 231235 155835 231238
rect 190453 231235 190519 231238
rect 220169 231298 220235 231301
rect 233509 231298 233575 231301
rect 220169 231296 233575 231298
rect 220169 231240 220174 231296
rect 220230 231240 233514 231296
rect 233570 231240 233575 231296
rect 220169 231238 233575 231240
rect 220169 231235 220235 231238
rect 233509 231235 233575 231238
rect 119889 231162 119955 231165
rect 162209 231162 162275 231165
rect 119889 231160 162275 231162
rect 119889 231104 119894 231160
rect 119950 231104 162214 231160
rect 162270 231104 162275 231160
rect 119889 231102 162275 231104
rect 119889 231099 119955 231102
rect 161430 230621 161490 231102
rect 162209 231099 162275 231102
rect 225781 231162 225847 231165
rect 257429 231162 257495 231165
rect 225781 231160 257495 231162
rect 225781 231104 225786 231160
rect 225842 231104 257434 231160
rect 257490 231104 257495 231160
rect 225781 231102 257495 231104
rect 258030 231162 258090 231646
rect 262305 231162 262371 231165
rect 373257 231162 373323 231165
rect 258030 231160 373323 231162
rect 258030 231104 262310 231160
rect 262366 231104 373262 231160
rect 373318 231104 373323 231160
rect 258030 231102 373323 231104
rect 225781 231099 225847 231102
rect 257429 231099 257495 231102
rect 262305 231099 262371 231102
rect 373257 231099 373323 231102
rect 161381 230616 161490 230621
rect 161381 230560 161386 230616
rect 161442 230560 161490 230616
rect 161381 230558 161490 230560
rect 161381 230555 161447 230558
rect 58985 230482 59051 230485
rect 138013 230482 138079 230485
rect 58985 230480 138079 230482
rect 58985 230424 58990 230480
rect 59046 230424 138018 230480
rect 138074 230424 138079 230480
rect 58985 230422 138079 230424
rect 58985 230419 59051 230422
rect 138013 230419 138079 230422
rect 160093 230482 160159 230485
rect 161289 230482 161355 230485
rect 240685 230482 240751 230485
rect 160093 230480 240751 230482
rect 160093 230424 160098 230480
rect 160154 230424 161294 230480
rect 161350 230424 240690 230480
rect 240746 230424 240751 230480
rect 160093 230422 240751 230424
rect 160093 230419 160159 230422
rect 161289 230419 161355 230422
rect 240685 230419 240751 230422
rect 111793 230346 111859 230349
rect 113081 230346 113147 230349
rect 160870 230346 160876 230348
rect 111793 230344 160876 230346
rect 111793 230288 111798 230344
rect 111854 230288 113086 230344
rect 113142 230288 160876 230344
rect 111793 230286 160876 230288
rect 111793 230283 111859 230286
rect 113081 230283 113147 230286
rect 160870 230284 160876 230286
rect 160940 230284 160946 230348
rect 218145 230346 218211 230349
rect 218973 230346 219039 230349
rect 218145 230344 219039 230346
rect 218145 230288 218150 230344
rect 218206 230288 218978 230344
rect 219034 230288 219039 230344
rect 218145 230286 219039 230288
rect 218145 230283 218211 230286
rect 218973 230283 219039 230286
rect 238293 230346 238359 230349
rect 316125 230346 316191 230349
rect 316677 230346 316743 230349
rect 238293 230344 316743 230346
rect 238293 230288 238298 230344
rect 238354 230288 316130 230344
rect 316186 230288 316682 230344
rect 316738 230288 316743 230344
rect 238293 230286 316743 230288
rect 238293 230283 238359 230286
rect 316125 230283 316191 230286
rect 316677 230283 316743 230286
rect 135253 230210 135319 230213
rect 136541 230210 136607 230213
rect 175774 230210 175780 230212
rect 135253 230208 175780 230210
rect 135253 230152 135258 230208
rect 135314 230152 136546 230208
rect 136602 230152 175780 230208
rect 135253 230150 175780 230152
rect 135253 230147 135319 230150
rect 136541 230147 136607 230150
rect 175774 230148 175780 230150
rect 175844 230148 175850 230212
rect 97349 229802 97415 229805
rect 109677 229802 109743 229805
rect 97349 229800 109743 229802
rect 97349 229744 97354 229800
rect 97410 229744 109682 229800
rect 109738 229744 109743 229800
rect 97349 229742 109743 229744
rect 97349 229739 97415 229742
rect 109677 229739 109743 229742
rect 184289 229802 184355 229805
rect 198457 229802 198523 229805
rect 231894 229802 231900 229804
rect 184289 229800 231900 229802
rect 184289 229744 184294 229800
rect 184350 229744 198462 229800
rect 198518 229744 231900 229800
rect 184289 229742 231900 229744
rect 184289 229739 184355 229742
rect 198457 229739 198523 229742
rect 231894 229740 231900 229742
rect 231964 229740 231970 229804
rect 295333 229802 295399 229805
rect 412398 229802 412404 229804
rect 295333 229800 412404 229802
rect 295333 229744 295338 229800
rect 295394 229744 412404 229800
rect 295333 229742 412404 229744
rect 295333 229739 295399 229742
rect 412398 229740 412404 229742
rect 412468 229740 412474 229804
rect 11697 229122 11763 229125
rect 93853 229122 93919 229125
rect 94497 229122 94563 229125
rect 11697 229120 94563 229122
rect 11697 229064 11702 229120
rect 11758 229064 93858 229120
rect 93914 229064 94502 229120
rect 94558 229064 94563 229120
rect 11697 229062 94563 229064
rect 11697 229059 11763 229062
rect 93853 229059 93919 229062
rect 94497 229059 94563 229062
rect 142153 229122 142219 229125
rect 218145 229122 218211 229125
rect 142153 229120 218211 229122
rect 142153 229064 142158 229120
rect 142214 229064 218150 229120
rect 218206 229064 218211 229120
rect 142153 229062 218211 229064
rect 142153 229059 142219 229062
rect 218145 229059 218211 229062
rect 92381 228850 92447 228853
rect 157333 228850 157399 228853
rect 92381 228848 157399 228850
rect 92381 228792 92386 228848
rect 92442 228792 157338 228848
rect 157394 228792 157399 228848
rect 92381 228790 157399 228792
rect 92381 228787 92447 228790
rect 157333 228787 157399 228790
rect 199377 228850 199443 228853
rect 204437 228850 204503 228853
rect 199377 228848 204503 228850
rect 199377 228792 199382 228848
rect 199438 228792 204442 228848
rect 204498 228792 204503 228848
rect 199377 228790 204503 228792
rect 199377 228787 199443 228790
rect 204437 228787 204503 228790
rect 144177 228714 144243 228717
rect 193806 228714 193812 228716
rect 144177 228712 193812 228714
rect 144177 228656 144182 228712
rect 144238 228656 193812 228712
rect 144177 228654 193812 228656
rect 144177 228651 144243 228654
rect 193806 228652 193812 228654
rect 193876 228652 193882 228716
rect 145005 228578 145071 228581
rect 239397 228578 239463 228581
rect 145005 228576 239463 228578
rect 145005 228520 145010 228576
rect 145066 228520 239402 228576
rect 239458 228520 239463 228576
rect 145005 228518 239463 228520
rect 145005 228515 145071 228518
rect 239397 228515 239463 228518
rect 178033 228442 178099 228445
rect 179270 228442 179276 228444
rect 178033 228440 179276 228442
rect 178033 228384 178038 228440
rect 178094 228384 179276 228440
rect 178033 228382 179276 228384
rect 178033 228379 178099 228382
rect 179270 228380 179276 228382
rect 179340 228380 179346 228444
rect 191046 228380 191052 228444
rect 191116 228442 191122 228444
rect 244222 228442 244228 228444
rect 191116 228382 244228 228442
rect 191116 228380 191122 228382
rect 244222 228380 244228 228382
rect 244292 228380 244298 228444
rect 66662 228244 66668 228308
rect 66732 228306 66738 228308
rect 87597 228306 87663 228309
rect 66732 228304 87663 228306
rect 66732 228248 87602 228304
rect 87658 228248 87663 228304
rect 66732 228246 87663 228248
rect 66732 228244 66738 228246
rect 87597 228243 87663 228246
rect 102133 228306 102199 228309
rect 103421 228306 103487 228309
rect 144729 228306 144795 228309
rect 102133 228304 144795 228306
rect 102133 228248 102138 228304
rect 102194 228248 103426 228304
rect 103482 228248 144734 228304
rect 144790 228248 144795 228304
rect 102133 228246 144795 228248
rect 102133 228243 102199 228246
rect 103421 228243 103487 228246
rect 144729 228243 144795 228246
rect 218145 228306 218211 228309
rect 285765 228306 285831 228309
rect 218145 228304 285831 228306
rect 218145 228248 218150 228304
rect 218206 228248 285770 228304
rect 285826 228248 285831 228304
rect 218145 228246 285831 228248
rect 218145 228243 218211 228246
rect 285765 228243 285831 228246
rect -960 227884 480 228124
rect 91185 227762 91251 227765
rect 92381 227762 92447 227765
rect 91185 227760 92447 227762
rect 91185 227704 91190 227760
rect 91246 227704 92386 227760
rect 92442 227704 92447 227760
rect 91185 227702 92447 227704
rect 91185 227699 91251 227702
rect 92381 227699 92447 227702
rect 204437 227762 204503 227765
rect 204989 227762 205055 227765
rect 204437 227760 205055 227762
rect 204437 227704 204442 227760
rect 204498 227704 204994 227760
rect 205050 227704 205055 227760
rect 204437 227702 205055 227704
rect 204437 227699 204503 227702
rect 204989 227699 205055 227702
rect 144085 227626 144151 227629
rect 153009 227626 153075 227629
rect 208945 227626 209011 227629
rect 144085 227624 209011 227626
rect 144085 227568 144090 227624
rect 144146 227568 153014 227624
rect 153070 227568 208950 227624
rect 209006 227568 209011 227624
rect 144085 227566 209011 227568
rect 144085 227563 144151 227566
rect 153009 227563 153075 227566
rect 208945 227563 209011 227566
rect 10961 227082 11027 227085
rect 202321 227082 202387 227085
rect 10961 227080 202387 227082
rect 10961 227024 10966 227080
rect 11022 227024 202326 227080
rect 202382 227024 202387 227080
rect 10961 227022 202387 227024
rect 10961 227019 11027 227022
rect 202321 227019 202387 227022
rect 202505 227082 202571 227085
rect 414238 227082 414244 227084
rect 202505 227080 414244 227082
rect 202505 227024 202510 227080
rect 202566 227024 414244 227080
rect 202505 227022 414244 227024
rect 202505 227019 202571 227022
rect 414238 227020 414244 227022
rect 414308 227020 414314 227084
rect 66069 226946 66135 226949
rect 397453 226946 397519 226949
rect 66069 226944 397519 226946
rect 66069 226888 66074 226944
rect 66130 226888 397458 226944
rect 397514 226888 397519 226944
rect 66069 226886 397519 226888
rect 66069 226883 66135 226886
rect 397453 226883 397519 226886
rect 115933 226266 115999 226269
rect 143441 226266 143507 226269
rect 234061 226266 234127 226269
rect 115933 226264 122850 226266
rect 115933 226208 115938 226264
rect 115994 226208 122850 226264
rect 115933 226206 122850 226208
rect 115933 226203 115999 226206
rect 122790 226130 122850 226206
rect 143441 226264 234127 226266
rect 143441 226208 143446 226264
rect 143502 226208 234066 226264
rect 234122 226208 234127 226264
rect 143441 226206 234127 226208
rect 143441 226203 143507 226206
rect 234061 226203 234127 226206
rect 160686 226130 160692 226132
rect 122790 226070 160692 226130
rect 160686 226068 160692 226070
rect 160756 226068 160762 226132
rect 149145 225994 149211 225997
rect 184790 225994 184796 225996
rect 149145 225992 184796 225994
rect 149145 225936 149150 225992
rect 149206 225936 184796 225992
rect 149145 225934 184796 225936
rect 149145 225931 149211 225934
rect 184790 225932 184796 225934
rect 184860 225932 184866 225996
rect 221641 225722 221707 225725
rect 251817 225722 251883 225725
rect 221641 225720 251883 225722
rect 221641 225664 221646 225720
rect 221702 225664 251822 225720
rect 251878 225664 251883 225720
rect 221641 225662 251883 225664
rect 221641 225659 221707 225662
rect 251817 225659 251883 225662
rect 96521 225586 96587 225589
rect 147765 225586 147831 225589
rect 96521 225584 147831 225586
rect 96521 225528 96526 225584
rect 96582 225528 147770 225584
rect 147826 225528 147831 225584
rect 96521 225526 147831 225528
rect 96521 225523 96587 225526
rect 147765 225523 147831 225526
rect 184790 225524 184796 225588
rect 184860 225586 184866 225588
rect 298134 225586 298140 225588
rect 184860 225526 298140 225586
rect 184860 225524 184866 225526
rect 298134 225524 298140 225526
rect 298204 225586 298210 225588
rect 298461 225586 298527 225589
rect 298204 225584 298527 225586
rect 298204 225528 298466 225584
rect 298522 225528 298527 225584
rect 298204 225526 298527 225528
rect 298204 225524 298210 225526
rect 298461 225523 298527 225526
rect 95233 225042 95299 225045
rect 96521 225042 96587 225045
rect 95233 225040 96587 225042
rect 95233 224984 95238 225040
rect 95294 224984 96526 225040
rect 96582 224984 96587 225040
rect 95233 224982 96587 224984
rect 95233 224979 95299 224982
rect 96521 224979 96587 224982
rect 115933 225042 115999 225045
rect 117129 225042 117195 225045
rect 115933 225040 117195 225042
rect 115933 224984 115938 225040
rect 115994 224984 117134 225040
rect 117190 224984 117195 225040
rect 115933 224982 117195 224984
rect 115933 224979 115999 224982
rect 117129 224979 117195 224982
rect 215937 225042 216003 225045
rect 216070 225042 216076 225044
rect 215937 225040 216076 225042
rect 215937 224984 215942 225040
rect 215998 224984 216076 225040
rect 215937 224982 216076 224984
rect 215937 224979 216003 224982
rect 216070 224980 216076 224982
rect 216140 224980 216146 225044
rect 73061 224906 73127 224909
rect 159449 224906 159515 224909
rect 73061 224904 159515 224906
rect 73061 224848 73066 224904
rect 73122 224848 159454 224904
rect 159510 224848 159515 224904
rect 73061 224846 159515 224848
rect 73061 224843 73127 224846
rect 159449 224843 159515 224846
rect 195789 224906 195855 224909
rect 284937 224906 285003 224909
rect 195789 224904 285003 224906
rect 195789 224848 195794 224904
rect 195850 224848 284942 224904
rect 284998 224848 285003 224904
rect 195789 224846 285003 224848
rect 195789 224843 195855 224846
rect 284937 224843 285003 224846
rect 89529 224770 89595 224773
rect 166809 224770 166875 224773
rect 89529 224768 166875 224770
rect 89529 224712 89534 224768
rect 89590 224712 166814 224768
rect 166870 224712 166875 224768
rect 89529 224710 166875 224712
rect 89529 224707 89595 224710
rect 166809 224707 166875 224710
rect 129733 224634 129799 224637
rect 131021 224634 131087 224637
rect 171961 224634 172027 224637
rect 129733 224632 172027 224634
rect 129733 224576 129738 224632
rect 129794 224576 131026 224632
rect 131082 224576 171966 224632
rect 172022 224576 172027 224632
rect 129733 224574 172027 224576
rect 129733 224571 129799 224574
rect 131021 224571 131087 224574
rect 171961 224571 172027 224574
rect 171777 224362 171843 224365
rect 295977 224362 296043 224365
rect 171777 224360 296043 224362
rect 171777 224304 171782 224360
rect 171838 224304 295982 224360
rect 296038 224304 296043 224360
rect 171777 224302 296043 224304
rect 171777 224299 171843 224302
rect 295977 224299 296043 224302
rect 166809 224226 166875 224229
rect 323577 224226 323643 224229
rect 166809 224224 323643 224226
rect 166809 224168 166814 224224
rect 166870 224168 323582 224224
rect 323638 224168 323643 224224
rect 166809 224166 323643 224168
rect 166809 224163 166875 224166
rect 323577 224163 323643 224166
rect 115013 223546 115079 223549
rect 247217 223546 247283 223549
rect 115013 223544 247283 223546
rect 115013 223488 115018 223544
rect 115074 223488 247222 223544
rect 247278 223488 247283 223544
rect 115013 223486 247283 223488
rect 115013 223483 115079 223486
rect 247217 223483 247283 223486
rect 60365 223410 60431 223413
rect 169150 223410 169156 223412
rect 60365 223408 169156 223410
rect 60365 223352 60370 223408
rect 60426 223352 169156 223408
rect 60365 223350 169156 223352
rect 60365 223347 60431 223350
rect 169150 223348 169156 223350
rect 169220 223348 169226 223412
rect 199326 222940 199332 223004
rect 199396 223002 199402 223004
rect 296713 223002 296779 223005
rect 297909 223002 297975 223005
rect 199396 223000 297975 223002
rect 199396 222944 296718 223000
rect 296774 222944 297914 223000
rect 297970 222944 297975 223000
rect 199396 222942 297975 222944
rect 199396 222940 199402 222942
rect 296713 222939 296779 222942
rect 297909 222939 297975 222942
rect 67265 222866 67331 222869
rect 583569 222866 583635 222869
rect 67265 222864 583635 222866
rect 67265 222808 67270 222864
rect 67326 222808 583574 222864
rect 583630 222808 583635 222864
rect 67265 222806 583635 222808
rect 67265 222803 67331 222806
rect 583569 222803 583635 222806
rect 59077 222186 59143 222189
rect 235349 222186 235415 222189
rect 59077 222184 235415 222186
rect 59077 222128 59082 222184
rect 59138 222128 235354 222184
rect 235410 222128 235415 222184
rect 59077 222126 235415 222128
rect 59077 222123 59143 222126
rect 235349 222123 235415 222126
rect 56409 222050 56475 222053
rect 218053 222050 218119 222053
rect 56409 222048 218119 222050
rect 56409 221992 56414 222048
rect 56470 221992 218058 222048
rect 218114 221992 218119 222048
rect 56409 221990 218119 221992
rect 56409 221987 56475 221990
rect 218053 221987 218119 221990
rect 228173 222050 228239 222053
rect 267733 222050 267799 222053
rect 269021 222050 269087 222053
rect 228173 222048 269087 222050
rect 228173 221992 228178 222048
rect 228234 221992 267738 222048
rect 267794 221992 269026 222048
rect 269082 221992 269087 222048
rect 228173 221990 269087 221992
rect 228173 221987 228239 221990
rect 267733 221987 267799 221990
rect 269021 221987 269087 221990
rect 94497 221914 94563 221917
rect 195421 221914 195487 221917
rect 195830 221914 195836 221916
rect 94497 221912 195836 221914
rect 94497 221856 94502 221912
rect 94558 221856 195426 221912
rect 195482 221856 195836 221912
rect 94497 221854 195836 221856
rect 94497 221851 94563 221854
rect 195421 221851 195487 221854
rect 195830 221852 195836 221854
rect 195900 221852 195906 221916
rect 208945 221914 209011 221917
rect 320173 221914 320239 221917
rect 320633 221914 320699 221917
rect 208945 221912 320699 221914
rect 208945 221856 208950 221912
rect 209006 221856 320178 221912
rect 320234 221856 320638 221912
rect 320694 221856 320699 221912
rect 208945 221854 320699 221856
rect 208945 221851 209011 221854
rect 320173 221851 320239 221854
rect 320633 221851 320699 221854
rect 122097 220826 122163 220829
rect 233417 220826 233483 220829
rect 122097 220824 233483 220826
rect 122097 220768 122102 220824
rect 122158 220768 233422 220824
rect 233478 220768 233483 220824
rect 122097 220766 233483 220768
rect 122097 220763 122163 220766
rect 233417 220763 233483 220766
rect 76557 220690 76623 220693
rect 156505 220690 156571 220693
rect 76557 220688 156571 220690
rect 76557 220632 76562 220688
rect 76618 220632 156510 220688
rect 156566 220632 156571 220688
rect 76557 220630 156571 220632
rect 76557 220627 76623 220630
rect 156505 220627 156571 220630
rect 138657 220554 138723 220557
rect 190177 220554 190243 220557
rect 138657 220552 190243 220554
rect 138657 220496 138662 220552
rect 138718 220496 190182 220552
rect 190238 220496 190243 220552
rect 138657 220494 190243 220496
rect 138657 220491 138723 220494
rect 190177 220491 190243 220494
rect 192937 220282 193003 220285
rect 238753 220282 238819 220285
rect 192937 220280 238819 220282
rect 192937 220224 192942 220280
rect 192998 220224 238758 220280
rect 238814 220224 238819 220280
rect 192937 220222 238819 220224
rect 192937 220219 193003 220222
rect 238753 220219 238819 220222
rect 190310 220084 190316 220148
rect 190380 220146 190386 220148
rect 195421 220146 195487 220149
rect 190380 220144 195487 220146
rect 190380 220088 195426 220144
rect 195482 220088 195487 220144
rect 190380 220086 195487 220088
rect 190380 220084 190386 220086
rect 195421 220083 195487 220086
rect 210417 220146 210483 220149
rect 444373 220146 444439 220149
rect 210417 220144 444439 220146
rect 210417 220088 210422 220144
rect 210478 220088 444378 220144
rect 444434 220088 444439 220144
rect 210417 220086 444439 220088
rect 210417 220083 210483 220086
rect 444373 220083 444439 220086
rect 190177 219466 190243 219469
rect 192477 219466 192543 219469
rect 190177 219464 192543 219466
rect 190177 219408 190182 219464
rect 190238 219408 192482 219464
rect 192538 219408 192543 219464
rect 190177 219406 192543 219408
rect 190177 219403 190243 219406
rect 192477 219403 192543 219406
rect 56501 219330 56567 219333
rect 227621 219330 227687 219333
rect 56501 219328 227687 219330
rect 56501 219272 56506 219328
rect 56562 219272 227626 219328
rect 227682 219272 227687 219328
rect 56501 219270 227687 219272
rect 56501 219267 56567 219270
rect 227621 219267 227687 219270
rect 117405 219194 117471 219197
rect 170949 219194 171015 219197
rect 195237 219194 195303 219197
rect 267825 219194 267891 219197
rect 117405 219192 171150 219194
rect 117405 219136 117410 219192
rect 117466 219136 170954 219192
rect 171010 219136 171150 219192
rect 117405 219134 171150 219136
rect 117405 219131 117471 219134
rect 170949 219131 171015 219134
rect 171090 218650 171150 219134
rect 195237 219192 267891 219194
rect 195237 219136 195242 219192
rect 195298 219136 267830 219192
rect 267886 219136 267891 219192
rect 195237 219134 267891 219136
rect 195237 219131 195303 219134
rect 267690 218786 267750 219134
rect 267825 219131 267891 219134
rect 583293 219058 583359 219061
rect 583520 219058 584960 219148
rect 583293 219056 584960 219058
rect 583293 219000 583298 219056
rect 583354 219000 584960 219056
rect 583293 218998 584960 219000
rect 583293 218995 583359 218998
rect 583520 218908 584960 218998
rect 298737 218786 298803 218789
rect 267690 218784 298803 218786
rect 267690 218728 298742 218784
rect 298798 218728 298803 218784
rect 267690 218726 298803 218728
rect 298737 218723 298803 218726
rect 192569 218650 192635 218653
rect 171090 218648 192635 218650
rect 171090 218592 192574 218648
rect 192630 218592 192635 218648
rect 171090 218590 192635 218592
rect 192569 218587 192635 218590
rect 218053 218650 218119 218653
rect 234654 218650 234660 218652
rect 218053 218648 234660 218650
rect 218053 218592 218058 218648
rect 218114 218592 234660 218648
rect 218053 218590 234660 218592
rect 218053 218587 218119 218590
rect 234654 218588 234660 218590
rect 234724 218588 234730 218652
rect 263777 218650 263843 218653
rect 408585 218650 408651 218653
rect 263777 218648 408651 218650
rect 263777 218592 263782 218648
rect 263838 218592 408590 218648
rect 408646 218592 408651 218648
rect 263777 218590 408651 218592
rect 263777 218587 263843 218590
rect 408585 218587 408651 218590
rect 227069 218106 227135 218109
rect 227621 218106 227687 218109
rect 227069 218104 227687 218106
rect 227069 218048 227074 218104
rect 227130 218048 227626 218104
rect 227682 218048 227687 218104
rect 227069 218046 227687 218048
rect 227069 218043 227135 218046
rect 227621 218043 227687 218046
rect 176009 217970 176075 217973
rect 225229 217970 225295 217973
rect 176009 217968 225295 217970
rect 176009 217912 176014 217968
rect 176070 217912 225234 217968
rect 225290 217912 225295 217968
rect 176009 217910 225295 217912
rect 176009 217907 176075 217910
rect 225229 217907 225295 217910
rect 150341 217562 150407 217565
rect 169017 217562 169083 217565
rect 150341 217560 169083 217562
rect 150341 217504 150346 217560
rect 150402 217504 169022 217560
rect 169078 217504 169083 217560
rect 150341 217502 169083 217504
rect 150341 217499 150407 217502
rect 169017 217499 169083 217502
rect 77937 217426 78003 217429
rect 213821 217426 213887 217429
rect 77937 217424 213887 217426
rect 77937 217368 77942 217424
rect 77998 217368 213826 217424
rect 213882 217368 213887 217424
rect 77937 217366 213887 217368
rect 77937 217363 78003 217366
rect 213821 217363 213887 217366
rect 225597 217426 225663 217429
rect 231945 217426 232011 217429
rect 225597 217424 232011 217426
rect 225597 217368 225602 217424
rect 225658 217368 231950 217424
rect 232006 217368 232011 217424
rect 225597 217366 232011 217368
rect 225597 217363 225663 217366
rect 231945 217363 232011 217366
rect 112989 217290 113055 217293
rect 253054 217290 253060 217292
rect 112989 217288 253060 217290
rect 112989 217232 112994 217288
rect 113050 217232 253060 217288
rect 112989 217230 253060 217232
rect 112989 217227 113055 217230
rect 253054 217228 253060 217230
rect 253124 217228 253130 217292
rect 142797 216610 142863 216613
rect 272609 216610 272675 216613
rect 142797 216608 272675 216610
rect 142797 216552 142802 216608
rect 142858 216552 272614 216608
rect 272670 216552 272675 216608
rect 142797 216550 272675 216552
rect 142797 216547 142863 216550
rect 272609 216547 272675 216550
rect 109677 216474 109743 216477
rect 207105 216474 207171 216477
rect 109677 216472 207171 216474
rect 109677 216416 109682 216472
rect 109738 216416 207110 216472
rect 207166 216416 207171 216472
rect 109677 216414 207171 216416
rect 109677 216411 109743 216414
rect 207105 216411 207171 216414
rect 69606 216276 69612 216340
rect 69676 216338 69682 216340
rect 158069 216338 158135 216341
rect 69676 216336 158135 216338
rect 69676 216280 158074 216336
rect 158130 216280 158135 216336
rect 69676 216278 158135 216280
rect 69676 216276 69682 216278
rect 158069 216275 158135 216278
rect 207933 216066 207999 216069
rect 215293 216066 215359 216069
rect 207933 216064 215359 216066
rect 207933 216008 207938 216064
rect 207994 216008 215298 216064
rect 215354 216008 215359 216064
rect 207933 216006 215359 216008
rect 207933 216003 207999 216006
rect 215293 216003 215359 216006
rect 217133 216066 217199 216069
rect 233182 216066 233188 216068
rect 217133 216064 233188 216066
rect 217133 216008 217138 216064
rect 217194 216008 233188 216064
rect 217133 216006 233188 216008
rect 217133 216003 217199 216006
rect 233182 216004 233188 216006
rect 233252 216004 233258 216068
rect 86861 215930 86927 215933
rect 141417 215930 141483 215933
rect 86861 215928 141483 215930
rect 86861 215872 86866 215928
rect 86922 215872 141422 215928
rect 141478 215872 141483 215928
rect 86861 215870 141483 215872
rect 86861 215867 86927 215870
rect 141417 215867 141483 215870
rect 193857 215930 193923 215933
rect 224401 215930 224467 215933
rect 193857 215928 224467 215930
rect 193857 215872 193862 215928
rect 193918 215872 224406 215928
rect 224462 215872 224467 215928
rect 193857 215870 224467 215872
rect 193857 215867 193923 215870
rect 224401 215867 224467 215870
rect 225229 215930 225295 215933
rect 338849 215930 338915 215933
rect 225229 215928 338915 215930
rect 225229 215872 225234 215928
rect 225290 215872 338854 215928
rect 338910 215872 338915 215928
rect 225229 215870 338915 215872
rect 225229 215867 225295 215870
rect 338849 215867 338915 215870
rect 207105 215386 207171 215389
rect 207749 215386 207815 215389
rect 207105 215384 207815 215386
rect 207105 215328 207110 215384
rect 207166 215328 207754 215384
rect 207810 215328 207815 215384
rect 207105 215326 207815 215328
rect 207105 215323 207171 215326
rect 207749 215323 207815 215326
rect 272609 215386 272675 215389
rect 274081 215386 274147 215389
rect 272609 215384 274147 215386
rect 272609 215328 272614 215384
rect 272670 215328 274086 215384
rect 274142 215328 274147 215384
rect 272609 215326 274147 215328
rect 272609 215323 272675 215326
rect 274081 215323 274147 215326
rect 71037 215250 71103 215253
rect 209773 215250 209839 215253
rect 210509 215250 210575 215253
rect 222377 215252 222443 215253
rect 222326 215250 222332 215252
rect 71037 215248 210575 215250
rect 71037 215192 71042 215248
rect 71098 215192 209778 215248
rect 209834 215192 210514 215248
rect 210570 215192 210575 215248
rect 71037 215190 210575 215192
rect 222286 215190 222332 215250
rect 222396 215248 222443 215252
rect 222438 215192 222443 215248
rect 71037 215187 71103 215190
rect 209773 215187 209839 215190
rect 210509 215187 210575 215190
rect 222326 215188 222332 215190
rect 222396 215188 222443 215192
rect 222377 215187 222443 215188
rect 100937 215114 101003 215117
rect 102041 215114 102107 215117
rect 128261 215114 128327 215117
rect 228449 215114 228515 215117
rect 100937 215112 103530 215114
rect -960 214978 480 215068
rect 100937 215056 100942 215112
rect 100998 215056 102046 215112
rect 102102 215056 103530 215112
rect 100937 215054 103530 215056
rect 100937 215051 101003 215054
rect 102041 215051 102107 215054
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect 103470 214978 103530 215054
rect 128261 215112 228515 215114
rect 128261 215056 128266 215112
rect 128322 215056 228454 215112
rect 228510 215056 228515 215112
rect 128261 215054 228515 215056
rect 128261 215051 128327 215054
rect 228449 215051 228515 215054
rect 161974 214978 161980 214980
rect 103470 214918 161980 214978
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 161974 214916 161980 214918
rect 162044 214916 162050 214980
rect 232998 214780 233004 214844
rect 233068 214842 233074 214844
rect 245745 214842 245811 214845
rect 233068 214840 245811 214842
rect 233068 214784 245750 214840
rect 245806 214784 245811 214840
rect 233068 214782 245811 214784
rect 233068 214780 233074 214782
rect 245745 214779 245811 214782
rect 196709 214706 196775 214709
rect 400213 214706 400279 214709
rect 196709 214704 400279 214706
rect 196709 214648 196714 214704
rect 196770 214648 400218 214704
rect 400274 214648 400279 214704
rect 196709 214646 400279 214648
rect 196709 214643 196775 214646
rect 400213 214643 400279 214646
rect 215293 214570 215359 214573
rect 420177 214570 420243 214573
rect 215293 214568 420243 214570
rect 215293 214512 215298 214568
rect 215354 214512 420182 214568
rect 420238 214512 420243 214568
rect 215293 214510 420243 214512
rect 215293 214507 215359 214510
rect 420177 214507 420243 214510
rect 232078 214372 232084 214436
rect 232148 214434 232154 214436
rect 232497 214434 232563 214437
rect 232148 214432 232563 214434
rect 232148 214376 232502 214432
rect 232558 214376 232563 214432
rect 232148 214374 232563 214376
rect 232148 214372 232154 214374
rect 232497 214371 232563 214374
rect 229645 213890 229711 213893
rect 254025 213890 254091 213893
rect 229645 213888 254091 213890
rect 229645 213832 229650 213888
rect 229706 213832 254030 213888
rect 254086 213832 254091 213888
rect 229645 213830 254091 213832
rect 229645 213827 229711 213830
rect 254025 213827 254091 213830
rect 108297 213754 108363 213757
rect 150341 213754 150407 213757
rect 151077 213754 151143 213757
rect 108297 213752 151143 213754
rect 108297 213696 108302 213752
rect 108358 213696 150346 213752
rect 150402 213696 151082 213752
rect 151138 213696 151143 213752
rect 108297 213694 151143 213696
rect 108297 213691 108363 213694
rect 150341 213691 150407 213694
rect 151077 213691 151143 213694
rect 129641 213618 129707 213621
rect 230473 213618 230539 213621
rect 129641 213616 230539 213618
rect 129641 213560 129646 213616
rect 129702 213560 230478 213616
rect 230534 213560 230539 213616
rect 129641 213558 230539 213560
rect 129641 213555 129707 213558
rect 230473 213555 230539 213558
rect 15837 213210 15903 213213
rect 170397 213210 170463 213213
rect 250529 213210 250595 213213
rect 15837 213208 250595 213210
rect 15837 213152 15842 213208
rect 15898 213152 170402 213208
rect 170458 213152 250534 213208
rect 250590 213152 250595 213208
rect 15837 213150 250595 213152
rect 15837 213147 15903 213150
rect 170397 213147 170463 213150
rect 250529 213147 250595 213150
rect 85665 212530 85731 212533
rect 86861 212530 86927 212533
rect 178534 212530 178540 212532
rect 85665 212528 178540 212530
rect 85665 212472 85670 212528
rect 85726 212472 86866 212528
rect 86922 212472 178540 212528
rect 85665 212470 178540 212472
rect 85665 212467 85731 212470
rect 86861 212467 86927 212470
rect 178534 212468 178540 212470
rect 178604 212468 178610 212532
rect 100661 212394 100727 212397
rect 188981 212394 189047 212397
rect 100661 212392 190470 212394
rect 100661 212336 100666 212392
rect 100722 212336 188986 212392
rect 189042 212336 190470 212392
rect 100661 212334 190470 212336
rect 100661 212331 100727 212334
rect 188981 212331 189047 212334
rect 190410 212122 190470 212334
rect 301497 212122 301563 212125
rect 190410 212120 301563 212122
rect 190410 212064 301502 212120
rect 301558 212064 301563 212120
rect 190410 212062 301563 212064
rect 301497 212059 301563 212062
rect 187417 211986 187483 211989
rect 345749 211986 345815 211989
rect 187417 211984 345815 211986
rect 187417 211928 187422 211984
rect 187478 211928 345754 211984
rect 345810 211928 345815 211984
rect 187417 211926 345815 211928
rect 187417 211923 187483 211926
rect 345749 211923 345815 211926
rect 204989 211850 205055 211853
rect 439129 211850 439195 211853
rect 204989 211848 439195 211850
rect 204989 211792 204994 211848
rect 205050 211792 439134 211848
rect 439190 211792 439195 211848
rect 204989 211790 439195 211792
rect 204989 211787 205055 211790
rect 439129 211787 439195 211790
rect 223389 211170 223455 211173
rect 223614 211170 223620 211172
rect 223389 211168 223620 211170
rect 223389 211112 223394 211168
rect 223450 211112 223620 211168
rect 223389 211110 223620 211112
rect 223389 211107 223455 211110
rect 223614 211108 223620 211110
rect 223684 211108 223690 211172
rect 133689 211034 133755 211037
rect 163773 211034 163839 211037
rect 133689 211032 163839 211034
rect 133689 210976 133694 211032
rect 133750 210976 163778 211032
rect 163834 210976 163839 211032
rect 133689 210974 163839 210976
rect 133689 210971 133755 210974
rect 163773 210971 163839 210974
rect 213821 211034 213887 211037
rect 276749 211034 276815 211037
rect 213821 211032 276815 211034
rect 213821 210976 213826 211032
rect 213882 210976 276754 211032
rect 276810 210976 276815 211032
rect 213821 210974 276815 210976
rect 213821 210971 213887 210974
rect 276749 210971 276815 210974
rect 158713 210490 158779 210493
rect 237557 210490 237623 210493
rect 244365 210490 244431 210493
rect 158713 210488 244431 210490
rect 158713 210432 158718 210488
rect 158774 210432 237562 210488
rect 237618 210432 244370 210488
rect 244426 210432 244431 210488
rect 158713 210430 244431 210432
rect 158713 210427 158779 210430
rect 237557 210427 237623 210430
rect 244365 210427 244431 210430
rect 117313 210354 117379 210357
rect 223389 210354 223455 210357
rect 117313 210352 223455 210354
rect 117313 210296 117318 210352
rect 117374 210296 223394 210352
rect 223450 210296 223455 210352
rect 117313 210294 223455 210296
rect 117313 210291 117379 210294
rect 223389 210291 223455 210294
rect 396717 210354 396783 210357
rect 433374 210354 433380 210356
rect 396717 210352 433380 210354
rect 396717 210296 396722 210352
rect 396778 210296 433380 210352
rect 396717 210294 433380 210296
rect 396717 210291 396783 210294
rect 433374 210292 433380 210294
rect 433444 210292 433450 210356
rect 123477 209674 123543 209677
rect 242985 209674 243051 209677
rect 123477 209672 243051 209674
rect 123477 209616 123482 209672
rect 123538 209616 242990 209672
rect 243046 209616 243051 209672
rect 123477 209614 243051 209616
rect 123477 209611 123543 209614
rect 242985 209611 243051 209614
rect 122833 209538 122899 209541
rect 225689 209538 225755 209541
rect 122833 209536 225755 209538
rect 122833 209480 122838 209536
rect 122894 209480 225694 209536
rect 225750 209480 225755 209536
rect 122833 209478 225755 209480
rect 122833 209475 122899 209478
rect 225689 209475 225755 209478
rect 89713 209402 89779 209405
rect 91001 209402 91067 209405
rect 173014 209402 173020 209404
rect 89713 209400 173020 209402
rect 89713 209344 89718 209400
rect 89774 209344 91006 209400
rect 91062 209344 173020 209400
rect 89713 209342 173020 209344
rect 89713 209339 89779 209342
rect 91001 209339 91067 209342
rect 173014 209340 173020 209342
rect 173084 209340 173090 209404
rect 173801 208450 173867 208453
rect 423673 208450 423739 208453
rect 173801 208448 423739 208450
rect 173801 208392 173806 208448
rect 173862 208392 423678 208448
rect 423734 208392 423739 208448
rect 173801 208390 423739 208392
rect 173801 208387 173867 208390
rect 423673 208387 423739 208390
rect 63309 208314 63375 208317
rect 213177 208314 213243 208317
rect 63309 208312 213243 208314
rect 63309 208256 63314 208312
rect 63370 208256 213182 208312
rect 213238 208256 213243 208312
rect 63309 208254 213243 208256
rect 63309 208251 63375 208254
rect 213177 208251 213243 208254
rect 99281 208178 99347 208181
rect 99281 208176 238770 208178
rect 99281 208120 99286 208176
rect 99342 208120 238770 208176
rect 99281 208118 238770 208120
rect 99281 208115 99347 208118
rect 238710 207634 238770 208118
rect 240358 207634 240364 207636
rect 238710 207574 240364 207634
rect 240358 207572 240364 207574
rect 240428 207634 240434 207636
rect 251817 207634 251883 207637
rect 240428 207632 251883 207634
rect 240428 207576 251822 207632
rect 251878 207576 251883 207632
rect 240428 207574 251883 207576
rect 240428 207572 240434 207574
rect 251817 207571 251883 207574
rect 440233 207090 440299 207093
rect 216078 207088 440299 207090
rect 216078 207032 440238 207088
rect 440294 207032 440299 207088
rect 216078 207030 440299 207032
rect 216078 206957 216138 207030
rect 440233 207027 440299 207030
rect 69657 206954 69723 206957
rect 216029 206954 216138 206957
rect 69657 206952 216138 206954
rect 69657 206896 69662 206952
rect 69718 206896 216034 206952
rect 216090 206896 216138 206952
rect 69657 206894 216138 206896
rect 235901 206954 235967 206957
rect 264973 206954 265039 206957
rect 235901 206952 265039 206954
rect 235901 206896 235906 206952
rect 235962 206896 264978 206952
rect 265034 206896 265039 206952
rect 235901 206894 265039 206896
rect 69657 206891 69723 206894
rect 216029 206891 216095 206894
rect 235901 206891 235967 206894
rect 264973 206891 265039 206894
rect 182173 206818 182239 206821
rect 230381 206818 230447 206821
rect 232129 206818 232195 206821
rect 182173 206816 232195 206818
rect 182173 206760 182178 206816
rect 182234 206760 230386 206816
rect 230442 206760 232134 206816
rect 232190 206760 232195 206816
rect 182173 206758 232195 206760
rect 182173 206755 182239 206758
rect 230381 206755 230447 206758
rect 232129 206755 232195 206758
rect 91093 206274 91159 206277
rect 207289 206274 207355 206277
rect 209037 206274 209103 206277
rect 91093 206272 209103 206274
rect 91093 206216 91098 206272
rect 91154 206216 207294 206272
rect 207350 206216 209042 206272
rect 209098 206216 209103 206272
rect 91093 206214 209103 206216
rect 91093 206211 91159 206214
rect 207289 206211 207355 206214
rect 209037 206211 209103 206214
rect 209221 206274 209287 206277
rect 422937 206274 423003 206277
rect 209221 206272 423003 206274
rect 209221 206216 209226 206272
rect 209282 206216 422942 206272
rect 422998 206216 423003 206272
rect 209221 206214 423003 206216
rect 209221 206211 209287 206214
rect 422937 206211 423003 206214
rect 214465 205732 214531 205733
rect 214414 205730 214420 205732
rect 214374 205670 214420 205730
rect 214484 205728 214531 205732
rect 214526 205672 214531 205728
rect 214414 205668 214420 205670
rect 214484 205668 214531 205672
rect 214465 205667 214531 205668
rect 583385 205730 583451 205733
rect 583520 205730 584960 205820
rect 583385 205728 584960 205730
rect 583385 205672 583390 205728
rect 583446 205672 584960 205728
rect 583385 205670 584960 205672
rect 583385 205667 583451 205670
rect 83457 205594 83523 205597
rect 239397 205594 239463 205597
rect 239765 205594 239831 205597
rect 83457 205592 239831 205594
rect 83457 205536 83462 205592
rect 83518 205536 239402 205592
rect 239458 205536 239770 205592
rect 239826 205536 239831 205592
rect 583520 205580 584960 205670
rect 83457 205534 239831 205536
rect 83457 205531 83523 205534
rect 239397 205531 239463 205534
rect 239765 205531 239831 205534
rect 133137 205458 133203 205461
rect 209957 205458 210023 205461
rect 210417 205458 210483 205461
rect 133137 205456 210483 205458
rect 133137 205400 133142 205456
rect 133198 205400 209962 205456
rect 210018 205400 210422 205456
rect 210478 205400 210483 205456
rect 133137 205398 210483 205400
rect 133137 205395 133203 205398
rect 209957 205395 210023 205398
rect 210417 205395 210483 205398
rect 216438 205396 216444 205460
rect 216508 205458 216514 205460
rect 216508 205398 238770 205458
rect 216508 205396 216514 205398
rect 147581 205322 147647 205325
rect 147581 205320 161490 205322
rect 147581 205264 147586 205320
rect 147642 205264 161490 205320
rect 147581 205262 161490 205264
rect 147581 205259 147647 205262
rect 161430 204914 161490 205262
rect 238710 205050 238770 205398
rect 251265 205050 251331 205053
rect 320909 205050 320975 205053
rect 238710 205048 320975 205050
rect 238710 204992 251270 205048
rect 251326 204992 320914 205048
rect 320970 204992 320975 205048
rect 238710 204990 320975 204992
rect 251265 204987 251331 204990
rect 320909 204987 320975 204990
rect 172421 204914 172487 204917
rect 418889 204914 418955 204917
rect 161430 204912 418955 204914
rect 161430 204856 172426 204912
rect 172482 204856 418894 204912
rect 418950 204856 418955 204912
rect 161430 204854 418955 204856
rect 172421 204851 172487 204854
rect 418889 204851 418955 204854
rect 144913 204234 144979 204237
rect 238017 204234 238083 204237
rect 144913 204232 238083 204234
rect 144913 204176 144918 204232
rect 144974 204176 238022 204232
rect 238078 204176 238083 204232
rect 144913 204174 238083 204176
rect 144913 204171 144979 204174
rect 238017 204171 238083 204174
rect 227069 203690 227135 203693
rect 411253 203690 411319 203693
rect 227069 203688 411319 203690
rect 227069 203632 227074 203688
rect 227130 203632 411258 203688
rect 411314 203632 411319 203688
rect 227069 203630 411319 203632
rect 227069 203627 227135 203630
rect 411253 203627 411319 203630
rect 92381 203554 92447 203557
rect 209037 203554 209103 203557
rect 92381 203552 209103 203554
rect 92381 203496 92386 203552
rect 92442 203496 209042 203552
rect 209098 203496 209103 203552
rect 92381 203494 209103 203496
rect 92381 203491 92447 203494
rect 209037 203491 209103 203494
rect 210509 203554 210575 203557
rect 426433 203554 426499 203557
rect 210509 203552 426499 203554
rect 210509 203496 210514 203552
rect 210570 203496 426438 203552
rect 426494 203496 426499 203552
rect 210509 203494 426499 203496
rect 210509 203491 210575 203494
rect 426433 203491 426499 203494
rect 120073 202874 120139 202877
rect 156597 202874 156663 202877
rect 120073 202872 156663 202874
rect 120073 202816 120078 202872
rect 120134 202816 156602 202872
rect 156658 202816 156663 202872
rect 120073 202814 156663 202816
rect 120073 202811 120139 202814
rect 156597 202811 156663 202814
rect 177757 202876 177823 202877
rect 177757 202872 177804 202876
rect 177868 202874 177874 202876
rect 177757 202816 177762 202872
rect 177757 202812 177804 202816
rect 177868 202814 177914 202874
rect 177868 202812 177874 202814
rect 177757 202811 177823 202812
rect 91001 202330 91067 202333
rect 295926 202330 295932 202332
rect 91001 202328 295932 202330
rect 91001 202272 91006 202328
rect 91062 202272 295932 202328
rect 91001 202270 295932 202272
rect 91001 202267 91067 202270
rect 295926 202268 295932 202270
rect 295996 202268 296002 202332
rect 141417 202194 141483 202197
rect 191833 202194 191899 202197
rect 141417 202192 191899 202194
rect 141417 202136 141422 202192
rect 141478 202136 191838 202192
rect 191894 202136 191899 202192
rect 141417 202134 191899 202136
rect 141417 202131 141483 202134
rect 191833 202131 191899 202134
rect 195237 202194 195303 202197
rect 404997 202194 405063 202197
rect 195237 202192 405063 202194
rect 195237 202136 195242 202192
rect 195298 202136 405002 202192
rect 405058 202136 405063 202192
rect 195237 202134 405063 202136
rect 195237 202131 195303 202134
rect 404997 202131 405063 202134
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 216765 200970 216831 200973
rect 225689 200970 225755 200973
rect 216765 200968 225755 200970
rect 216765 200912 216770 200968
rect 216826 200912 225694 200968
rect 225750 200912 225755 200968
rect 216765 200910 225755 200912
rect 216765 200907 216831 200910
rect 225689 200907 225755 200910
rect 136541 200834 136607 200837
rect 316769 200834 316835 200837
rect 136541 200832 316835 200834
rect 136541 200776 136546 200832
rect 136602 200776 316774 200832
rect 316830 200776 316835 200832
rect 136541 200774 316835 200776
rect 136541 200771 136607 200774
rect 316769 200771 316835 200774
rect 81341 200698 81407 200701
rect 169017 200698 169083 200701
rect 81341 200696 169083 200698
rect 81341 200640 81346 200696
rect 81402 200640 169022 200696
rect 169078 200640 169083 200696
rect 81341 200638 169083 200640
rect 81341 200635 81407 200638
rect 169017 200635 169083 200638
rect 181621 200698 181687 200701
rect 369117 200698 369183 200701
rect 181621 200696 369183 200698
rect 181621 200640 181626 200696
rect 181682 200640 369122 200696
rect 369178 200640 369183 200696
rect 181621 200638 369183 200640
rect 181621 200635 181687 200638
rect 369117 200635 369183 200638
rect 121361 200018 121427 200021
rect 157926 200018 157932 200020
rect 121361 200016 157932 200018
rect 121361 199960 121366 200016
rect 121422 199960 157932 200016
rect 121361 199958 157932 199960
rect 121361 199955 121427 199958
rect 157926 199956 157932 199958
rect 157996 199956 158002 200020
rect 103421 199474 103487 199477
rect 195145 199474 195211 199477
rect 103421 199472 195211 199474
rect 103421 199416 103426 199472
rect 103482 199416 195150 199472
rect 195206 199416 195211 199472
rect 103421 199414 195211 199416
rect 103421 199411 103487 199414
rect 195145 199411 195211 199414
rect 216029 199474 216095 199477
rect 230606 199474 230612 199476
rect 216029 199472 230612 199474
rect 216029 199416 216034 199472
rect 216090 199416 230612 199472
rect 216029 199414 230612 199416
rect 216029 199411 216095 199414
rect 230606 199412 230612 199414
rect 230676 199412 230682 199476
rect 153101 199338 153167 199341
rect 309869 199338 309935 199341
rect 153101 199336 309935 199338
rect 153101 199280 153106 199336
rect 153162 199280 309874 199336
rect 309930 199280 309935 199336
rect 153101 199278 309935 199280
rect 153101 199275 153167 199278
rect 309869 199275 309935 199278
rect 195237 198794 195303 198797
rect 244222 198794 244228 198796
rect 195237 198792 244228 198794
rect 195237 198736 195242 198792
rect 195298 198736 244228 198792
rect 195237 198734 244228 198736
rect 195237 198731 195303 198734
rect 244222 198732 244228 198734
rect 244292 198732 244298 198796
rect 86861 198250 86927 198253
rect 177389 198250 177455 198253
rect 86861 198248 177455 198250
rect 86861 198192 86866 198248
rect 86922 198192 177394 198248
rect 177450 198192 177455 198248
rect 86861 198190 177455 198192
rect 86861 198187 86927 198190
rect 177389 198187 177455 198190
rect 119981 198114 120047 198117
rect 240726 198114 240732 198116
rect 119981 198112 240732 198114
rect 119981 198056 119986 198112
rect 120042 198056 240732 198112
rect 119981 198054 240732 198056
rect 119981 198051 120047 198054
rect 240726 198052 240732 198054
rect 240796 198052 240802 198116
rect 166901 197978 166967 197981
rect 429193 197978 429259 197981
rect 166901 197976 429259 197978
rect 166901 197920 166906 197976
rect 166962 197920 429198 197976
rect 429254 197920 429259 197976
rect 166901 197918 429259 197920
rect 166901 197915 166967 197918
rect 429193 197915 429259 197918
rect 191833 197298 191899 197301
rect 191833 197296 258090 197298
rect 191833 197240 191838 197296
rect 191894 197240 258090 197296
rect 191833 197238 258090 197240
rect 191833 197235 191899 197238
rect 113081 196754 113147 196757
rect 193857 196754 193923 196757
rect 113081 196752 193923 196754
rect 113081 196696 113086 196752
rect 113142 196696 193862 196752
rect 193918 196696 193923 196752
rect 113081 196694 193923 196696
rect 258030 196754 258090 197238
rect 260833 196754 260899 196757
rect 292665 196754 292731 196757
rect 258030 196752 292731 196754
rect 258030 196696 260838 196752
rect 260894 196696 292670 196752
rect 292726 196696 292731 196752
rect 258030 196694 292731 196696
rect 113081 196691 113147 196694
rect 193857 196691 193923 196694
rect 260833 196691 260899 196694
rect 292665 196691 292731 196694
rect 87597 196618 87663 196621
rect 583753 196618 583819 196621
rect 87597 196616 583819 196618
rect 87597 196560 87602 196616
rect 87658 196560 583758 196616
rect 583814 196560 583819 196616
rect 87597 196558 583819 196560
rect 87597 196555 87663 196558
rect 583753 196555 583819 196558
rect 117221 195938 117287 195941
rect 245694 195938 245700 195940
rect 117221 195936 245700 195938
rect 117221 195880 117226 195936
rect 117282 195880 245700 195936
rect 117221 195878 245700 195880
rect 117221 195875 117287 195878
rect 245694 195876 245700 195878
rect 245764 195876 245770 195940
rect 198365 195394 198431 195397
rect 278998 195394 279004 195396
rect 198365 195392 279004 195394
rect 198365 195336 198370 195392
rect 198426 195336 279004 195392
rect 198365 195334 279004 195336
rect 198365 195331 198431 195334
rect 278998 195332 279004 195334
rect 279068 195332 279074 195396
rect 72417 195258 72483 195261
rect 351177 195258 351243 195261
rect 72417 195256 351243 195258
rect 72417 195200 72422 195256
rect 72478 195200 351182 195256
rect 351238 195200 351243 195256
rect 72417 195198 351243 195200
rect 72417 195195 72483 195198
rect 351177 195195 351243 195198
rect 279417 194578 279483 194581
rect 284334 194578 284340 194580
rect 279417 194576 284340 194578
rect 279417 194520 279422 194576
rect 279478 194520 284340 194576
rect 279417 194518 284340 194520
rect 279417 194515 279483 194518
rect 284334 194516 284340 194518
rect 284404 194516 284410 194580
rect 90357 194170 90423 194173
rect 173157 194170 173223 194173
rect 90357 194168 173223 194170
rect 90357 194112 90362 194168
rect 90418 194112 173162 194168
rect 173218 194112 173223 194168
rect 90357 194110 173223 194112
rect 90357 194107 90423 194110
rect 173157 194107 173223 194110
rect 160829 194034 160895 194037
rect 280429 194034 280495 194037
rect 160829 194032 280495 194034
rect 160829 193976 160834 194032
rect 160890 193976 280434 194032
rect 280490 193976 280495 194032
rect 160829 193974 280495 193976
rect 160829 193971 160895 193974
rect 280429 193971 280495 193974
rect 104801 193898 104867 193901
rect 315297 193898 315363 193901
rect 104801 193896 315363 193898
rect 104801 193840 104806 193896
rect 104862 193840 315302 193896
rect 315358 193840 315363 193896
rect 104801 193838 315363 193840
rect 104801 193835 104867 193838
rect 315297 193835 315363 193838
rect 142061 193218 142127 193221
rect 378133 193218 378199 193221
rect 378869 193218 378935 193221
rect 142061 193216 378935 193218
rect 142061 193160 142066 193216
rect 142122 193160 378138 193216
rect 378194 193160 378874 193216
rect 378930 193160 378935 193216
rect 142061 193158 378935 193160
rect 142061 193155 142127 193158
rect 378133 193155 378199 193158
rect 378869 193155 378935 193158
rect 78673 193082 78739 193085
rect 284293 193082 284359 193085
rect 78673 193080 287070 193082
rect 78673 193024 78678 193080
rect 78734 193024 284298 193080
rect 284354 193024 287070 193080
rect 78673 193022 287070 193024
rect 78673 193019 78739 193022
rect 284293 193019 284359 193022
rect 287010 192674 287070 193022
rect 291142 192674 291148 192676
rect 287010 192614 291148 192674
rect 291142 192612 291148 192614
rect 291212 192612 291218 192676
rect 244222 192476 244228 192540
rect 244292 192538 244298 192540
rect 392669 192538 392735 192541
rect 244292 192536 392735 192538
rect 244292 192480 392674 192536
rect 392730 192480 392735 192536
rect 244292 192478 392735 192480
rect 244292 192476 244298 192478
rect 392669 192475 392735 192478
rect 583201 192538 583267 192541
rect 583520 192538 584960 192628
rect 583201 192536 584960 192538
rect 583201 192480 583206 192536
rect 583262 192480 584960 192536
rect 583201 192478 584960 192480
rect 583201 192475 583267 192478
rect 583520 192388 584960 192478
rect 29637 191722 29703 191725
rect 30281 191722 30347 191725
rect 29637 191720 30347 191722
rect 29637 191664 29642 191720
rect 29698 191664 30286 191720
rect 30342 191664 30347 191720
rect 29637 191662 30347 191664
rect 29637 191659 29703 191662
rect 30281 191659 30347 191662
rect 184657 191178 184723 191181
rect 245694 191178 245700 191180
rect 184657 191176 245700 191178
rect 184657 191120 184662 191176
rect 184718 191120 245700 191176
rect 184657 191118 245700 191120
rect 184657 191115 184723 191118
rect 245694 191116 245700 191118
rect 245764 191116 245770 191180
rect 107561 191042 107627 191045
rect 287646 191042 287652 191044
rect 107561 191040 287652 191042
rect 107561 190984 107566 191040
rect 107622 190984 287652 191040
rect 107561 190982 287652 190984
rect 107561 190979 107627 190982
rect 287646 190980 287652 190982
rect 287716 190980 287722 191044
rect 29637 190498 29703 190501
rect 374729 190498 374795 190501
rect 29637 190496 374795 190498
rect 29637 190440 29642 190496
rect 29698 190440 374734 190496
rect 374790 190440 374795 190496
rect 29637 190438 374795 190440
rect 29637 190435 29703 190438
rect 374729 190435 374795 190438
rect 17861 190362 17927 190365
rect 162117 190362 162183 190365
rect 17861 190360 162183 190362
rect 17861 190304 17866 190360
rect 17922 190304 162122 190360
rect 162178 190304 162183 190360
rect 17861 190302 162183 190304
rect 17861 190299 17927 190302
rect 162117 190299 162183 190302
rect 200614 189892 200620 189956
rect 200684 189954 200690 189956
rect 278313 189954 278379 189957
rect 200684 189952 278379 189954
rect 200684 189896 278318 189952
rect 278374 189896 278379 189952
rect 200684 189894 278379 189896
rect 200684 189892 200690 189894
rect 278313 189891 278379 189894
rect 154481 189818 154547 189821
rect 316677 189818 316743 189821
rect 154481 189816 316743 189818
rect 154481 189760 154486 189816
rect 154542 189760 316682 189816
rect 316738 189760 316743 189816
rect 154481 189758 316743 189760
rect 154481 189755 154547 189758
rect 316677 189755 316743 189758
rect 96521 189682 96587 189685
rect 449985 189682 450051 189685
rect 96521 189680 450051 189682
rect 96521 189624 96526 189680
rect 96582 189624 449990 189680
rect 450046 189624 450051 189680
rect 96521 189622 450051 189624
rect 96521 189619 96587 189622
rect 449985 189619 450051 189622
rect 17217 189138 17283 189141
rect 17861 189138 17927 189141
rect 17217 189136 17927 189138
rect 17217 189080 17222 189136
rect 17278 189080 17866 189136
rect 17922 189080 17927 189136
rect 17217 189078 17927 189080
rect 17217 189075 17283 189078
rect 17861 189075 17927 189078
rect -960 188866 480 188956
rect 2773 188866 2839 188869
rect -960 188864 2839 188866
rect -960 188808 2778 188864
rect 2834 188808 2839 188864
rect -960 188806 2839 188808
rect -960 188716 480 188806
rect 2773 188803 2839 188806
rect 161381 188458 161447 188461
rect 187049 188458 187115 188461
rect 161381 188456 187115 188458
rect 161381 188400 161386 188456
rect 161442 188400 187054 188456
rect 187110 188400 187115 188456
rect 161381 188398 187115 188400
rect 161381 188395 161447 188398
rect 187049 188395 187115 188398
rect 188337 188458 188403 188461
rect 301037 188458 301103 188461
rect 188337 188456 301103 188458
rect 188337 188400 188342 188456
rect 188398 188400 301042 188456
rect 301098 188400 301103 188456
rect 188337 188398 301103 188400
rect 188337 188395 188403 188398
rect 301037 188395 301103 188398
rect 75678 188260 75684 188324
rect 75748 188322 75754 188324
rect 443085 188322 443151 188325
rect 75748 188320 443151 188322
rect 75748 188264 443090 188320
rect 443146 188264 443151 188320
rect 75748 188262 443151 188264
rect 75748 188260 75754 188262
rect 443085 188259 443151 188262
rect 218789 187778 218855 187781
rect 248505 187778 248571 187781
rect 218789 187776 248571 187778
rect 218789 187720 218794 187776
rect 218850 187720 248510 187776
rect 248566 187720 248571 187776
rect 218789 187718 248571 187720
rect 218789 187715 218855 187718
rect 248505 187715 248571 187718
rect 163589 187234 163655 187237
rect 207013 187234 207079 187237
rect 163589 187232 207079 187234
rect 163589 187176 163594 187232
rect 163650 187176 207018 187232
rect 207074 187176 207079 187232
rect 163589 187174 207079 187176
rect 163589 187171 163655 187174
rect 207013 187171 207079 187174
rect 151077 187098 151143 187101
rect 305494 187098 305500 187100
rect 151077 187096 305500 187098
rect 151077 187040 151082 187096
rect 151138 187040 305500 187096
rect 151077 187038 305500 187040
rect 151077 187035 151143 187038
rect 305494 187036 305500 187038
rect 305564 187036 305570 187100
rect 95141 186962 95207 186965
rect 299606 186962 299612 186964
rect 95141 186960 299612 186962
rect 95141 186904 95146 186960
rect 95202 186904 299612 186960
rect 95141 186902 299612 186904
rect 95141 186899 95207 186902
rect 299606 186900 299612 186902
rect 299676 186900 299682 186964
rect 269757 186418 269823 186421
rect 277158 186418 277164 186420
rect 269757 186416 277164 186418
rect 269757 186360 269762 186416
rect 269818 186360 277164 186416
rect 269757 186358 277164 186360
rect 269757 186355 269823 186358
rect 277158 186356 277164 186358
rect 277228 186356 277234 186420
rect 278037 186418 278103 186421
rect 285622 186418 285628 186420
rect 278037 186416 285628 186418
rect 278037 186360 278042 186416
rect 278098 186360 285628 186416
rect 278037 186358 285628 186360
rect 278037 186355 278103 186358
rect 285622 186356 285628 186358
rect 285692 186356 285698 186420
rect 54845 186282 54911 186285
rect 197997 186282 198063 186285
rect 54845 186280 198063 186282
rect 54845 186224 54850 186280
rect 54906 186224 198002 186280
rect 198058 186224 198063 186280
rect 54845 186222 198063 186224
rect 54845 186219 54911 186222
rect 197997 186219 198063 186222
rect 217317 185874 217383 185877
rect 227662 185874 227668 185876
rect 217317 185872 227668 185874
rect 217317 185816 217322 185872
rect 217378 185816 227668 185872
rect 217317 185814 227668 185816
rect 217317 185811 217383 185814
rect 227662 185812 227668 185814
rect 227732 185812 227738 185876
rect 211797 185738 211863 185741
rect 237414 185738 237420 185740
rect 211797 185736 237420 185738
rect 211797 185680 211802 185736
rect 211858 185680 237420 185736
rect 211797 185678 237420 185680
rect 211797 185675 211863 185678
rect 237414 185676 237420 185678
rect 237484 185676 237490 185740
rect 278129 185738 278195 185741
rect 281758 185738 281764 185740
rect 278129 185736 281764 185738
rect 278129 185680 278134 185736
rect 278190 185680 281764 185736
rect 278129 185678 281764 185680
rect 278129 185675 278195 185678
rect 281758 185676 281764 185678
rect 281828 185676 281834 185740
rect 170857 185602 170923 185605
rect 188838 185602 188844 185604
rect 170857 185600 188844 185602
rect 170857 185544 170862 185600
rect 170918 185544 188844 185600
rect 170857 185542 188844 185544
rect 170857 185539 170923 185542
rect 188838 185540 188844 185542
rect 188908 185602 188914 185604
rect 202229 185602 202295 185605
rect 295333 185602 295399 185605
rect 188908 185542 190470 185602
rect 188908 185540 188914 185542
rect 106181 185194 106247 185197
rect 167637 185194 167703 185197
rect 106181 185192 167703 185194
rect 106181 185136 106186 185192
rect 106242 185136 167642 185192
rect 167698 185136 167703 185192
rect 106181 185134 167703 185136
rect 106181 185131 106247 185134
rect 167637 185131 167703 185134
rect 100661 185058 100727 185061
rect 180149 185058 180215 185061
rect 100661 185056 180215 185058
rect 100661 185000 100666 185056
rect 100722 185000 180154 185056
rect 180210 185000 180215 185056
rect 100661 184998 180215 185000
rect 190410 185058 190470 185542
rect 202229 185600 295399 185602
rect 202229 185544 202234 185600
rect 202290 185544 295338 185600
rect 295394 185544 295399 185600
rect 202229 185542 295399 185544
rect 202229 185539 202295 185542
rect 295333 185539 295399 185542
rect 249885 185468 249951 185469
rect 249885 185466 249932 185468
rect 249840 185464 249932 185466
rect 249840 185408 249890 185464
rect 249840 185406 249932 185408
rect 249885 185404 249932 185406
rect 249996 185404 250002 185468
rect 249885 185403 249951 185404
rect 215293 185058 215359 185061
rect 190410 185056 215359 185058
rect 190410 185000 215298 185056
rect 215354 185000 215359 185056
rect 190410 184998 215359 185000
rect 100661 184995 100727 184998
rect 180149 184995 180215 184998
rect 215293 184995 215359 184998
rect 227805 185058 227871 185061
rect 398598 185058 398604 185060
rect 227805 185056 398604 185058
rect 227805 185000 227810 185056
rect 227866 185000 398604 185056
rect 227805 184998 398604 185000
rect 227805 184995 227871 184998
rect 398598 184996 398604 184998
rect 398668 184996 398674 185060
rect 225689 184514 225755 184517
rect 270309 184514 270375 184517
rect 225689 184512 270375 184514
rect 225689 184456 225694 184512
rect 225750 184456 270314 184512
rect 270370 184456 270375 184512
rect 225689 184454 270375 184456
rect 225689 184451 225755 184454
rect 270309 184451 270375 184454
rect 162158 184316 162164 184380
rect 162228 184378 162234 184380
rect 334709 184378 334775 184381
rect 162228 184376 334775 184378
rect 162228 184320 334714 184376
rect 334770 184320 334775 184376
rect 162228 184318 334775 184320
rect 162228 184316 162234 184318
rect 334709 184315 334775 184318
rect 117129 184242 117195 184245
rect 293217 184242 293283 184245
rect 117129 184240 293283 184242
rect 117129 184184 117134 184240
rect 117190 184184 293222 184240
rect 293278 184184 293283 184240
rect 117129 184182 293283 184184
rect 117129 184179 117195 184182
rect 293217 184179 293283 184182
rect 102041 183698 102107 183701
rect 169109 183698 169175 183701
rect 102041 183696 169175 183698
rect 102041 183640 102046 183696
rect 102102 183640 169114 183696
rect 169170 183640 169175 183696
rect 102041 183638 169175 183640
rect 102041 183635 102107 183638
rect 169109 183635 169175 183638
rect 131021 183154 131087 183157
rect 288566 183154 288572 183156
rect 131021 183152 288572 183154
rect 131021 183096 131026 183152
rect 131082 183096 288572 183152
rect 131021 183094 288572 183096
rect 131021 183091 131087 183094
rect 288566 183092 288572 183094
rect 288636 183092 288642 183156
rect 159950 182956 159956 183020
rect 160020 183018 160026 183020
rect 393405 183018 393471 183021
rect 160020 183016 393471 183018
rect 160020 182960 393410 183016
rect 393466 182960 393471 183016
rect 160020 182958 393471 182960
rect 160020 182956 160026 182958
rect 393405 182955 393471 182958
rect 186221 182882 186287 182885
rect 445937 182882 446003 182885
rect 186221 182880 446003 182882
rect 186221 182824 186226 182880
rect 186282 182824 445942 182880
rect 445998 182824 446003 182880
rect 186221 182822 446003 182824
rect 186221 182819 186287 182822
rect 445937 182819 446003 182822
rect 98821 182202 98887 182205
rect 178861 182202 178927 182205
rect 98821 182200 178927 182202
rect 98821 182144 98826 182200
rect 98882 182144 178866 182200
rect 178922 182144 178927 182200
rect 98821 182142 178927 182144
rect 98821 182139 98887 182142
rect 178861 182139 178927 182142
rect 93761 182066 93827 182069
rect 175089 182066 175155 182069
rect 93761 182064 175155 182066
rect 93761 182008 93766 182064
rect 93822 182008 175094 182064
rect 175150 182008 175155 182064
rect 93761 182006 175155 182008
rect 93761 182003 93827 182006
rect 175089 182003 175155 182006
rect 206553 181658 206619 181661
rect 237598 181658 237604 181660
rect 206553 181656 237604 181658
rect 206553 181600 206558 181656
rect 206614 181600 237604 181656
rect 206553 181598 237604 181600
rect 206553 181595 206619 181598
rect 237598 181596 237604 181598
rect 237668 181596 237674 181660
rect 155861 181522 155927 181525
rect 298686 181522 298692 181524
rect 155861 181520 298692 181522
rect 155861 181464 155866 181520
rect 155922 181464 298692 181520
rect 155861 181462 298692 181464
rect 155861 181459 155927 181462
rect 298686 181460 298692 181462
rect 298756 181460 298762 181524
rect 175089 181386 175155 181389
rect 400305 181386 400371 181389
rect 175089 181384 400371 181386
rect 175089 181328 175094 181384
rect 175150 181328 400310 181384
rect 400366 181328 400371 181384
rect 175089 181326 400371 181328
rect 175089 181323 175155 181326
rect 400305 181323 400371 181326
rect 108113 180842 108179 180845
rect 173341 180842 173407 180845
rect 108113 180840 173407 180842
rect 108113 180784 108118 180840
rect 108174 180784 173346 180840
rect 173402 180784 173407 180840
rect 108113 180782 173407 180784
rect 108113 180779 108179 180782
rect 173341 180779 173407 180782
rect 227069 180298 227135 180301
rect 238845 180298 238911 180301
rect 227069 180296 238911 180298
rect 227069 180240 227074 180296
rect 227130 180240 238850 180296
rect 238906 180240 238911 180296
rect 227069 180238 238911 180240
rect 227069 180235 227135 180238
rect 238845 180235 238911 180238
rect 197169 180162 197235 180165
rect 226333 180162 226399 180165
rect 197169 180160 226399 180162
rect 197169 180104 197174 180160
rect 197230 180104 226338 180160
rect 226394 180104 226399 180160
rect 197169 180102 226399 180104
rect 197169 180099 197235 180102
rect 226333 180099 226399 180102
rect 274081 180162 274147 180165
rect 290590 180162 290596 180164
rect 274081 180160 290596 180162
rect 274081 180104 274086 180160
rect 274142 180104 290596 180160
rect 274081 180102 290596 180104
rect 274081 180099 274147 180102
rect 290590 180100 290596 180102
rect 290660 180100 290666 180164
rect 166257 180026 166323 180029
rect 441705 180026 441771 180029
rect 166257 180024 441771 180026
rect 166257 179968 166262 180024
rect 166318 179968 441710 180024
rect 441766 179968 441771 180024
rect 166257 179966 441771 179968
rect 166257 179963 166323 179966
rect 441705 179963 441771 179966
rect 110689 179618 110755 179621
rect 166441 179618 166507 179621
rect 110689 179616 166507 179618
rect 110689 179560 110694 179616
rect 110750 179560 166446 179616
rect 166502 179560 166507 179616
rect 110689 179558 166507 179560
rect 110689 179555 110755 179558
rect 166441 179555 166507 179558
rect 97257 179482 97323 179485
rect 170397 179482 170463 179485
rect 97257 179480 170463 179482
rect 97257 179424 97262 179480
rect 97318 179424 170402 179480
rect 170458 179424 170463 179480
rect 97257 179422 170463 179424
rect 97257 179419 97323 179422
rect 170397 179419 170463 179422
rect 216765 179482 216831 179485
rect 255405 179482 255471 179485
rect 216765 179480 255471 179482
rect 216765 179424 216770 179480
rect 216826 179424 255410 179480
rect 255466 179424 255471 179480
rect 216765 179422 255471 179424
rect 216765 179419 216831 179422
rect 255405 179419 255471 179422
rect 148961 179346 149027 179349
rect 230381 179346 230447 179349
rect 148961 179344 230447 179346
rect 148961 179288 148966 179344
rect 149022 179288 230386 179344
rect 230442 179288 230447 179344
rect 148961 179286 230447 179288
rect 148961 179283 149027 179286
rect 230381 179283 230447 179286
rect 583520 179210 584960 179300
rect 583342 179150 584960 179210
rect 583342 179074 583402 179150
rect 583520 179074 584960 179150
rect 583342 179060 584960 179074
rect 583342 179014 583586 179060
rect 180006 178740 180012 178804
rect 180076 178802 180082 178804
rect 196617 178802 196683 178805
rect 180076 178800 196683 178802
rect 180076 178744 196622 178800
rect 196678 178744 196683 178800
rect 180076 178742 196683 178744
rect 180076 178740 180082 178742
rect 196617 178739 196683 178742
rect 276657 178802 276723 178805
rect 279969 178802 280035 178805
rect 276657 178800 280035 178802
rect 276657 178744 276662 178800
rect 276718 178744 279974 178800
rect 280030 178744 280035 178800
rect 276657 178742 280035 178744
rect 276657 178739 276723 178742
rect 279969 178739 280035 178742
rect 583526 178669 583586 179014
rect 193121 178666 193187 178669
rect 245653 178666 245719 178669
rect 193121 178664 245719 178666
rect 193121 178608 193126 178664
rect 193182 178608 245658 178664
rect 245714 178608 245719 178664
rect 193121 178606 245719 178608
rect 193121 178603 193187 178606
rect 245653 178603 245719 178606
rect 259269 178666 259335 178669
rect 274633 178666 274699 178669
rect 259269 178664 274699 178666
rect 259269 178608 259274 178664
rect 259330 178608 274638 178664
rect 274694 178608 274699 178664
rect 259269 178606 274699 178608
rect 259269 178603 259335 178606
rect 274633 178603 274699 178606
rect 278313 178666 278379 178669
rect 291469 178666 291535 178669
rect 278313 178664 291535 178666
rect 278313 178608 278318 178664
rect 278374 178608 291474 178664
rect 291530 178608 291535 178664
rect 278313 178606 291535 178608
rect 278313 178603 278379 178606
rect 291469 178603 291535 178606
rect 583477 178664 583586 178669
rect 583477 178608 583482 178664
rect 583538 178608 583586 178664
rect 583477 178606 583586 178608
rect 583477 178603 583543 178606
rect 231761 178258 231827 178261
rect 233366 178258 233372 178260
rect 231761 178256 233372 178258
rect 231761 178200 231766 178256
rect 231822 178200 233372 178256
rect 231761 178198 233372 178200
rect 231761 178195 231827 178198
rect 233366 178196 233372 178198
rect 233436 178196 233442 178260
rect 176101 178122 176167 178125
rect 113130 178120 176167 178122
rect 113130 178064 176106 178120
rect 176162 178064 176167 178120
rect 113130 178062 176167 178064
rect 112110 177924 112116 177988
rect 112180 177986 112186 177988
rect 113130 177986 113190 178062
rect 176101 178059 176167 178062
rect 216673 178122 216739 178125
rect 240777 178122 240843 178125
rect 216673 178120 240843 178122
rect 216673 178064 216678 178120
rect 216734 178064 240782 178120
rect 240838 178064 240843 178120
rect 216673 178062 240843 178064
rect 216673 178059 216739 178062
rect 240777 178059 240843 178062
rect 275277 178122 275343 178125
rect 278814 178122 278820 178124
rect 275277 178120 278820 178122
rect 275277 178064 275282 178120
rect 275338 178064 278820 178120
rect 275277 178062 278820 178064
rect 275277 178059 275343 178062
rect 278814 178060 278820 178062
rect 278884 178060 278890 178124
rect 279601 178122 279667 178125
rect 280470 178122 280476 178124
rect 279601 178120 280476 178122
rect 279601 178064 279606 178120
rect 279662 178064 280476 178120
rect 279601 178062 280476 178064
rect 279601 178059 279667 178062
rect 280470 178060 280476 178062
rect 280540 178060 280546 178124
rect 112180 177926 113190 177986
rect 284293 177986 284359 177989
rect 284518 177986 284524 177988
rect 284293 177984 284524 177986
rect 284293 177928 284298 177984
rect 284354 177928 284524 177984
rect 284293 177926 284524 177928
rect 112180 177924 112186 177926
rect 284293 177923 284359 177926
rect 284518 177924 284524 177926
rect 284588 177924 284594 177988
rect 98310 177516 98316 177580
rect 98380 177578 98386 177580
rect 98821 177578 98887 177581
rect 98380 177576 98887 177578
rect 98380 177520 98826 177576
rect 98882 177520 98887 177576
rect 98380 177518 98887 177520
rect 98380 177516 98386 177518
rect 98821 177515 98887 177518
rect 100702 177516 100708 177580
rect 100772 177578 100778 177580
rect 102041 177578 102107 177581
rect 100772 177576 102107 177578
rect 100772 177520 102046 177576
rect 102102 177520 102107 177576
rect 100772 177518 102107 177520
rect 100772 177516 100778 177518
rect 102041 177515 102107 177518
rect 105670 177516 105676 177580
rect 105740 177578 105746 177580
rect 106181 177578 106247 177581
rect 108113 177580 108179 177581
rect 108062 177578 108068 177580
rect 105740 177576 106247 177578
rect 105740 177520 106186 177576
rect 106242 177520 106247 177576
rect 105740 177518 106247 177520
rect 108022 177518 108068 177578
rect 108132 177576 108179 177580
rect 108174 177520 108179 177576
rect 105740 177516 105746 177518
rect 106181 177515 106247 177518
rect 108062 177516 108068 177518
rect 108132 177516 108179 177520
rect 109534 177516 109540 177580
rect 109604 177578 109610 177580
rect 110321 177578 110387 177581
rect 114369 177580 114435 177581
rect 114318 177578 114324 177580
rect 109604 177576 110387 177578
rect 109604 177520 110326 177576
rect 110382 177520 110387 177576
rect 109604 177518 110387 177520
rect 114278 177518 114324 177578
rect 114388 177576 114435 177580
rect 114430 177520 114435 177576
rect 109604 177516 109610 177518
rect 108113 177515 108179 177516
rect 110321 177515 110387 177518
rect 114318 177516 114324 177518
rect 114388 177516 114435 177520
rect 121862 177516 121868 177580
rect 121932 177578 121938 177580
rect 122741 177578 122807 177581
rect 121932 177576 122807 177578
rect 121932 177520 122746 177576
rect 122802 177520 122807 177576
rect 121932 177518 122807 177520
rect 121932 177516 121938 177518
rect 114369 177515 114435 177516
rect 122741 177515 122807 177518
rect 123150 177516 123156 177580
rect 123220 177578 123226 177580
rect 124029 177578 124095 177581
rect 123220 177576 124095 177578
rect 123220 177520 124034 177576
rect 124090 177520 124095 177576
rect 123220 177518 124095 177520
rect 123220 177516 123226 177518
rect 124029 177515 124095 177518
rect 124438 177516 124444 177580
rect 124508 177578 124514 177580
rect 125501 177578 125567 177581
rect 124508 177576 125567 177578
rect 124508 177520 125506 177576
rect 125562 177520 125567 177576
rect 124508 177518 125567 177520
rect 124508 177516 124514 177518
rect 125501 177515 125567 177518
rect 125726 177516 125732 177580
rect 125796 177578 125802 177580
rect 126881 177578 126947 177581
rect 125796 177576 126947 177578
rect 125796 177520 126886 177576
rect 126942 177520 126947 177576
rect 125796 177518 126947 177520
rect 125796 177516 125802 177518
rect 126881 177515 126947 177518
rect 130694 177516 130700 177580
rect 130764 177578 130770 177580
rect 130929 177578 130995 177581
rect 132401 177580 132467 177581
rect 132350 177578 132356 177580
rect 130764 177576 130995 177578
rect 130764 177520 130934 177576
rect 130990 177520 130995 177576
rect 130764 177518 130995 177520
rect 132310 177518 132356 177578
rect 132420 177576 132467 177580
rect 132462 177520 132467 177576
rect 130764 177516 130770 177518
rect 130929 177515 130995 177518
rect 132350 177516 132356 177518
rect 132420 177516 132467 177520
rect 133086 177516 133092 177580
rect 133156 177578 133162 177580
rect 133781 177578 133847 177581
rect 133156 177576 133847 177578
rect 133156 177520 133786 177576
rect 133842 177520 133847 177576
rect 133156 177518 133847 177520
rect 133156 177516 133162 177518
rect 132401 177515 132467 177516
rect 133781 177515 133847 177518
rect 148174 177516 148180 177580
rect 148244 177578 148250 177580
rect 148869 177578 148935 177581
rect 148244 177576 148935 177578
rect 148244 177520 148874 177576
rect 148930 177520 148935 177576
rect 148244 177518 148935 177520
rect 148244 177516 148250 177518
rect 148869 177515 148935 177518
rect 216029 177578 216095 177581
rect 236085 177578 236151 177581
rect 216029 177576 236151 177578
rect 216029 177520 216034 177576
rect 216090 177520 236090 177576
rect 236146 177520 236151 177576
rect 216029 177518 236151 177520
rect 216029 177515 216095 177518
rect 236085 177515 236151 177518
rect 272517 177578 272583 177581
rect 287329 177578 287395 177581
rect 272517 177576 287395 177578
rect 272517 177520 272522 177576
rect 272578 177520 287334 177576
rect 287390 177520 287395 177576
rect 272517 177518 287395 177520
rect 272517 177515 272583 177518
rect 287329 177515 287395 177518
rect 118366 177380 118372 177444
rect 118436 177442 118442 177444
rect 118601 177442 118667 177445
rect 118436 177440 118667 177442
rect 118436 177384 118606 177440
rect 118662 177384 118667 177440
rect 118436 177382 118667 177384
rect 118436 177380 118442 177382
rect 118601 177379 118667 177382
rect 207749 177442 207815 177445
rect 284661 177442 284727 177445
rect 207749 177440 284727 177442
rect 207749 177384 207754 177440
rect 207810 177384 284666 177440
rect 284722 177384 284727 177440
rect 207749 177382 284727 177384
rect 207749 177379 207815 177382
rect 284661 177379 284727 177382
rect 104566 177244 104572 177308
rect 104636 177306 104642 177308
rect 177573 177306 177639 177309
rect 229461 177306 229527 177309
rect 104636 177246 113190 177306
rect 104636 177244 104642 177246
rect 110689 177172 110755 177173
rect 110638 177170 110644 177172
rect 110598 177110 110644 177170
rect 110708 177168 110755 177172
rect 110750 177112 110755 177168
rect 110638 177108 110644 177110
rect 110708 177108 110755 177112
rect 113130 177170 113190 177246
rect 177573 177304 229527 177306
rect 177573 177248 177578 177304
rect 177634 177248 229466 177304
rect 229522 177248 229527 177304
rect 177573 177246 229527 177248
rect 177573 177243 177639 177246
rect 229461 177243 229527 177246
rect 274633 177306 274699 177309
rect 445845 177306 445911 177309
rect 274633 177304 445911 177306
rect 274633 177248 274638 177304
rect 274694 177248 445850 177304
rect 445906 177248 445911 177304
rect 274633 177246 445911 177248
rect 274633 177243 274699 177246
rect 445845 177243 445911 177246
rect 214557 177170 214623 177173
rect 113130 177168 214623 177170
rect 113130 177112 214562 177168
rect 214618 177112 214623 177168
rect 113130 177110 214623 177112
rect 110689 177107 110755 177108
rect 214557 177107 214623 177110
rect 106958 176972 106964 177036
rect 107028 177034 107034 177036
rect 164550 177034 164556 177036
rect 107028 176974 164556 177034
rect 107028 176972 107034 176974
rect 164550 176972 164556 176974
rect 164620 176972 164626 177036
rect 97022 176836 97028 176900
rect 97092 176898 97098 176900
rect 97257 176898 97323 176901
rect 97092 176896 97323 176898
rect 97092 176840 97262 176896
rect 97318 176840 97323 176896
rect 97092 176838 97323 176840
rect 97092 176836 97098 176838
rect 97257 176835 97323 176838
rect 101990 176836 101996 176900
rect 102060 176898 102066 176900
rect 180241 176898 180307 176901
rect 102060 176896 180307 176898
rect 102060 176840 180246 176896
rect 180302 176840 180307 176896
rect 102060 176838 180307 176840
rect 102060 176836 102066 176838
rect 180241 176835 180307 176838
rect 100661 176762 100727 176765
rect 103329 176762 103395 176765
rect 99422 176760 100727 176762
rect 99422 176704 100666 176760
rect 100722 176704 100727 176760
rect 99422 176702 100727 176704
rect 99422 176492 99482 176702
rect 100661 176699 100727 176702
rect 103286 176760 103395 176762
rect 103286 176704 103334 176760
rect 103390 176704 103395 176760
rect 103286 176699 103395 176704
rect 113214 176700 113220 176764
rect 113284 176762 113290 176764
rect 113725 176762 113791 176765
rect 115841 176764 115907 176765
rect 119521 176764 119587 176765
rect 120809 176764 120875 176765
rect 127065 176764 127131 176765
rect 129457 176764 129523 176765
rect 115790 176762 115796 176764
rect 113284 176760 113791 176762
rect 113284 176704 113730 176760
rect 113786 176704 113791 176760
rect 113284 176702 113791 176704
rect 115750 176702 115796 176762
rect 115860 176760 115907 176764
rect 119470 176762 119476 176764
rect 115902 176704 115907 176760
rect 113284 176700 113290 176702
rect 113725 176699 113791 176702
rect 115790 176700 115796 176702
rect 115860 176700 115907 176704
rect 119430 176702 119476 176762
rect 119540 176760 119587 176764
rect 120758 176762 120764 176764
rect 119582 176704 119587 176760
rect 119470 176700 119476 176702
rect 119540 176700 119587 176704
rect 120718 176702 120764 176762
rect 120828 176760 120875 176764
rect 127014 176762 127020 176764
rect 120870 176704 120875 176760
rect 120758 176700 120764 176702
rect 120828 176700 120875 176704
rect 126974 176702 127020 176762
rect 127084 176760 127131 176764
rect 129406 176762 129412 176764
rect 127126 176704 127131 176760
rect 127014 176700 127020 176702
rect 127084 176700 127131 176704
rect 129366 176702 129412 176762
rect 129476 176760 129523 176764
rect 129518 176704 129523 176760
rect 129406 176700 129412 176702
rect 129476 176700 129523 176704
rect 158846 176700 158852 176764
rect 158916 176762 158922 176764
rect 158989 176762 159055 176765
rect 158916 176760 159055 176762
rect 158916 176704 158994 176760
rect 159050 176704 159055 176760
rect 158916 176702 159055 176704
rect 158916 176700 158922 176702
rect 115841 176699 115907 176700
rect 119521 176699 119587 176700
rect 120809 176699 120875 176700
rect 127065 176699 127131 176700
rect 129457 176699 129523 176700
rect 158989 176699 159055 176702
rect 226241 176762 226307 176765
rect 229134 176762 229140 176764
rect 226241 176760 229140 176762
rect 226241 176704 226246 176760
rect 226302 176704 229140 176760
rect 226241 176702 229140 176704
rect 226241 176699 226307 176702
rect 229134 176700 229140 176702
rect 229204 176700 229210 176764
rect 103286 176492 103346 176699
rect 163497 176626 163563 176629
rect 216673 176626 216739 176629
rect 163497 176624 216739 176626
rect 163497 176568 163502 176624
rect 163558 176568 216678 176624
rect 216734 176568 216739 176624
rect 163497 176566 216739 176568
rect 163497 176563 163563 176566
rect 216673 176563 216739 176566
rect 226926 176564 226932 176628
rect 226996 176626 227002 176628
rect 230013 176626 230079 176629
rect 226996 176624 230079 176626
rect 226996 176568 230018 176624
rect 230074 176568 230079 176624
rect 226996 176566 230079 176568
rect 226996 176564 227002 176566
rect 230013 176563 230079 176566
rect 99414 176428 99420 176492
rect 99484 176428 99490 176492
rect 103278 176428 103284 176492
rect 103348 176428 103354 176492
rect 227662 176428 227668 176492
rect 227732 176490 227738 176492
rect 229185 176490 229251 176493
rect 227732 176488 229251 176490
rect 227732 176432 229190 176488
rect 229246 176432 229251 176488
rect 227732 176430 229251 176432
rect 227732 176428 227738 176430
rect 229185 176427 229251 176430
rect 228214 176292 228220 176356
rect 228284 176354 228290 176356
rect 229369 176354 229435 176357
rect 228284 176352 229435 176354
rect 228284 176296 229374 176352
rect 229430 176296 229435 176352
rect 228284 176294 229435 176296
rect 228284 176292 228290 176294
rect 229369 176291 229435 176294
rect 227713 176218 227779 176221
rect 227713 176216 228282 176218
rect 227713 176160 227718 176216
rect 227774 176160 228282 176216
rect 227713 176158 228282 176160
rect 227713 176155 227779 176158
rect -960 175796 480 176036
rect 215477 175946 215543 175949
rect 226241 175946 226307 175949
rect 215477 175944 226307 175946
rect 215477 175888 215482 175944
rect 215538 175888 226246 175944
rect 226302 175888 226307 175944
rect 215477 175886 226307 175888
rect 215477 175883 215543 175886
rect 226241 175883 226307 175886
rect 128118 175612 128124 175676
rect 128188 175674 128194 175676
rect 213913 175674 213979 175677
rect 128188 175614 200130 175674
rect 128188 175612 128194 175614
rect 116894 175476 116900 175540
rect 116964 175538 116970 175540
rect 167729 175538 167795 175541
rect 116964 175536 167795 175538
rect 116964 175480 167734 175536
rect 167790 175480 167795 175536
rect 116964 175478 167795 175480
rect 200070 175538 200130 175614
rect 213913 175672 217028 175674
rect 213913 175616 213918 175672
rect 213974 175616 217028 175672
rect 228222 175644 228282 176158
rect 229001 175946 229067 175949
rect 229001 175944 229110 175946
rect 229001 175888 229006 175944
rect 229062 175888 229110 175944
rect 229001 175883 229110 175888
rect 229050 175810 229110 175883
rect 244222 175810 244228 175812
rect 229050 175750 244228 175810
rect 244222 175748 244228 175750
rect 244292 175748 244298 175812
rect 277342 175748 277348 175812
rect 277412 175810 277418 175812
rect 279417 175810 279483 175813
rect 277412 175808 279483 175810
rect 277412 175752 279422 175808
rect 279478 175752 279483 175808
rect 277412 175750 279483 175752
rect 277412 175748 277418 175750
rect 279417 175747 279483 175750
rect 264973 175674 265039 175677
rect 264973 175672 268180 175674
rect 213913 175614 217028 175616
rect 264973 175616 264978 175672
rect 265034 175616 268180 175672
rect 264973 175614 268180 175616
rect 213913 175611 213979 175614
rect 264973 175611 265039 175614
rect 214097 175538 214163 175541
rect 281533 175538 281599 175541
rect 200070 175536 214163 175538
rect 200070 175480 214102 175536
rect 214158 175480 214163 175536
rect 200070 175478 214163 175480
rect 279956 175536 281599 175538
rect 279956 175480 281538 175536
rect 281594 175480 281599 175536
rect 279956 175478 281599 175480
rect 116964 175476 116970 175478
rect 167729 175475 167795 175478
rect 214097 175475 214163 175478
rect 281533 175475 281599 175478
rect 134425 175404 134491 175405
rect 135713 175404 135779 175405
rect 134374 175402 134380 175404
rect 134334 175342 134380 175402
rect 134444 175400 134491 175404
rect 135662 175402 135668 175404
rect 134486 175344 134491 175400
rect 134374 175340 134380 175342
rect 134444 175340 134491 175344
rect 135622 175342 135668 175402
rect 135732 175400 135779 175404
rect 135774 175344 135779 175400
rect 135662 175340 135668 175342
rect 135732 175340 135779 175344
rect 134425 175339 134491 175340
rect 135713 175339 135779 175340
rect 229093 175266 229159 175269
rect 228988 175264 229159 175266
rect 228988 175208 229098 175264
rect 229154 175208 229159 175264
rect 228988 175206 229159 175208
rect 229093 175203 229159 175206
rect 265065 175266 265131 175269
rect 265065 175264 268180 175266
rect 265065 175208 265070 175264
rect 265126 175208 268180 175264
rect 265065 175206 268180 175208
rect 265065 175203 265131 175206
rect 164550 174932 164556 174996
rect 164620 174994 164626 174996
rect 165521 174994 165587 174997
rect 164620 174992 165587 174994
rect 164620 174936 165526 174992
rect 165582 174936 165587 174992
rect 164620 174934 165587 174936
rect 164620 174932 164626 174934
rect 165521 174931 165587 174934
rect 213913 174994 213979 174997
rect 213913 174992 217028 174994
rect 213913 174936 213918 174992
rect 213974 174936 217028 174992
rect 213913 174934 217028 174936
rect 213913 174931 213979 174934
rect 264973 174858 265039 174861
rect 264973 174856 268180 174858
rect 264973 174800 264978 174856
rect 265034 174800 268180 174856
rect 264973 174798 268180 174800
rect 264973 174795 265039 174798
rect 229093 174722 229159 174725
rect 230473 174722 230539 174725
rect 280429 174722 280495 174725
rect 228988 174720 230539 174722
rect 228988 174664 229098 174720
rect 229154 174664 230478 174720
rect 230534 174664 230539 174720
rect 228988 174662 230539 174664
rect 279956 174720 280495 174722
rect 279956 174664 280434 174720
rect 280490 174664 280495 174720
rect 279956 174662 280495 174664
rect 229093 174659 229159 174662
rect 230473 174659 230539 174662
rect 280429 174659 280495 174662
rect 165429 174586 165495 174589
rect 210509 174586 210575 174589
rect 165429 174584 210575 174586
rect 165429 174528 165434 174584
rect 165490 174528 210514 174584
rect 210570 174528 210575 174584
rect 165429 174526 210575 174528
rect 165429 174523 165495 174526
rect 210509 174523 210575 174526
rect 261477 174450 261543 174453
rect 261477 174448 268180 174450
rect 261477 174392 261482 174448
rect 261538 174392 268180 174448
rect 261477 174390 268180 174392
rect 261477 174387 261543 174390
rect 214005 174314 214071 174317
rect 257337 174314 257403 174317
rect 214005 174312 217028 174314
rect 214005 174256 214010 174312
rect 214066 174256 217028 174312
rect 214005 174254 217028 174256
rect 228988 174312 257403 174314
rect 228988 174256 257342 174312
rect 257398 174256 257403 174312
rect 228988 174254 257403 174256
rect 214005 174251 214071 174254
rect 257337 174251 257403 174254
rect 229461 174042 229527 174045
rect 241697 174042 241763 174045
rect 229461 174040 241763 174042
rect 229461 173984 229466 174040
rect 229522 173984 241702 174040
rect 241758 173984 241763 174040
rect 229461 173982 241763 173984
rect 229461 173979 229527 173982
rect 241697 173979 241763 173982
rect 265249 174042 265315 174045
rect 281809 174042 281875 174045
rect 265249 174040 268180 174042
rect 265249 173984 265254 174040
rect 265310 173984 268180 174040
rect 265249 173982 268180 173984
rect 279956 174040 281875 174042
rect 279956 173984 281814 174040
rect 281870 173984 281875 174040
rect 279956 173982 281875 173984
rect 265249 173979 265315 173982
rect 281809 173979 281875 173982
rect 175917 173906 175983 173909
rect 215385 173906 215451 173909
rect 175917 173904 215451 173906
rect 175917 173848 175922 173904
rect 175978 173848 215390 173904
rect 215446 173848 215451 173904
rect 175917 173846 215451 173848
rect 175917 173843 175983 173846
rect 215385 173843 215451 173846
rect 230565 173770 230631 173773
rect 228988 173768 230631 173770
rect 228988 173712 230570 173768
rect 230626 173712 230631 173768
rect 228988 173710 230631 173712
rect 230565 173707 230631 173710
rect 279325 173770 279391 173773
rect 279325 173768 279434 173770
rect 279325 173712 279330 173768
rect 279386 173712 279434 173768
rect 279325 173707 279434 173712
rect 214465 173634 214531 173637
rect 265065 173634 265131 173637
rect 214465 173632 217028 173634
rect 214465 173576 214470 173632
rect 214526 173576 217028 173632
rect 214465 173574 217028 173576
rect 265065 173632 268180 173634
rect 265065 173576 265070 173632
rect 265126 173576 268180 173632
rect 265065 173574 268180 173576
rect 214465 173571 214531 173574
rect 265065 173571 265131 173574
rect 229369 173362 229435 173365
rect 228988 173360 229435 173362
rect 228988 173304 229374 173360
rect 229430 173304 229435 173360
rect 228988 173302 229435 173304
rect 229369 173299 229435 173302
rect 164969 173226 165035 173229
rect 215201 173226 215267 173229
rect 164969 173224 215267 173226
rect 164969 173168 164974 173224
rect 165030 173168 215206 173224
rect 215262 173168 215267 173224
rect 279374 173196 279434 173707
rect 164969 173166 215267 173168
rect 164969 173163 165035 173166
rect 215201 173163 215267 173166
rect 213913 172954 213979 172957
rect 213913 172952 217028 172954
rect 213913 172896 213918 172952
rect 213974 172896 217028 172952
rect 213913 172894 217028 172896
rect 213913 172891 213979 172894
rect 245929 172818 245995 172821
rect 228988 172816 245995 172818
rect 228988 172760 245934 172816
rect 245990 172760 245995 172816
rect 228988 172758 245995 172760
rect 245929 172755 245995 172758
rect 253289 172818 253355 172821
rect 268150 172818 268210 173060
rect 253289 172816 268210 172818
rect 253289 172760 253294 172816
rect 253350 172760 268210 172816
rect 253289 172758 268210 172760
rect 253289 172755 253355 172758
rect 264973 172682 265039 172685
rect 264973 172680 268180 172682
rect 264973 172624 264978 172680
rect 265034 172624 268180 172680
rect 264973 172622 268180 172624
rect 264973 172619 265039 172622
rect 280286 172546 280292 172548
rect 279956 172486 280292 172546
rect 280286 172484 280292 172486
rect 280356 172484 280362 172548
rect 173249 172410 173315 172413
rect 215477 172410 215543 172413
rect 231669 172410 231735 172413
rect 173249 172408 215543 172410
rect 173249 172352 173254 172408
rect 173310 172352 215482 172408
rect 215538 172352 215543 172408
rect 173249 172350 215543 172352
rect 228988 172408 231735 172410
rect 228988 172352 231674 172408
rect 231730 172352 231735 172408
rect 228988 172350 231735 172352
rect 173249 172347 173315 172350
rect 215477 172347 215543 172350
rect 231669 172347 231735 172350
rect 264237 172410 264303 172413
rect 265249 172410 265315 172413
rect 264237 172408 265315 172410
rect 264237 172352 264242 172408
rect 264298 172352 265254 172408
rect 265310 172352 265315 172408
rect 264237 172350 265315 172352
rect 264237 172347 264303 172350
rect 265249 172347 265315 172350
rect 214189 172274 214255 172277
rect 265065 172274 265131 172277
rect 279417 172274 279483 172277
rect 214189 172272 217028 172274
rect 214189 172216 214194 172272
rect 214250 172216 217028 172272
rect 214189 172214 217028 172216
rect 265065 172272 268180 172274
rect 265065 172216 265070 172272
rect 265126 172216 268180 172272
rect 265065 172214 268180 172216
rect 279374 172272 279483 172274
rect 279374 172216 279422 172272
rect 279478 172216 279483 172272
rect 214189 172211 214255 172214
rect 265065 172211 265131 172214
rect 279374 172211 279483 172216
rect 231393 171866 231459 171869
rect 228988 171864 231459 171866
rect 228988 171808 231398 171864
rect 231454 171808 231459 171864
rect 228988 171806 231459 171808
rect 231393 171803 231459 171806
rect 265157 171866 265223 171869
rect 265157 171864 268180 171866
rect 265157 171808 265162 171864
rect 265218 171808 268180 171864
rect 265157 171806 268180 171808
rect 265157 171803 265223 171806
rect 246297 171730 246363 171733
rect 255313 171730 255379 171733
rect 246297 171728 255379 171730
rect 246297 171672 246302 171728
rect 246358 171672 255318 171728
rect 255374 171672 255379 171728
rect 279374 171700 279434 172211
rect 246297 171670 255379 171672
rect 246297 171667 246363 171670
rect 255313 171667 255379 171670
rect 164724 171594 165354 171600
rect 167821 171594 167887 171597
rect 164724 171592 167887 171594
rect 164724 171540 167826 171592
rect 165294 171536 167826 171540
rect 167882 171536 167887 171592
rect 165294 171534 167887 171536
rect 167821 171531 167887 171534
rect 214097 171594 214163 171597
rect 214097 171592 217028 171594
rect 214097 171536 214102 171592
rect 214158 171536 217028 171592
rect 214097 171534 217028 171536
rect 214097 171531 214163 171534
rect 231761 171458 231827 171461
rect 228988 171456 231827 171458
rect 228988 171400 231766 171456
rect 231822 171400 231827 171456
rect 228988 171398 231827 171400
rect 231761 171395 231827 171398
rect 264973 171458 265039 171461
rect 264973 171456 268180 171458
rect 264973 171400 264978 171456
rect 265034 171400 268180 171456
rect 264973 171398 268180 171400
rect 264973 171395 265039 171398
rect 183185 171050 183251 171053
rect 214005 171050 214071 171053
rect 265065 171050 265131 171053
rect 280061 171050 280127 171053
rect 183185 171048 200130 171050
rect 183185 170992 183190 171048
rect 183246 170992 200130 171048
rect 183185 170990 200130 170992
rect 183185 170987 183251 170990
rect 200070 170914 200130 170990
rect 214005 171048 217028 171050
rect 214005 170992 214010 171048
rect 214066 170992 217028 171048
rect 214005 170990 217028 170992
rect 265065 171048 268180 171050
rect 265065 170992 265070 171048
rect 265126 170992 268180 171048
rect 265065 170990 268180 170992
rect 279926 171048 280127 171050
rect 279926 170992 280066 171048
rect 280122 170992 280127 171048
rect 279926 170990 280127 170992
rect 214005 170987 214071 170990
rect 265065 170987 265131 170990
rect 215937 170914 216003 170917
rect 229185 170914 229251 170917
rect 200070 170912 216003 170914
rect 200070 170856 215942 170912
rect 215998 170856 216003 170912
rect 200070 170854 216003 170856
rect 228988 170912 229251 170914
rect 228988 170856 229190 170912
rect 229246 170856 229251 170912
rect 279926 170884 279986 170990
rect 280061 170987 280127 170990
rect 228988 170854 229251 170856
rect 215937 170851 216003 170854
rect 229185 170851 229251 170854
rect 230749 170506 230815 170509
rect 228988 170504 230815 170506
rect 228988 170448 230754 170504
rect 230810 170448 230815 170504
rect 228988 170446 230815 170448
rect 230749 170443 230815 170446
rect 235349 170506 235415 170509
rect 242985 170506 243051 170509
rect 235349 170504 243051 170506
rect 235349 170448 235354 170504
rect 235410 170448 242990 170504
rect 243046 170448 243051 170504
rect 279325 170506 279391 170509
rect 279325 170504 279434 170506
rect 235349 170446 243051 170448
rect 235349 170443 235415 170446
rect 242985 170443 243051 170446
rect 213913 170370 213979 170373
rect 231669 170370 231735 170373
rect 240317 170370 240383 170373
rect 213913 170368 217028 170370
rect 213913 170312 213918 170368
rect 213974 170312 217028 170368
rect 213913 170310 217028 170312
rect 231669 170368 240383 170370
rect 231669 170312 231674 170368
rect 231730 170312 240322 170368
rect 240378 170312 240383 170368
rect 231669 170310 240383 170312
rect 213913 170307 213979 170310
rect 231669 170307 231735 170310
rect 240317 170307 240383 170310
rect 260097 170234 260163 170237
rect 268150 170234 268210 170476
rect 279325 170448 279330 170504
rect 279386 170448 279434 170504
rect 279325 170443 279434 170448
rect 260097 170232 268210 170234
rect 260097 170176 260102 170232
rect 260158 170176 268210 170232
rect 279374 170204 279434 170443
rect 260097 170174 268210 170176
rect 260097 170171 260163 170174
rect 264973 170098 265039 170101
rect 264973 170096 268180 170098
rect 264973 170040 264978 170096
rect 265034 170040 268180 170096
rect 264973 170038 268180 170040
rect 264973 170035 265039 170038
rect 230841 169962 230907 169965
rect 228988 169960 230907 169962
rect 228988 169904 230846 169960
rect 230902 169904 230907 169960
rect 228988 169902 230907 169904
rect 230841 169899 230907 169902
rect 240777 169826 240843 169829
rect 244365 169826 244431 169829
rect 240777 169824 244431 169826
rect 240777 169768 240782 169824
rect 240838 169768 244370 169824
rect 244426 169768 244431 169824
rect 240777 169766 244431 169768
rect 240777 169763 240843 169766
rect 244365 169763 244431 169766
rect 258717 169826 258783 169829
rect 265157 169826 265223 169829
rect 258717 169824 265223 169826
rect 258717 169768 258722 169824
rect 258778 169768 265162 169824
rect 265218 169768 265223 169824
rect 258717 169766 265223 169768
rect 258717 169763 258783 169766
rect 265157 169763 265223 169766
rect 213913 169690 213979 169693
rect 265065 169690 265131 169693
rect 213913 169688 217028 169690
rect 213913 169632 213918 169688
rect 213974 169632 217028 169688
rect 213913 169630 217028 169632
rect 265065 169688 268180 169690
rect 265065 169632 265070 169688
rect 265126 169632 268180 169688
rect 265065 169630 268180 169632
rect 213913 169627 213979 169630
rect 265065 169627 265131 169630
rect 231761 169554 231827 169557
rect 228988 169552 231827 169554
rect 228988 169496 231766 169552
rect 231822 169496 231827 169552
rect 228988 169494 231827 169496
rect 231761 169491 231827 169494
rect 281901 169418 281967 169421
rect 279956 169416 281967 169418
rect 279956 169360 281906 169416
rect 281962 169360 281967 169416
rect 279956 169358 281967 169360
rect 281901 169355 281967 169358
rect 214005 169010 214071 169013
rect 231761 169010 231827 169013
rect 214005 169008 217028 169010
rect 214005 168952 214010 169008
rect 214066 168952 217028 169008
rect 214005 168950 217028 168952
rect 228988 169008 231827 169010
rect 228988 168952 231766 169008
rect 231822 168952 231827 169008
rect 228988 168950 231827 168952
rect 214005 168947 214071 168950
rect 231761 168947 231827 168950
rect 252093 169010 252159 169013
rect 268150 169010 268210 169252
rect 252093 169008 268210 169010
rect 252093 168952 252098 169008
rect 252154 168952 268210 169008
rect 252093 168950 268210 168952
rect 252093 168947 252159 168950
rect 264973 168874 265039 168877
rect 264973 168872 268180 168874
rect 264973 168816 264978 168872
rect 265034 168816 268180 168872
rect 264973 168814 268180 168816
rect 264973 168811 265039 168814
rect 281533 168738 281599 168741
rect 279956 168736 281599 168738
rect 279956 168680 281538 168736
rect 281594 168680 281599 168736
rect 279956 168678 281599 168680
rect 281533 168675 281599 168678
rect 230933 168602 230999 168605
rect 228988 168600 230999 168602
rect 228988 168544 230938 168600
rect 230994 168544 230999 168600
rect 228988 168542 230999 168544
rect 230933 168539 230999 168542
rect 240777 168466 240843 168469
rect 241646 168466 241652 168468
rect 240777 168464 241652 168466
rect 240777 168408 240782 168464
rect 240838 168408 241652 168464
rect 240777 168406 241652 168408
rect 240777 168403 240843 168406
rect 241646 168404 241652 168406
rect 241716 168404 241722 168468
rect 265433 168466 265499 168469
rect 265433 168464 268180 168466
rect 265433 168408 265438 168464
rect 265494 168408 268180 168464
rect 265433 168406 268180 168408
rect 265433 168403 265499 168406
rect 213913 168330 213979 168333
rect 213913 168328 217028 168330
rect 213913 168272 213918 168328
rect 213974 168272 217028 168328
rect 213913 168270 217028 168272
rect 213913 168267 213979 168270
rect 231761 168058 231827 168061
rect 228988 168056 231827 168058
rect 228988 168000 231766 168056
rect 231822 168000 231827 168056
rect 228988 167998 231827 168000
rect 231761 167995 231827 167998
rect 265341 167922 265407 167925
rect 280470 167922 280476 167924
rect 265341 167920 268180 167922
rect 265341 167864 265346 167920
rect 265402 167864 268180 167920
rect 265341 167862 268180 167864
rect 279956 167862 280476 167922
rect 265341 167859 265407 167862
rect 280470 167860 280476 167862
rect 280540 167860 280546 167924
rect 214005 167650 214071 167653
rect 231485 167650 231551 167653
rect 214005 167648 217028 167650
rect 214005 167592 214010 167648
rect 214066 167592 217028 167648
rect 214005 167590 217028 167592
rect 228988 167648 231551 167650
rect 228988 167592 231490 167648
rect 231546 167592 231551 167648
rect 228988 167590 231551 167592
rect 214005 167587 214071 167590
rect 231485 167587 231551 167590
rect 279366 167588 279372 167652
rect 279436 167588 279442 167652
rect 264973 167514 265039 167517
rect 264973 167512 268180 167514
rect 264973 167456 264978 167512
rect 265034 167456 268180 167512
rect 264973 167454 268180 167456
rect 264973 167451 265039 167454
rect 262121 167242 262187 167245
rect 265617 167242 265683 167245
rect 262121 167240 265683 167242
rect 262121 167184 262126 167240
rect 262182 167184 265622 167240
rect 265678 167184 265683 167240
rect 262121 167182 265683 167184
rect 262121 167179 262187 167182
rect 265617 167179 265683 167182
rect 242893 167106 242959 167109
rect 228988 167104 242959 167106
rect 228988 167048 242898 167104
rect 242954 167048 242959 167104
rect 228988 167046 242959 167048
rect 242893 167043 242959 167046
rect 243629 167106 243695 167109
rect 243629 167104 268180 167106
rect 243629 167048 243634 167104
rect 243690 167048 268180 167104
rect 279374 167076 279434 167588
rect 243629 167046 268180 167048
rect 243629 167043 243695 167046
rect 213913 166970 213979 166973
rect 213913 166968 217028 166970
rect 213913 166912 213918 166968
rect 213974 166912 217028 166968
rect 213913 166910 217028 166912
rect 213913 166907 213979 166910
rect 234613 166834 234679 166837
rect 236494 166834 236500 166836
rect 234613 166832 236500 166834
rect 234613 166776 234618 166832
rect 234674 166776 236500 166832
rect 234613 166774 236500 166776
rect 234613 166771 234679 166774
rect 236494 166772 236500 166774
rect 236564 166772 236570 166836
rect 231761 166698 231827 166701
rect 228988 166696 231827 166698
rect 228988 166640 231766 166696
rect 231822 166640 231827 166696
rect 228988 166638 231827 166640
rect 231761 166635 231827 166638
rect 265065 166698 265131 166701
rect 265065 166696 268180 166698
rect 265065 166640 265070 166696
rect 265126 166640 268180 166696
rect 265065 166638 268180 166640
rect 265065 166635 265131 166638
rect 214005 166426 214071 166429
rect 281901 166426 281967 166429
rect 214005 166424 217028 166426
rect 214005 166368 214010 166424
rect 214066 166368 217028 166424
rect 214005 166366 217028 166368
rect 279956 166424 281967 166426
rect 279956 166368 281906 166424
rect 281962 166368 281967 166424
rect 279956 166366 281967 166368
rect 214005 166363 214071 166366
rect 281901 166363 281967 166366
rect 264973 166290 265039 166293
rect 371877 166290 371943 166293
rect 438894 166290 438900 166292
rect 264973 166288 268180 166290
rect 264973 166232 264978 166288
rect 265034 166232 268180 166288
rect 264973 166230 268180 166232
rect 371877 166288 438900 166290
rect 371877 166232 371882 166288
rect 371938 166232 438900 166288
rect 371877 166230 438900 166232
rect 264973 166227 265039 166230
rect 371877 166227 371943 166230
rect 438894 166228 438900 166230
rect 438964 166228 438970 166292
rect 231301 166154 231367 166157
rect 228988 166152 231367 166154
rect 228988 166096 231306 166152
rect 231362 166096 231367 166152
rect 228988 166094 231367 166096
rect 231301 166091 231367 166094
rect 265157 165882 265223 165885
rect 580901 165882 580967 165885
rect 583520 165882 584960 165972
rect 265157 165880 268180 165882
rect 265157 165824 265162 165880
rect 265218 165824 268180 165880
rect 265157 165822 268180 165824
rect 580901 165880 584960 165882
rect 580901 165824 580906 165880
rect 580962 165824 584960 165880
rect 580901 165822 584960 165824
rect 265157 165819 265223 165822
rect 580901 165819 580967 165822
rect 167729 165746 167795 165749
rect 233182 165746 233188 165748
rect 167729 165744 217028 165746
rect 167729 165688 167734 165744
rect 167790 165688 217028 165744
rect 167729 165686 217028 165688
rect 228988 165686 233188 165746
rect 167729 165683 167795 165686
rect 233182 165684 233188 165686
rect 233252 165684 233258 165748
rect 583520 165732 584960 165822
rect 281625 165610 281691 165613
rect 279956 165608 281691 165610
rect 279956 165552 281630 165608
rect 281686 165552 281691 165608
rect 279956 165550 281691 165552
rect 281625 165547 281691 165550
rect 265065 165338 265131 165341
rect 265065 165336 268180 165338
rect 265065 165280 265070 165336
rect 265126 165280 268180 165336
rect 265065 165278 268180 165280
rect 265065 165275 265131 165278
rect 231485 165202 231551 165205
rect 228988 165200 231551 165202
rect 228988 165144 231490 165200
rect 231546 165144 231551 165200
rect 228988 165142 231551 165144
rect 231485 165139 231551 165142
rect 213913 165066 213979 165069
rect 231393 165066 231459 165069
rect 244457 165066 244523 165069
rect 213913 165064 217028 165066
rect 213913 165008 213918 165064
rect 213974 165008 217028 165064
rect 213913 165006 217028 165008
rect 231393 165064 244523 165066
rect 231393 165008 231398 165064
rect 231454 165008 244462 165064
rect 244518 165008 244523 165064
rect 231393 165006 244523 165008
rect 213913 165003 213979 165006
rect 231393 165003 231459 165006
rect 244457 165003 244523 165006
rect 232497 164930 232563 164933
rect 265157 164930 265223 164933
rect 232497 164928 265223 164930
rect 232497 164872 232502 164928
rect 232558 164872 265162 164928
rect 265218 164872 265223 164928
rect 232497 164870 265223 164872
rect 232497 164867 232563 164870
rect 265157 164867 265223 164870
rect 265617 164930 265683 164933
rect 282821 164930 282887 164933
rect 265617 164928 268180 164930
rect 265617 164872 265622 164928
rect 265678 164872 268180 164928
rect 265617 164870 268180 164872
rect 279956 164928 282887 164930
rect 279956 164872 282826 164928
rect 282882 164872 282887 164928
rect 279956 164870 282887 164872
rect 265617 164867 265683 164870
rect 282821 164867 282887 164870
rect 231669 164794 231735 164797
rect 228988 164792 231735 164794
rect 228988 164736 231674 164792
rect 231730 164736 231735 164792
rect 228988 164734 231735 164736
rect 231669 164731 231735 164734
rect 264973 164522 265039 164525
rect 264973 164520 268180 164522
rect 264973 164464 264978 164520
rect 265034 164464 268180 164520
rect 264973 164462 268180 164464
rect 264973 164459 265039 164462
rect 215201 164386 215267 164389
rect 230933 164386 230999 164389
rect 215201 164384 217028 164386
rect 215201 164328 215206 164384
rect 215262 164328 217028 164384
rect 215201 164326 217028 164328
rect 228988 164384 230999 164386
rect 228988 164328 230938 164384
rect 230994 164328 230999 164384
rect 228988 164326 230999 164328
rect 215201 164323 215267 164326
rect 230933 164323 230999 164326
rect 265249 164114 265315 164117
rect 282821 164114 282887 164117
rect 265249 164112 268180 164114
rect 265249 164056 265254 164112
rect 265310 164056 268180 164112
rect 265249 164054 268180 164056
rect 279956 164112 282887 164114
rect 279956 164056 282826 164112
rect 282882 164056 282887 164112
rect 279956 164054 282887 164056
rect 265249 164051 265315 164054
rect 282821 164051 282887 164054
rect 231025 163842 231091 163845
rect 228988 163840 231091 163842
rect 228988 163784 231030 163840
rect 231086 163784 231091 163840
rect 228988 163782 231091 163784
rect 231025 163779 231091 163782
rect 213913 163706 213979 163709
rect 265065 163706 265131 163709
rect 213913 163704 217028 163706
rect 213913 163648 213918 163704
rect 213974 163648 217028 163704
rect 213913 163646 217028 163648
rect 265065 163704 268180 163706
rect 265065 163648 265070 163704
rect 265126 163648 268180 163704
rect 265065 163646 268180 163648
rect 213913 163643 213979 163646
rect 265065 163643 265131 163646
rect 229134 163434 229140 163436
rect 228988 163374 229140 163434
rect 229134 163372 229140 163374
rect 229204 163372 229210 163436
rect 234245 163434 234311 163437
rect 263593 163434 263659 163437
rect 234245 163432 263659 163434
rect 234245 163376 234250 163432
rect 234306 163376 263598 163432
rect 263654 163376 263659 163432
rect 234245 163374 263659 163376
rect 234245 163371 234311 163374
rect 263593 163371 263659 163374
rect 262857 163298 262923 163301
rect 281758 163298 281764 163300
rect 262857 163296 268180 163298
rect 262857 163240 262862 163296
rect 262918 163240 268180 163296
rect 262857 163238 268180 163240
rect 279956 163238 281764 163298
rect 262857 163235 262923 163238
rect 281758 163236 281764 163238
rect 281828 163236 281834 163300
rect 214005 163026 214071 163029
rect 214005 163024 217028 163026
rect -960 162890 480 162980
rect 214005 162968 214010 163024
rect 214066 162968 217028 163024
rect 214005 162966 217028 162968
rect 214005 162963 214071 162966
rect 3325 162890 3391 162893
rect 231117 162890 231183 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect 228988 162888 231183 162890
rect 228988 162832 231122 162888
rect 231178 162832 231183 162888
rect 228988 162830 231183 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 231117 162827 231183 162830
rect 264973 162890 265039 162893
rect 264973 162888 268180 162890
rect 264973 162832 264978 162888
rect 265034 162832 268180 162888
rect 264973 162830 268180 162832
rect 264973 162827 265039 162830
rect 281625 162618 281691 162621
rect 279956 162616 281691 162618
rect 279956 162560 281630 162616
rect 281686 162560 281691 162616
rect 279956 162558 281691 162560
rect 281625 162555 281691 162558
rect 237557 162482 237623 162485
rect 228988 162480 237623 162482
rect 228988 162424 237562 162480
rect 237618 162424 237623 162480
rect 228988 162422 237623 162424
rect 237557 162419 237623 162422
rect 213913 162346 213979 162349
rect 265065 162346 265131 162349
rect 213913 162344 217028 162346
rect 213913 162288 213918 162344
rect 213974 162288 217028 162344
rect 213913 162286 217028 162288
rect 265065 162344 268180 162346
rect 265065 162288 265070 162344
rect 265126 162288 268180 162344
rect 265065 162286 268180 162288
rect 213913 162283 213979 162286
rect 265065 162283 265131 162286
rect 229553 161938 229619 161941
rect 228988 161936 229619 161938
rect 228988 161880 229558 161936
rect 229614 161880 229619 161936
rect 228988 161878 229619 161880
rect 229553 161875 229619 161878
rect 258030 161878 268180 161938
rect 214005 161802 214071 161805
rect 214005 161800 217028 161802
rect 214005 161744 214010 161800
rect 214066 161744 217028 161800
rect 214005 161742 217028 161744
rect 214005 161739 214071 161742
rect 249006 161740 249012 161804
rect 249076 161802 249082 161804
rect 258030 161802 258090 161878
rect 281901 161802 281967 161805
rect 249076 161742 258090 161802
rect 279956 161800 281967 161802
rect 279956 161744 281906 161800
rect 281962 161744 281967 161800
rect 279956 161742 281967 161744
rect 249076 161740 249082 161742
rect 281901 161739 281967 161742
rect 231669 161530 231735 161533
rect 228988 161528 231735 161530
rect 228988 161472 231674 161528
rect 231730 161472 231735 161528
rect 228988 161470 231735 161472
rect 231669 161467 231735 161470
rect 265157 161530 265223 161533
rect 265157 161528 268180 161530
rect 265157 161472 265162 161528
rect 265218 161472 268180 161528
rect 265157 161470 268180 161472
rect 265157 161467 265223 161470
rect 213913 161122 213979 161125
rect 264973 161122 265039 161125
rect 282821 161122 282887 161125
rect 213913 161120 217028 161122
rect 213913 161064 213918 161120
rect 213974 161064 217028 161120
rect 213913 161062 217028 161064
rect 264973 161120 268180 161122
rect 264973 161064 264978 161120
rect 265034 161064 268180 161120
rect 264973 161062 268180 161064
rect 279956 161120 282887 161122
rect 279956 161064 282826 161120
rect 282882 161064 282887 161120
rect 279956 161062 282887 161064
rect 213913 161059 213979 161062
rect 264973 161059 265039 161062
rect 282821 161059 282887 161062
rect 236085 160986 236151 160989
rect 228988 160984 236151 160986
rect 228988 160928 236090 160984
rect 236146 160928 236151 160984
rect 228988 160926 236151 160928
rect 236085 160923 236151 160926
rect 231761 160714 231827 160717
rect 248454 160714 248460 160716
rect 231761 160712 248460 160714
rect 231761 160656 231766 160712
rect 231822 160656 248460 160712
rect 231761 160654 248460 160656
rect 231761 160651 231827 160654
rect 248454 160652 248460 160654
rect 248524 160652 248530 160716
rect 231025 160578 231091 160581
rect 228988 160576 231091 160578
rect 228988 160520 231030 160576
rect 231086 160520 231091 160576
rect 228988 160518 231091 160520
rect 231025 160515 231091 160518
rect 214005 160442 214071 160445
rect 234153 160442 234219 160445
rect 268150 160442 268210 160684
rect 214005 160440 217028 160442
rect 214005 160384 214010 160440
rect 214066 160384 217028 160440
rect 214005 160382 217028 160384
rect 234153 160440 268210 160442
rect 234153 160384 234158 160440
rect 234214 160384 268210 160440
rect 234153 160382 268210 160384
rect 214005 160379 214071 160382
rect 234153 160379 234219 160382
rect 265433 160306 265499 160309
rect 282821 160306 282887 160309
rect 265433 160304 268180 160306
rect 265433 160248 265438 160304
rect 265494 160248 268180 160304
rect 265433 160246 268180 160248
rect 279956 160304 282887 160306
rect 279956 160248 282826 160304
rect 282882 160248 282887 160304
rect 279956 160246 282887 160248
rect 265433 160243 265499 160246
rect 282821 160243 282887 160246
rect 231761 160034 231827 160037
rect 228988 160032 231827 160034
rect 228988 159976 231766 160032
rect 231822 159976 231827 160032
rect 228988 159974 231827 159976
rect 231761 159971 231827 159974
rect 213913 159762 213979 159765
rect 264973 159762 265039 159765
rect 213913 159760 217028 159762
rect 213913 159704 213918 159760
rect 213974 159704 217028 159760
rect 213913 159702 217028 159704
rect 264973 159760 268180 159762
rect 264973 159704 264978 159760
rect 265034 159704 268180 159760
rect 264973 159702 268180 159704
rect 213913 159699 213979 159702
rect 264973 159699 265039 159702
rect 237465 159626 237531 159629
rect 228988 159624 237531 159626
rect 228988 159568 237470 159624
rect 237526 159568 237531 159624
rect 228988 159566 237531 159568
rect 237465 159563 237531 159566
rect 282821 159490 282887 159493
rect 279956 159488 282887 159490
rect 279956 159432 282826 159488
rect 282882 159432 282887 159488
rect 279956 159430 282887 159432
rect 282821 159427 282887 159430
rect 267273 159354 267339 159357
rect 410517 159354 410583 159357
rect 435030 159354 435036 159356
rect 267273 159352 268180 159354
rect 267273 159296 267278 159352
rect 267334 159296 268180 159352
rect 267273 159294 268180 159296
rect 410517 159352 435036 159354
rect 410517 159296 410522 159352
rect 410578 159296 435036 159352
rect 410517 159294 435036 159296
rect 267273 159291 267339 159294
rect 410517 159291 410583 159294
rect 435030 159292 435036 159294
rect 435100 159292 435106 159356
rect 214557 159082 214623 159085
rect 247217 159082 247283 159085
rect 214557 159080 217028 159082
rect 214557 159024 214562 159080
rect 214618 159024 217028 159080
rect 214557 159022 217028 159024
rect 228988 159080 247283 159082
rect 228988 159024 247222 159080
rect 247278 159024 247283 159080
rect 228988 159022 247283 159024
rect 214557 159019 214623 159022
rect 247217 159019 247283 159022
rect 260281 159082 260347 159085
rect 265157 159082 265223 159085
rect 260281 159080 265223 159082
rect 260281 159024 260286 159080
rect 260342 159024 265162 159080
rect 265218 159024 265223 159080
rect 260281 159022 265223 159024
rect 260281 159019 260347 159022
rect 265157 159019 265223 159022
rect 265157 158946 265223 158949
rect 265157 158944 268180 158946
rect 265157 158888 265162 158944
rect 265218 158888 268180 158944
rect 265157 158886 268180 158888
rect 265157 158883 265223 158886
rect 281809 158810 281875 158813
rect 279956 158808 281875 158810
rect 279956 158752 281814 158808
rect 281870 158752 281875 158808
rect 279956 158750 281875 158752
rect 281809 158747 281875 158750
rect 231761 158674 231827 158677
rect 228988 158672 231827 158674
rect 228988 158616 231766 158672
rect 231822 158616 231827 158672
rect 228988 158614 231827 158616
rect 231761 158611 231827 158614
rect 265065 158538 265131 158541
rect 265065 158536 268180 158538
rect 265065 158480 265070 158536
rect 265126 158480 268180 158536
rect 265065 158478 268180 158480
rect 265065 158475 265131 158478
rect 213913 158402 213979 158405
rect 213913 158400 217028 158402
rect 213913 158344 213918 158400
rect 213974 158344 217028 158400
rect 213913 158342 217028 158344
rect 213913 158339 213979 158342
rect 231485 158130 231551 158133
rect 228988 158128 231551 158130
rect 228988 158072 231490 158128
rect 231546 158072 231551 158128
rect 228988 158070 231551 158072
rect 231485 158067 231551 158070
rect 231669 157994 231735 157997
rect 246297 157994 246363 157997
rect 231669 157992 246363 157994
rect 231669 157936 231674 157992
rect 231730 157936 246302 157992
rect 246358 157936 246363 157992
rect 231669 157934 246363 157936
rect 231669 157931 231735 157934
rect 246297 157931 246363 157934
rect 229829 157858 229895 157861
rect 268150 157858 268210 158100
rect 282085 157994 282151 157997
rect 279956 157992 282151 157994
rect 279956 157936 282090 157992
rect 282146 157936 282151 157992
rect 279956 157934 282151 157936
rect 282085 157931 282151 157934
rect 229829 157856 268210 157858
rect 229829 157800 229834 157856
rect 229890 157800 268210 157856
rect 229829 157798 268210 157800
rect 229829 157795 229895 157798
rect 214005 157722 214071 157725
rect 230657 157722 230723 157725
rect 214005 157720 217028 157722
rect 214005 157664 214010 157720
rect 214066 157664 217028 157720
rect 214005 157662 217028 157664
rect 228988 157720 230723 157722
rect 228988 157664 230662 157720
rect 230718 157664 230723 157720
rect 228988 157662 230723 157664
rect 214005 157659 214071 157662
rect 230657 157659 230723 157662
rect 264973 157722 265039 157725
rect 264973 157720 268180 157722
rect 264973 157664 264978 157720
rect 265034 157664 268180 157720
rect 264973 157662 268180 157664
rect 264973 157659 265039 157662
rect 281717 157314 281783 157317
rect 279956 157312 281783 157314
rect 279956 157256 281722 157312
rect 281778 157256 281783 157312
rect 279956 157254 281783 157256
rect 281717 157251 281783 157254
rect 213913 157178 213979 157181
rect 231669 157178 231735 157181
rect 213913 157176 217028 157178
rect 213913 157120 213918 157176
rect 213974 157120 217028 157176
rect 213913 157118 217028 157120
rect 228988 157176 231735 157178
rect 228988 157120 231674 157176
rect 231730 157120 231735 157176
rect 228988 157118 231735 157120
rect 213913 157115 213979 157118
rect 231669 157115 231735 157118
rect 265065 157178 265131 157181
rect 265065 157176 268180 157178
rect 265065 157120 265070 157176
rect 265126 157120 268180 157176
rect 265065 157118 268180 157120
rect 265065 157115 265131 157118
rect 231761 156770 231827 156773
rect 253197 156770 253263 156773
rect 228988 156768 231827 156770
rect 228988 156712 231766 156768
rect 231822 156712 231827 156768
rect 228988 156710 231827 156712
rect 231761 156707 231827 156710
rect 231902 156768 253263 156770
rect 231902 156712 253202 156768
rect 253258 156712 253263 156768
rect 231902 156710 253263 156712
rect 231209 156634 231275 156637
rect 231902 156634 231962 156710
rect 253197 156707 253263 156710
rect 264973 156770 265039 156773
rect 264973 156768 268180 156770
rect 264973 156712 264978 156768
rect 265034 156712 268180 156768
rect 264973 156710 268180 156712
rect 264973 156707 265039 156710
rect 231209 156632 231962 156634
rect 231209 156576 231214 156632
rect 231270 156576 231962 156632
rect 231209 156574 231962 156576
rect 236729 156634 236795 156637
rect 265157 156634 265223 156637
rect 236729 156632 265223 156634
rect 236729 156576 236734 156632
rect 236790 156576 265162 156632
rect 265218 156576 265223 156632
rect 236729 156574 265223 156576
rect 231209 156571 231275 156574
rect 236729 156571 236795 156574
rect 265157 156571 265223 156574
rect 214005 156498 214071 156501
rect 281574 156498 281580 156500
rect 214005 156496 217028 156498
rect 214005 156440 214010 156496
rect 214066 156440 217028 156496
rect 214005 156438 217028 156440
rect 279956 156438 281580 156498
rect 214005 156435 214071 156438
rect 281574 156436 281580 156438
rect 281644 156436 281650 156500
rect 265157 156362 265223 156365
rect 265157 156360 268180 156362
rect 265157 156304 265162 156360
rect 265218 156304 268180 156360
rect 265157 156302 268180 156304
rect 265157 156299 265223 156302
rect 237598 156226 237604 156228
rect 228988 156166 237604 156226
rect 237598 156164 237604 156166
rect 237668 156164 237674 156228
rect 265065 155954 265131 155957
rect 265065 155952 268180 155954
rect 265065 155896 265070 155952
rect 265126 155896 268180 155952
rect 265065 155894 268180 155896
rect 265065 155891 265131 155894
rect 213913 155818 213979 155821
rect 231761 155818 231827 155821
rect 213913 155816 217028 155818
rect 213913 155760 213918 155816
rect 213974 155760 217028 155816
rect 213913 155758 217028 155760
rect 228988 155816 231827 155818
rect 228988 155760 231766 155816
rect 231822 155760 231827 155816
rect 228988 155758 231827 155760
rect 213913 155755 213979 155758
rect 231761 155755 231827 155758
rect 281533 155682 281599 155685
rect 279956 155680 281599 155682
rect 279956 155624 281538 155680
rect 281594 155624 281599 155680
rect 279956 155622 281599 155624
rect 281533 155619 281599 155622
rect 264973 155546 265039 155549
rect 264973 155544 268180 155546
rect 264973 155488 264978 155544
rect 265034 155488 268180 155544
rect 264973 155486 268180 155488
rect 264973 155483 265039 155486
rect 230565 155274 230631 155277
rect 228988 155272 230631 155274
rect 228988 155216 230570 155272
rect 230626 155216 230631 155272
rect 228988 155214 230631 155216
rect 230565 155211 230631 155214
rect 231761 155274 231827 155277
rect 243169 155274 243235 155277
rect 231761 155272 243235 155274
rect 231761 155216 231766 155272
rect 231822 155216 243174 155272
rect 243230 155216 243235 155272
rect 231761 155214 243235 155216
rect 231761 155211 231827 155214
rect 243169 155211 243235 155214
rect 214005 155138 214071 155141
rect 214005 155136 217028 155138
rect 214005 155080 214010 155136
rect 214066 155080 217028 155136
rect 214005 155078 217028 155080
rect 214005 155075 214071 155078
rect 231209 154866 231275 154869
rect 228988 154864 231275 154866
rect 228988 154808 231214 154864
rect 231270 154808 231275 154864
rect 228988 154806 231275 154808
rect 231209 154803 231275 154806
rect 243813 154866 243879 154869
rect 268150 154866 268210 155108
rect 282269 155002 282335 155005
rect 279956 155000 282335 155002
rect 279956 154944 282274 155000
rect 282330 154944 282335 155000
rect 279956 154942 282335 154944
rect 282269 154939 282335 154942
rect 243813 154864 268210 154866
rect 243813 154808 243818 154864
rect 243874 154808 268210 154864
rect 243813 154806 268210 154808
rect 243813 154803 243879 154806
rect 265709 154594 265775 154597
rect 265709 154592 268180 154594
rect 265709 154536 265714 154592
rect 265770 154536 268180 154592
rect 265709 154534 268180 154536
rect 265709 154531 265775 154534
rect 214005 154458 214071 154461
rect 231301 154458 231367 154461
rect 238518 154458 238524 154460
rect 214005 154456 217028 154458
rect 214005 154400 214010 154456
rect 214066 154400 217028 154456
rect 214005 154398 217028 154400
rect 231301 154456 238524 154458
rect 231301 154400 231306 154456
rect 231362 154400 238524 154456
rect 231301 154398 238524 154400
rect 214005 154395 214071 154398
rect 231301 154395 231367 154398
rect 238518 154396 238524 154398
rect 238588 154396 238594 154460
rect 231761 154322 231827 154325
rect 228988 154320 231827 154322
rect 228988 154264 231766 154320
rect 231822 154264 231827 154320
rect 228988 154262 231827 154264
rect 231761 154259 231827 154262
rect 264973 154186 265039 154189
rect 282085 154186 282151 154189
rect 264973 154184 268180 154186
rect 264973 154128 264978 154184
rect 265034 154128 268180 154184
rect 264973 154126 268180 154128
rect 279956 154184 282151 154186
rect 279956 154128 282090 154184
rect 282146 154128 282151 154184
rect 279956 154126 282151 154128
rect 264973 154123 265039 154126
rect 282085 154123 282151 154126
rect 231393 153914 231459 153917
rect 228988 153912 231459 153914
rect 228988 153856 231398 153912
rect 231454 153856 231459 153912
rect 228988 153854 231459 153856
rect 231393 153851 231459 153854
rect 231761 153914 231827 153917
rect 249926 153914 249932 153916
rect 231761 153912 249932 153914
rect 231761 153856 231766 153912
rect 231822 153856 249932 153912
rect 231761 153854 249932 153856
rect 231761 153851 231827 153854
rect 249926 153852 249932 153854
rect 249996 153852 250002 153916
rect 213913 153778 213979 153781
rect 246481 153778 246547 153781
rect 265157 153778 265223 153781
rect 213913 153776 217028 153778
rect 213913 153720 213918 153776
rect 213974 153720 217028 153776
rect 213913 153718 217028 153720
rect 246481 153776 265223 153778
rect 246481 153720 246486 153776
rect 246542 153720 265162 153776
rect 265218 153720 265223 153776
rect 246481 153718 265223 153720
rect 213913 153715 213979 153718
rect 246481 153715 246547 153718
rect 265157 153715 265223 153718
rect 264421 153506 264487 153509
rect 268150 153506 268210 153748
rect 282821 153506 282887 153509
rect 264421 153504 268210 153506
rect 264421 153448 264426 153504
rect 264482 153448 268210 153504
rect 264421 153446 268210 153448
rect 279956 153504 282887 153506
rect 279956 153448 282826 153504
rect 282882 153448 282887 153504
rect 279956 153446 282887 153448
rect 264421 153443 264487 153446
rect 282821 153443 282887 153446
rect 231209 153370 231275 153373
rect 228988 153368 231275 153370
rect 228988 153312 231214 153368
rect 231270 153312 231275 153368
rect 228988 153310 231275 153312
rect 231209 153307 231275 153310
rect 258030 153310 268180 153370
rect 239581 153234 239647 153237
rect 258030 153234 258090 153310
rect 239581 153232 258090 153234
rect 239581 153176 239586 153232
rect 239642 153176 258090 153232
rect 239581 153174 258090 153176
rect 239581 153171 239647 153174
rect 213913 153098 213979 153101
rect 230565 153098 230631 153101
rect 252553 153098 252619 153101
rect 213913 153096 217028 153098
rect 213913 153040 213918 153096
rect 213974 153040 217028 153096
rect 213913 153038 217028 153040
rect 230565 153096 252619 153098
rect 230565 153040 230570 153096
rect 230626 153040 252558 153096
rect 252614 153040 252619 153096
rect 230565 153038 252619 153040
rect 213913 153035 213979 153038
rect 230565 153035 230631 153038
rect 252553 153035 252619 153038
rect 231761 152962 231827 152965
rect 228988 152960 231827 152962
rect 228988 152904 231766 152960
rect 231822 152904 231827 152960
rect 228988 152902 231827 152904
rect 231761 152899 231827 152902
rect 265065 152962 265131 152965
rect 265065 152960 268180 152962
rect 265065 152904 265070 152960
rect 265126 152904 268180 152960
rect 265065 152902 268180 152904
rect 265065 152899 265131 152902
rect 282177 152690 282243 152693
rect 583520 152690 584960 152780
rect 279956 152688 282243 152690
rect 279956 152632 282182 152688
rect 282238 152632 282243 152688
rect 279956 152630 282243 152632
rect 282177 152627 282243 152630
rect 583342 152630 584960 152690
rect 214005 152554 214071 152557
rect 244222 152554 244228 152556
rect 214005 152552 217028 152554
rect 214005 152496 214010 152552
rect 214066 152496 217028 152552
rect 214005 152494 217028 152496
rect 228988 152494 244228 152554
rect 214005 152491 214071 152494
rect 244222 152492 244228 152494
rect 244292 152492 244298 152556
rect 264973 152554 265039 152557
rect 583342 152554 583402 152630
rect 583520 152554 584960 152630
rect 264973 152552 268180 152554
rect 264973 152496 264978 152552
rect 265034 152496 268180 152552
rect 264973 152494 268180 152496
rect 583342 152540 584960 152554
rect 583342 152494 583586 152540
rect 264973 152491 265039 152494
rect 583526 152282 583586 152494
rect 583661 152282 583727 152285
rect 583526 152280 583727 152282
rect 583526 152224 583666 152280
rect 583722 152224 583727 152280
rect 583526 152222 583727 152224
rect 583661 152219 583727 152222
rect 230565 152010 230631 152013
rect 228988 152008 230631 152010
rect 228988 151952 230570 152008
rect 230626 151952 230631 152008
rect 228988 151950 230631 151952
rect 230565 151947 230631 151950
rect 265801 152010 265867 152013
rect 265801 152008 268180 152010
rect 265801 151952 265806 152008
rect 265862 151952 268180 152008
rect 265801 151950 268180 151952
rect 265801 151947 265867 151950
rect 214557 151874 214623 151877
rect 280337 151874 280403 151877
rect 214557 151872 217028 151874
rect 214557 151816 214562 151872
rect 214618 151816 217028 151872
rect 214557 151814 217028 151816
rect 279956 151872 280403 151874
rect 279956 151816 280342 151872
rect 280398 151816 280403 151872
rect 279956 151814 280403 151816
rect 214557 151811 214623 151814
rect 280337 151811 280403 151814
rect 230473 151602 230539 151605
rect 228988 151600 230539 151602
rect 228988 151544 230478 151600
rect 230534 151544 230539 151600
rect 228988 151542 230539 151544
rect 230473 151539 230539 151542
rect 265341 151602 265407 151605
rect 265341 151600 268180 151602
rect 265341 151544 265346 151600
rect 265402 151544 268180 151600
rect 265341 151542 268180 151544
rect 265341 151539 265407 151542
rect 214005 151194 214071 151197
rect 281901 151194 281967 151197
rect 214005 151192 217028 151194
rect 214005 151136 214010 151192
rect 214066 151136 217028 151192
rect 279956 151192 281967 151194
rect 214005 151134 217028 151136
rect 214005 151131 214071 151134
rect 184841 151058 184907 151061
rect 215886 151058 215892 151060
rect 184841 151056 215892 151058
rect 184841 151000 184846 151056
rect 184902 151000 215892 151056
rect 184841 150998 215892 151000
rect 184841 150995 184907 150998
rect 215886 150996 215892 150998
rect 215956 150996 215962 151060
rect 230657 151058 230723 151061
rect 228988 151056 230723 151058
rect 228988 151000 230662 151056
rect 230718 151000 230723 151056
rect 228988 150998 230723 151000
rect 230657 150995 230723 150998
rect 231669 151058 231735 151061
rect 247125 151058 247191 151061
rect 231669 151056 247191 151058
rect 231669 151000 231674 151056
rect 231730 151000 247130 151056
rect 247186 151000 247191 151056
rect 231669 150998 247191 151000
rect 231669 150995 231735 150998
rect 247125 150995 247191 150998
rect 244917 150922 244983 150925
rect 268150 150922 268210 151164
rect 279956 151136 281906 151192
rect 281962 151136 281967 151192
rect 279956 151134 281967 151136
rect 281901 151131 281967 151134
rect 244917 150920 268210 150922
rect 244917 150864 244922 150920
rect 244978 150864 268210 150920
rect 244917 150862 268210 150864
rect 244917 150859 244983 150862
rect 265065 150786 265131 150789
rect 265065 150784 268180 150786
rect 265065 150728 265070 150784
rect 265126 150728 268180 150784
rect 265065 150726 268180 150728
rect 265065 150723 265131 150726
rect 230422 150650 230428 150652
rect 228988 150590 230428 150650
rect 230422 150588 230428 150590
rect 230492 150588 230498 150652
rect 213913 150514 213979 150517
rect 213913 150512 217028 150514
rect 213913 150456 213918 150512
rect 213974 150456 217028 150512
rect 213913 150454 217028 150456
rect 213913 150451 213979 150454
rect 282821 150378 282887 150381
rect 279956 150376 282887 150378
rect 241513 150106 241579 150109
rect 268150 150106 268210 150348
rect 279956 150320 282826 150376
rect 282882 150320 282887 150376
rect 279956 150318 282887 150320
rect 282821 150315 282887 150318
rect 228988 150104 241579 150106
rect 228988 150048 241518 150104
rect 241574 150048 241579 150104
rect 228988 150046 241579 150048
rect 241513 150043 241579 150046
rect 258030 150046 268210 150106
rect -960 149834 480 149924
rect 3601 149834 3667 149837
rect -960 149832 3667 149834
rect -960 149776 3606 149832
rect 3662 149776 3667 149832
rect -960 149774 3667 149776
rect -960 149684 480 149774
rect 3601 149771 3667 149774
rect 213913 149834 213979 149837
rect 213913 149832 217028 149834
rect 213913 149776 213918 149832
rect 213974 149776 217028 149832
rect 213913 149774 217028 149776
rect 213913 149771 213979 149774
rect 234654 149698 234660 149700
rect 228988 149638 234660 149698
rect 234654 149636 234660 149638
rect 234724 149636 234730 149700
rect 242341 149698 242407 149701
rect 258030 149698 258090 150046
rect 264973 149970 265039 149973
rect 264973 149968 268180 149970
rect 264973 149912 264978 149968
rect 265034 149912 268180 149968
rect 264973 149910 268180 149912
rect 264973 149907 265039 149910
rect 282729 149698 282795 149701
rect 242341 149696 258090 149698
rect 242341 149640 242346 149696
rect 242402 149640 258090 149696
rect 242341 149638 258090 149640
rect 279956 149696 282795 149698
rect 279956 149640 282734 149696
rect 282790 149640 282795 149696
rect 279956 149638 282795 149640
rect 242341 149635 242407 149638
rect 282729 149635 282795 149638
rect 214005 149154 214071 149157
rect 240133 149154 240199 149157
rect 268150 149154 268210 149532
rect 214005 149152 217028 149154
rect 214005 149096 214010 149152
rect 214066 149096 217028 149152
rect 214005 149094 217028 149096
rect 228988 149152 240199 149154
rect 228988 149096 240138 149152
rect 240194 149096 240199 149152
rect 228988 149094 240199 149096
rect 214005 149091 214071 149094
rect 240133 149091 240199 149094
rect 265022 149094 268210 149154
rect 295333 149154 295399 149157
rect 295926 149154 295932 149156
rect 295333 149152 295932 149154
rect 295333 149096 295338 149152
rect 295394 149096 295932 149152
rect 295333 149094 295932 149096
rect 264094 148956 264100 149020
rect 264164 149018 264170 149020
rect 265022 149018 265082 149094
rect 295333 149091 295399 149094
rect 295926 149092 295932 149094
rect 295996 149154 296002 149156
rect 425145 149154 425211 149157
rect 295996 149152 425211 149154
rect 295996 149096 425150 149152
rect 425206 149096 425211 149152
rect 295996 149094 425211 149096
rect 295996 149092 296002 149094
rect 425145 149091 425211 149094
rect 264164 148958 265082 149018
rect 265617 149018 265683 149021
rect 265617 149016 268180 149018
rect 265617 148960 265622 149016
rect 265678 148960 268180 149016
rect 265617 148958 268180 148960
rect 264164 148956 264170 148958
rect 265617 148955 265683 148958
rect 282821 148882 282887 148885
rect 279956 148880 282887 148882
rect 279956 148824 282826 148880
rect 282882 148824 282887 148880
rect 279956 148822 282887 148824
rect 282821 148819 282887 148822
rect 229093 148746 229159 148749
rect 228988 148744 229159 148746
rect 228988 148688 229098 148744
rect 229154 148688 229159 148744
rect 228988 148686 229159 148688
rect 229093 148683 229159 148686
rect 265157 148610 265223 148613
rect 265157 148608 268180 148610
rect 265157 148552 265162 148608
rect 265218 148552 268180 148608
rect 265157 148550 268180 148552
rect 265157 148547 265223 148550
rect 213913 148474 213979 148477
rect 213913 148472 217028 148474
rect 213913 148416 213918 148472
rect 213974 148416 217028 148472
rect 213913 148414 217028 148416
rect 213913 148411 213979 148414
rect 231485 148338 231551 148341
rect 237414 148338 237420 148340
rect 231485 148336 237420 148338
rect 231485 148280 231490 148336
rect 231546 148280 237420 148336
rect 231485 148278 237420 148280
rect 231485 148275 231551 148278
rect 237414 148276 237420 148278
rect 237484 148276 237490 148340
rect 253381 148338 253447 148341
rect 265065 148338 265131 148341
rect 253381 148336 265131 148338
rect 253381 148280 253386 148336
rect 253442 148280 265070 148336
rect 265126 148280 265131 148336
rect 253381 148278 265131 148280
rect 253381 148275 253447 148278
rect 265065 148275 265131 148278
rect 388437 148338 388503 148341
rect 443177 148338 443243 148341
rect 388437 148336 443243 148338
rect 388437 148280 388442 148336
rect 388498 148280 443182 148336
rect 443238 148280 443243 148336
rect 388437 148278 443243 148280
rect 388437 148275 388503 148278
rect 443177 148275 443243 148278
rect 245745 148202 245811 148205
rect 228988 148200 245811 148202
rect 228988 148144 245750 148200
rect 245806 148144 245811 148200
rect 228988 148142 245811 148144
rect 245745 148139 245811 148142
rect 265065 148202 265131 148205
rect 265065 148200 268180 148202
rect 265065 148144 265070 148200
rect 265126 148144 268180 148200
rect 265065 148142 268180 148144
rect 265065 148139 265131 148142
rect 282177 148066 282243 148069
rect 279956 148064 282243 148066
rect 279956 148008 282182 148064
rect 282238 148008 282243 148064
rect 279956 148006 282243 148008
rect 282177 148003 282243 148006
rect 213913 147930 213979 147933
rect 213913 147928 217028 147930
rect 213913 147872 213918 147928
rect 213974 147872 217028 147928
rect 213913 147870 217028 147872
rect 213913 147867 213979 147870
rect 230565 147794 230631 147797
rect 228988 147792 230631 147794
rect 228988 147736 230570 147792
rect 230626 147736 230631 147792
rect 228988 147734 230631 147736
rect 230565 147731 230631 147734
rect 264973 147794 265039 147797
rect 264973 147792 268180 147794
rect 264973 147736 264978 147792
rect 265034 147736 268180 147792
rect 264973 147734 268180 147736
rect 264973 147731 265039 147734
rect 265065 147386 265131 147389
rect 281717 147386 281783 147389
rect 265065 147384 268180 147386
rect 265065 147328 265070 147384
rect 265126 147328 268180 147384
rect 265065 147326 268180 147328
rect 279956 147384 281783 147386
rect 279956 147328 281722 147384
rect 281778 147328 281783 147384
rect 279956 147326 281783 147328
rect 265065 147323 265131 147326
rect 281717 147323 281783 147326
rect 214005 147250 214071 147253
rect 229737 147250 229803 147253
rect 214005 147248 217028 147250
rect 214005 147192 214010 147248
rect 214066 147192 217028 147248
rect 214005 147190 217028 147192
rect 228988 147248 229803 147250
rect 228988 147192 229742 147248
rect 229798 147192 229803 147248
rect 228988 147190 229803 147192
rect 214005 147187 214071 147190
rect 229737 147187 229803 147190
rect 236494 146916 236500 146980
rect 236564 146978 236570 146980
rect 236637 146978 236703 146981
rect 236564 146976 236703 146978
rect 236564 146920 236642 146976
rect 236698 146920 236703 146976
rect 406009 146978 406075 146981
rect 582649 146978 582715 146981
rect 406009 146976 582715 146978
rect 236564 146918 236703 146920
rect 236564 146916 236570 146918
rect 236637 146915 236703 146918
rect 231761 146842 231827 146845
rect 228988 146840 231827 146842
rect 228988 146784 231766 146840
rect 231822 146784 231827 146840
rect 228988 146782 231827 146784
rect 231761 146779 231827 146782
rect 236821 146706 236887 146709
rect 268150 146706 268210 146948
rect 406009 146920 406014 146976
rect 406070 146920 582654 146976
rect 582710 146920 582715 146976
rect 406009 146918 582715 146920
rect 406009 146915 406075 146918
rect 582649 146915 582715 146918
rect 236821 146704 268210 146706
rect 236821 146648 236826 146704
rect 236882 146648 268210 146704
rect 236821 146646 268210 146648
rect 236821 146643 236887 146646
rect 213913 146570 213979 146573
rect 282821 146570 282887 146573
rect 213913 146568 217028 146570
rect 213913 146512 213918 146568
rect 213974 146512 217028 146568
rect 213913 146510 217028 146512
rect 279956 146568 282887 146570
rect 279956 146512 282826 146568
rect 282882 146512 282887 146568
rect 279956 146510 282887 146512
rect 213913 146507 213979 146510
rect 282821 146507 282887 146510
rect 264973 146434 265039 146437
rect 264973 146432 268180 146434
rect 264973 146376 264978 146432
rect 265034 146376 268180 146432
rect 264973 146374 268180 146376
rect 264973 146371 265039 146374
rect 230565 146300 230631 146301
rect 230565 146298 230612 146300
rect 228988 146238 230306 146298
rect 230520 146296 230612 146298
rect 230520 146240 230570 146296
rect 230520 146238 230612 146240
rect 230246 146162 230306 146238
rect 230565 146236 230612 146238
rect 230676 146236 230682 146300
rect 395981 146298 396047 146301
rect 399569 146298 399635 146301
rect 395981 146296 399635 146298
rect 395981 146240 395986 146296
rect 396042 146240 399574 146296
rect 399630 146240 399635 146296
rect 395981 146238 399635 146240
rect 230565 146235 230631 146236
rect 395981 146235 396047 146238
rect 399569 146235 399635 146238
rect 231761 146162 231827 146165
rect 230246 146160 231827 146162
rect 230246 146104 231766 146160
rect 231822 146104 231827 146160
rect 230246 146102 231827 146104
rect 231761 146099 231827 146102
rect 265157 146026 265223 146029
rect 265157 146024 268180 146026
rect 265157 145968 265162 146024
rect 265218 145968 268180 146024
rect 265157 145966 268180 145968
rect 265157 145963 265223 145966
rect 242433 145890 242499 145893
rect 282821 145890 282887 145893
rect 228988 145888 242499 145890
rect 216998 145346 217058 145860
rect 228988 145832 242438 145888
rect 242494 145832 242499 145888
rect 228988 145830 242499 145832
rect 279956 145888 282887 145890
rect 279956 145832 282826 145888
rect 282882 145832 282887 145888
rect 279956 145830 282887 145832
rect 242433 145827 242499 145830
rect 282821 145827 282887 145830
rect 264973 145754 265039 145757
rect 258030 145752 265039 145754
rect 258030 145696 264978 145752
rect 265034 145696 265039 145752
rect 258030 145694 265039 145696
rect 232446 145556 232452 145620
rect 232516 145618 232522 145620
rect 258030 145618 258090 145694
rect 264973 145691 265039 145694
rect 232516 145558 258090 145618
rect 265065 145618 265131 145621
rect 265065 145616 268180 145618
rect 265065 145560 265070 145616
rect 265126 145560 268180 145616
rect 265065 145558 268180 145560
rect 232516 145556 232522 145558
rect 265065 145555 265131 145558
rect 231894 145346 231900 145348
rect 200070 145286 217058 145346
rect 228988 145286 231900 145346
rect 166206 144876 166212 144940
rect 166276 144938 166282 144940
rect 200070 144938 200130 145286
rect 231894 145284 231900 145286
rect 231964 145284 231970 145348
rect 213913 145210 213979 145213
rect 264973 145210 265039 145213
rect 213913 145208 217028 145210
rect 213913 145152 213918 145208
rect 213974 145152 217028 145208
rect 213913 145150 217028 145152
rect 264973 145208 268180 145210
rect 264973 145152 264978 145208
rect 265034 145152 268180 145208
rect 264973 145150 268180 145152
rect 213913 145147 213979 145150
rect 264973 145147 265039 145150
rect 280337 145074 280403 145077
rect 279956 145072 280403 145074
rect 279956 145016 280342 145072
rect 280398 145016 280403 145072
rect 279956 145014 280403 145016
rect 280337 145011 280403 145014
rect 231485 144938 231551 144941
rect 166276 144878 200130 144938
rect 228988 144936 231551 144938
rect 228988 144880 231490 144936
rect 231546 144880 231551 144936
rect 228988 144878 231551 144880
rect 166276 144876 166282 144878
rect 231485 144875 231551 144878
rect 249742 144802 249748 144804
rect 238710 144742 249748 144802
rect 214189 144530 214255 144533
rect 214189 144528 217028 144530
rect 214189 144472 214194 144528
rect 214250 144472 217028 144528
rect 214189 144470 217028 144472
rect 214189 144467 214255 144470
rect 238710 144394 238770 144742
rect 249742 144740 249748 144742
rect 249812 144740 249818 144804
rect 264973 144802 265039 144805
rect 264973 144800 268180 144802
rect 264973 144744 264978 144800
rect 265034 144744 268180 144800
rect 264973 144742 268180 144744
rect 264973 144739 265039 144742
rect 228988 144334 238770 144394
rect 265249 144394 265315 144397
rect 265249 144392 268180 144394
rect 265249 144336 265254 144392
rect 265310 144336 268180 144392
rect 265249 144334 268180 144336
rect 265249 144331 265315 144334
rect 282821 144258 282887 144261
rect 279956 144256 282887 144258
rect 279956 144200 282826 144256
rect 282882 144200 282887 144256
rect 279956 144198 282887 144200
rect 282821 144195 282887 144198
rect 231710 144060 231716 144124
rect 231780 144122 231786 144124
rect 251173 144122 251239 144125
rect 231780 144120 251239 144122
rect 231780 144064 251178 144120
rect 251234 144064 251239 144120
rect 231780 144062 251239 144064
rect 231780 144060 231786 144062
rect 251173 144059 251239 144062
rect 231761 143986 231827 143989
rect 228988 143984 231827 143986
rect 228988 143928 231766 143984
rect 231822 143928 231827 143984
rect 228988 143926 231827 143928
rect 231761 143923 231827 143926
rect 213913 143850 213979 143853
rect 264605 143850 264671 143853
rect 213913 143848 217028 143850
rect 213913 143792 213918 143848
rect 213974 143792 217028 143848
rect 213913 143790 217028 143792
rect 264605 143848 268180 143850
rect 264605 143792 264610 143848
rect 264666 143792 268180 143848
rect 264605 143790 268180 143792
rect 213913 143787 213979 143790
rect 264605 143787 264671 143790
rect 280797 143578 280863 143581
rect 279956 143576 280863 143578
rect 279956 143520 280802 143576
rect 280858 143520 280863 143576
rect 279956 143518 280863 143520
rect 280797 143515 280863 143518
rect 360929 143578 360995 143581
rect 433517 143578 433583 143581
rect 360929 143576 433583 143578
rect 360929 143520 360934 143576
rect 360990 143520 433522 143576
rect 433578 143520 433583 143576
rect 360929 143518 433583 143520
rect 360929 143515 360995 143518
rect 433517 143515 433583 143518
rect 231669 143442 231735 143445
rect 228988 143440 231735 143442
rect 228988 143384 231674 143440
rect 231730 143384 231735 143440
rect 228988 143382 231735 143384
rect 231669 143379 231735 143382
rect 265065 143442 265131 143445
rect 415393 143442 415459 143445
rect 416129 143442 416195 143445
rect 265065 143440 268180 143442
rect 265065 143384 265070 143440
rect 265126 143384 268180 143440
rect 265065 143382 268180 143384
rect 415393 143440 416195 143442
rect 415393 143384 415398 143440
rect 415454 143384 416134 143440
rect 416190 143384 416195 143440
rect 415393 143382 416195 143384
rect 265065 143379 265131 143382
rect 415393 143379 415459 143382
rect 416129 143379 416195 143382
rect 425053 143442 425119 143445
rect 425789 143442 425855 143445
rect 425053 143440 425855 143442
rect 425053 143384 425058 143440
rect 425114 143384 425794 143440
rect 425850 143384 425855 143440
rect 425053 143382 425855 143384
rect 425053 143379 425119 143382
rect 425789 143379 425855 143382
rect 214005 143306 214071 143309
rect 214005 143304 217028 143306
rect 214005 143248 214010 143304
rect 214066 143248 217028 143304
rect 214005 143246 217028 143248
rect 214005 143243 214071 143246
rect 247769 143170 247835 143173
rect 238710 143168 247835 143170
rect 238710 143112 247774 143168
rect 247830 143112 247835 143168
rect 238710 143110 247835 143112
rect 231710 143034 231716 143036
rect 228988 142974 231716 143034
rect 231710 142972 231716 142974
rect 231780 142972 231786 143036
rect 230974 142836 230980 142900
rect 231044 142898 231050 142900
rect 238710 142898 238770 143110
rect 247769 143107 247835 143110
rect 240777 143034 240843 143037
rect 249006 143034 249012 143036
rect 240777 143032 249012 143034
rect 240777 142976 240782 143032
rect 240838 142976 249012 143032
rect 240777 142974 249012 142976
rect 240777 142971 240843 142974
rect 249006 142972 249012 142974
rect 249076 142972 249082 143036
rect 265709 143034 265775 143037
rect 265709 143032 268180 143034
rect 265709 142976 265714 143032
rect 265770 142976 268180 143032
rect 265709 142974 268180 142976
rect 265709 142971 265775 142974
rect 231044 142838 238770 142898
rect 241513 142898 241579 142901
rect 242014 142898 242020 142900
rect 241513 142896 242020 142898
rect 241513 142840 241518 142896
rect 241574 142840 242020 142896
rect 241513 142838 242020 142840
rect 231044 142836 231050 142838
rect 241513 142835 241579 142838
rect 242014 142836 242020 142838
rect 242084 142836 242090 142900
rect 231158 142700 231164 142764
rect 231228 142762 231234 142764
rect 261477 142762 261543 142765
rect 283097 142762 283163 142765
rect 231228 142760 261543 142762
rect 231228 142704 261482 142760
rect 261538 142704 261543 142760
rect 231228 142702 261543 142704
rect 279956 142760 283163 142762
rect 279956 142704 283102 142760
rect 283158 142704 283163 142760
rect 279956 142702 283163 142704
rect 231228 142700 231234 142702
rect 261477 142699 261543 142702
rect 283097 142699 283163 142702
rect 395337 142762 395403 142765
rect 412633 142762 412699 142765
rect 415485 142762 415551 142765
rect 395337 142760 415551 142762
rect 395337 142704 395342 142760
rect 395398 142704 412638 142760
rect 412694 142704 415490 142760
rect 415546 142704 415551 142760
rect 395337 142702 415551 142704
rect 395337 142699 395403 142702
rect 412633 142699 412699 142702
rect 415485 142699 415551 142702
rect 213913 142626 213979 142629
rect 258809 142626 258875 142629
rect 213913 142624 217028 142626
rect 213913 142568 213918 142624
rect 213974 142568 217028 142624
rect 213913 142566 217028 142568
rect 258809 142624 268180 142626
rect 258809 142568 258814 142624
rect 258870 142568 268180 142624
rect 258809 142566 268180 142568
rect 213913 142563 213979 142566
rect 258809 142563 258875 142566
rect 231761 142490 231827 142493
rect 244273 142492 244339 142493
rect 244222 142490 244228 142492
rect 228988 142488 231827 142490
rect 228988 142432 231766 142488
rect 231822 142432 231827 142488
rect 228988 142430 231827 142432
rect 244182 142430 244228 142490
rect 244292 142488 244339 142492
rect 244334 142432 244339 142488
rect 231761 142427 231827 142430
rect 244222 142428 244228 142430
rect 244292 142428 244339 142432
rect 244273 142427 244339 142428
rect 399477 142354 399543 142357
rect 405733 142354 405799 142357
rect 399477 142352 405799 142354
rect 399477 142296 399482 142352
rect 399538 142296 405738 142352
rect 405794 142296 405799 142352
rect 399477 142294 405799 142296
rect 399477 142291 399543 142294
rect 405733 142291 405799 142294
rect 264973 142218 265039 142221
rect 349797 142218 349863 142221
rect 416129 142218 416195 142221
rect 264973 142216 268180 142218
rect 264973 142160 264978 142216
rect 265034 142160 268180 142216
rect 264973 142158 268180 142160
rect 349797 142216 416195 142218
rect 349797 142160 349802 142216
rect 349858 142160 416134 142216
rect 416190 142160 416195 142216
rect 349797 142158 416195 142160
rect 264973 142155 265039 142158
rect 349797 142155 349863 142158
rect 416129 142155 416195 142158
rect 424174 142156 424180 142220
rect 424244 142218 424250 142220
rect 427077 142218 427143 142221
rect 424244 142216 427143 142218
rect 424244 142160 427082 142216
rect 427138 142160 427143 142216
rect 424244 142158 427143 142160
rect 424244 142156 424250 142158
rect 427077 142155 427143 142158
rect 232078 142082 232084 142084
rect 228988 142022 232084 142082
rect 232078 142020 232084 142022
rect 232148 142020 232154 142084
rect 282821 142082 282887 142085
rect 279956 142080 282887 142082
rect 279956 142024 282826 142080
rect 282882 142024 282887 142080
rect 279956 142022 282887 142024
rect 282821 142019 282887 142022
rect 214005 141946 214071 141949
rect 214005 141944 217028 141946
rect 214005 141888 214010 141944
rect 214066 141888 217028 141944
rect 214005 141886 217028 141888
rect 214005 141883 214071 141886
rect 231209 141674 231275 141677
rect 228988 141672 231275 141674
rect 228988 141616 231214 141672
rect 231270 141616 231275 141672
rect 228988 141614 231275 141616
rect 231209 141611 231275 141614
rect 237966 141340 237972 141404
rect 238036 141402 238042 141404
rect 268150 141402 268210 141780
rect 238036 141342 268210 141402
rect 238036 141340 238042 141342
rect 213913 141266 213979 141269
rect 265249 141266 265315 141269
rect 281901 141266 281967 141269
rect 213913 141264 217028 141266
rect 213913 141208 213918 141264
rect 213974 141208 217028 141264
rect 213913 141206 217028 141208
rect 265249 141264 268180 141266
rect 265249 141208 265254 141264
rect 265310 141208 268180 141264
rect 265249 141206 268180 141208
rect 279956 141264 281967 141266
rect 279956 141208 281906 141264
rect 281962 141208 281967 141264
rect 279956 141206 281967 141208
rect 213913 141203 213979 141206
rect 265249 141203 265315 141206
rect 281901 141203 281967 141206
rect 236494 141130 236500 141132
rect 228988 141070 236500 141130
rect 236494 141068 236500 141070
rect 236564 141068 236570 141132
rect 261661 140858 261727 140861
rect 432597 140858 432663 140861
rect 440182 140858 440188 140860
rect 261661 140856 268180 140858
rect 261661 140800 261666 140856
rect 261722 140800 268180 140856
rect 261661 140798 268180 140800
rect 432597 140856 440188 140858
rect 432597 140800 432602 140856
rect 432658 140800 440188 140856
rect 432597 140798 440188 140800
rect 261661 140795 261727 140798
rect 432597 140795 432663 140798
rect 440182 140796 440188 140798
rect 440252 140796 440258 140860
rect 243537 140722 243603 140725
rect 228988 140720 243603 140722
rect 228988 140664 243542 140720
rect 243598 140664 243603 140720
rect 228988 140662 243603 140664
rect 243537 140659 243603 140662
rect 389173 140722 389239 140725
rect 389173 140720 400138 140722
rect 389173 140664 389178 140720
rect 389234 140664 400138 140720
rect 389173 140662 400138 140664
rect 389173 140659 389239 140662
rect 213913 140586 213979 140589
rect 213913 140584 217028 140586
rect 213913 140528 213918 140584
rect 213974 140528 217028 140584
rect 213913 140526 217028 140528
rect 213913 140523 213979 140526
rect 282821 140450 282887 140453
rect 279956 140448 282887 140450
rect 230565 140178 230631 140181
rect 228988 140176 230631 140178
rect 228988 140120 230570 140176
rect 230626 140120 230631 140176
rect 228988 140118 230631 140120
rect 230565 140115 230631 140118
rect 242014 140116 242020 140180
rect 242084 140178 242090 140180
rect 268150 140178 268210 140420
rect 279956 140392 282826 140448
rect 282882 140392 282887 140448
rect 279956 140390 282887 140392
rect 282821 140387 282887 140390
rect 242084 140118 268210 140178
rect 242084 140116 242090 140118
rect 264973 140042 265039 140045
rect 342989 140042 343055 140045
rect 389173 140042 389239 140045
rect 264973 140040 268180 140042
rect 264973 139984 264978 140040
rect 265034 139984 268180 140040
rect 264973 139982 268180 139984
rect 342989 140040 389239 140042
rect 342989 139984 342994 140040
rect 343050 139984 389178 140040
rect 389234 139984 389239 140040
rect 342989 139982 389239 139984
rect 264973 139979 265039 139982
rect 342989 139979 343055 139982
rect 389173 139979 389239 139982
rect 214557 139906 214623 139909
rect 214557 139904 217028 139906
rect 214557 139848 214562 139904
rect 214618 139848 217028 139904
rect 214557 139846 217028 139848
rect 214557 139843 214623 139846
rect 253933 139770 253999 139773
rect 282729 139770 282795 139773
rect 228988 139768 253999 139770
rect 228988 139712 253938 139768
rect 253994 139712 253999 139768
rect 228988 139710 253999 139712
rect 279956 139768 282795 139770
rect 279956 139712 282734 139768
rect 282790 139712 282795 139768
rect 279956 139710 282795 139712
rect 253933 139707 253999 139710
rect 282729 139707 282795 139710
rect 265801 139634 265867 139637
rect 265801 139632 268180 139634
rect 265801 139576 265806 139632
rect 265862 139576 268180 139632
rect 400078 139604 400138 140662
rect 407941 140042 408007 140045
rect 441654 140042 441660 140044
rect 407941 140040 441660 140042
rect 407941 139984 407946 140040
rect 408002 139984 441660 140040
rect 407941 139982 441660 139984
rect 407941 139979 408007 139982
rect 441654 139980 441660 139982
rect 441724 139980 441730 140044
rect 265801 139574 268180 139576
rect 265801 139571 265867 139574
rect 419625 139498 419691 139501
rect 425513 139500 425579 139501
rect 420862 139498 420868 139500
rect 419625 139496 420868 139498
rect 419625 139440 419630 139496
rect 419686 139440 420868 139496
rect 419625 139438 420868 139440
rect 419625 139435 419691 139438
rect 420862 139436 420868 139438
rect 420932 139436 420938 139500
rect 425462 139436 425468 139500
rect 425532 139498 425579 139500
rect 425532 139496 425624 139498
rect 425574 139440 425624 139496
rect 425532 139438 425624 139440
rect 425532 139436 425579 139438
rect 426382 139436 426388 139500
rect 426452 139498 426458 139500
rect 427445 139498 427511 139501
rect 426452 139496 427511 139498
rect 426452 139440 427450 139496
rect 427506 139440 427511 139496
rect 426452 139438 427511 139440
rect 426452 139436 426458 139438
rect 425513 139435 425579 139436
rect 427445 139435 427511 139438
rect 430614 139436 430620 139500
rect 430684 139498 430690 139500
rect 431309 139498 431375 139501
rect 430684 139496 431375 139498
rect 430684 139440 431314 139496
rect 431370 139440 431375 139496
rect 430684 139438 431375 139440
rect 430684 139436 430690 139438
rect 431309 139435 431375 139438
rect 436369 139498 436435 139501
rect 436686 139498 436692 139500
rect 436369 139496 436692 139498
rect 436369 139440 436374 139496
rect 436430 139440 436692 139496
rect 436369 139438 436692 139440
rect 436369 139435 436435 139438
rect 436686 139436 436692 139438
rect 436756 139436 436762 139500
rect 438853 139362 438919 139365
rect 439078 139362 439084 139364
rect 438853 139360 439084 139362
rect 438853 139304 438858 139360
rect 438914 139304 439084 139360
rect 438853 139302 439084 139304
rect 438853 139299 438919 139302
rect 439078 139300 439084 139302
rect 439148 139300 439154 139364
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 213913 139226 213979 139229
rect 233366 139226 233372 139228
rect 213913 139224 217028 139226
rect 213913 139168 213918 139224
rect 213974 139168 217028 139224
rect 213913 139166 217028 139168
rect 228988 139166 233372 139226
rect 213913 139163 213979 139166
rect 233366 139164 233372 139166
rect 233436 139164 233442 139228
rect 265065 139226 265131 139229
rect 265065 139224 268180 139226
rect 265065 139168 265070 139224
rect 265126 139168 268180 139224
rect 583520 139212 584960 139302
rect 265065 139166 268180 139168
rect 265065 139163 265131 139166
rect 282821 138954 282887 138957
rect 441889 138954 441955 138957
rect 442022 138954 442028 138956
rect 279956 138952 282887 138954
rect 279956 138896 282826 138952
rect 282882 138896 282887 138952
rect 279956 138894 282887 138896
rect 439852 138952 442028 138954
rect 439852 138896 441894 138952
rect 441950 138896 442028 138952
rect 439852 138894 442028 138896
rect 282821 138891 282887 138894
rect 441889 138891 441955 138894
rect 442022 138892 442028 138894
rect 442092 138892 442098 138956
rect 245653 138818 245719 138821
rect 393405 138818 393471 138821
rect 228988 138816 245719 138818
rect 228988 138760 245658 138816
rect 245714 138760 245719 138816
rect 228988 138758 245719 138760
rect 245653 138755 245719 138758
rect 393270 138816 400108 138818
rect 393270 138760 393410 138816
rect 393466 138760 400108 138816
rect 393270 138758 400108 138760
rect 214097 138682 214163 138685
rect 383009 138682 383075 138685
rect 393270 138682 393330 138758
rect 393405 138755 393471 138758
rect 214097 138680 217028 138682
rect 214097 138624 214102 138680
rect 214158 138624 217028 138680
rect 383009 138680 393330 138682
rect 214097 138622 217028 138624
rect 214097 138619 214163 138622
rect 236637 138410 236703 138413
rect 268150 138410 268210 138652
rect 383009 138624 383014 138680
rect 383070 138624 393330 138680
rect 383009 138622 393330 138624
rect 383009 138619 383075 138622
rect 439589 138546 439655 138549
rect 439589 138544 439698 138546
rect 439589 138488 439594 138544
rect 439650 138488 439698 138544
rect 439589 138483 439698 138488
rect 236637 138408 268210 138410
rect 236637 138352 236642 138408
rect 236698 138352 268210 138408
rect 236637 138350 268210 138352
rect 236637 138347 236703 138350
rect 231761 138274 231827 138277
rect 228988 138272 231827 138274
rect 228988 138216 231766 138272
rect 231822 138216 231827 138272
rect 228988 138214 231827 138216
rect 231761 138211 231827 138214
rect 264973 138274 265039 138277
rect 282821 138274 282887 138277
rect 264973 138272 268180 138274
rect 264973 138216 264978 138272
rect 265034 138216 268180 138272
rect 264973 138214 268180 138216
rect 279956 138272 282887 138274
rect 279956 138216 282826 138272
rect 282882 138216 282887 138272
rect 279956 138214 282887 138216
rect 264973 138211 265039 138214
rect 282821 138211 282887 138214
rect 439638 138138 439698 138483
rect 441981 138138 442047 138141
rect 439638 138136 442047 138138
rect 439638 138108 441986 138136
rect 439668 138080 441986 138108
rect 442042 138080 442047 138136
rect 439668 138078 442047 138080
rect 441981 138075 442047 138078
rect 213361 138002 213427 138005
rect 213361 138000 217028 138002
rect 213361 137944 213366 138000
rect 213422 137944 217028 138000
rect 213361 137942 217028 137944
rect 213361 137939 213427 137942
rect 245694 137866 245700 137868
rect 228988 137806 245700 137866
rect 245694 137804 245700 137806
rect 245764 137804 245770 137868
rect 264973 137866 265039 137869
rect 264973 137864 268180 137866
rect 264973 137808 264978 137864
rect 265034 137808 268180 137864
rect 264973 137806 268180 137808
rect 264973 137803 265039 137806
rect 358077 137730 358143 137733
rect 399845 137730 399911 137733
rect 358077 137728 399911 137730
rect 358077 137672 358082 137728
rect 358138 137672 399850 137728
rect 399906 137672 399911 137728
rect 358077 137670 399911 137672
rect 358077 137667 358143 137670
rect 399845 137667 399911 137670
rect 397545 137594 397611 137597
rect 397545 137592 400108 137594
rect 397545 137536 397550 137592
rect 397606 137536 400108 137592
rect 397545 137534 400108 137536
rect 397545 137531 397611 137534
rect 176009 137458 176075 137461
rect 216806 137458 216812 137460
rect 176009 137456 216812 137458
rect 176009 137400 176014 137456
rect 176070 137400 216812 137456
rect 176009 137398 216812 137400
rect 176009 137395 176075 137398
rect 216806 137396 216812 137398
rect 216876 137396 216882 137460
rect 281625 137458 281691 137461
rect 440417 137458 440483 137461
rect 279956 137456 281691 137458
rect 229686 137322 229692 137324
rect -960 136778 480 136868
rect 3325 136778 3391 136781
rect -960 136776 3391 136778
rect -960 136720 3330 136776
rect 3386 136720 3391 136776
rect -960 136718 3391 136720
rect -960 136628 480 136718
rect 3325 136715 3391 136718
rect 206369 136778 206435 136781
rect 216998 136778 217058 137292
rect 228988 137262 229692 137322
rect 229686 137260 229692 137262
rect 229756 137260 229762 137324
rect 246573 137186 246639 137189
rect 268150 137186 268210 137428
rect 279956 137400 281630 137456
rect 281686 137400 281691 137456
rect 279956 137398 281691 137400
rect 439852 137456 440483 137458
rect 439852 137400 440422 137456
rect 440478 137400 440483 137456
rect 439852 137398 440483 137400
rect 281625 137395 281691 137398
rect 440417 137395 440483 137398
rect 246573 137184 268210 137186
rect 246573 137128 246578 137184
rect 246634 137128 268210 137184
rect 246573 137126 268210 137128
rect 246573 137123 246639 137126
rect 235257 137050 235323 137053
rect 235257 137048 268180 137050
rect 235257 136992 235262 137048
rect 235318 136992 268180 137048
rect 235257 136990 268180 136992
rect 235257 136987 235323 136990
rect 231577 136914 231643 136917
rect 228988 136912 231643 136914
rect 228988 136856 231582 136912
rect 231638 136856 231643 136912
rect 228988 136854 231643 136856
rect 231577 136851 231643 136854
rect 279325 136914 279391 136917
rect 279325 136912 279434 136914
rect 279325 136856 279330 136912
rect 279386 136856 279434 136912
rect 279325 136851 279434 136856
rect 206369 136776 217058 136778
rect 206369 136720 206374 136776
rect 206430 136720 217058 136776
rect 206369 136718 217058 136720
rect 206369 136715 206435 136718
rect 215937 136642 216003 136645
rect 265065 136642 265131 136645
rect 215937 136640 217028 136642
rect 215937 136584 215942 136640
rect 215998 136584 217028 136640
rect 215937 136582 217028 136584
rect 265065 136640 268180 136642
rect 265065 136584 265070 136640
rect 265126 136584 268180 136640
rect 279374 136612 279434 136851
rect 397545 136778 397611 136781
rect 442901 136778 442967 136781
rect 397545 136776 400108 136778
rect 397545 136720 397550 136776
rect 397606 136720 400108 136776
rect 397545 136718 400108 136720
rect 439852 136776 442967 136778
rect 439852 136720 442906 136776
rect 442962 136720 442967 136776
rect 439852 136718 442967 136720
rect 397545 136715 397611 136718
rect 442901 136715 442967 136718
rect 265065 136582 268180 136584
rect 215937 136579 216003 136582
rect 265065 136579 265131 136582
rect 231761 136370 231827 136373
rect 228988 136368 231827 136370
rect 228988 136312 231766 136368
rect 231822 136312 231827 136368
rect 228988 136310 231827 136312
rect 231761 136307 231827 136310
rect 214005 135962 214071 135965
rect 231301 135962 231367 135965
rect 214005 135960 217028 135962
rect 214005 135904 214010 135960
rect 214066 135904 217028 135960
rect 214005 135902 217028 135904
rect 228988 135960 231367 135962
rect 228988 135904 231306 135960
rect 231362 135904 231367 135960
rect 228988 135902 231367 135904
rect 214005 135899 214071 135902
rect 231301 135899 231367 135902
rect 233734 135764 233740 135828
rect 233804 135826 233810 135828
rect 268150 135826 268210 136204
rect 398598 136172 398604 136236
rect 398668 136234 398674 136236
rect 441705 136234 441771 136237
rect 398668 136174 400108 136234
rect 439852 136232 441771 136234
rect 439852 136176 441710 136232
rect 441766 136176 441771 136232
rect 439852 136174 441771 136176
rect 398668 136172 398674 136174
rect 441705 136171 441771 136174
rect 282269 135962 282335 135965
rect 279956 135960 282335 135962
rect 279956 135904 282274 135960
rect 282330 135904 282335 135960
rect 279956 135902 282335 135904
rect 282269 135899 282335 135902
rect 305494 135900 305500 135964
rect 305564 135962 305570 135964
rect 327073 135962 327139 135965
rect 328361 135962 328427 135965
rect 305564 135960 328427 135962
rect 305564 135904 327078 135960
rect 327134 135904 328366 135960
rect 328422 135904 328427 135960
rect 305564 135902 328427 135904
rect 305564 135900 305570 135902
rect 327073 135899 327139 135902
rect 328361 135899 328427 135902
rect 439497 135826 439563 135829
rect 233804 135766 268210 135826
rect 439454 135824 439563 135826
rect 439454 135768 439502 135824
rect 439558 135768 439563 135824
rect 233804 135764 233810 135766
rect 439454 135763 439563 135768
rect 264973 135690 265039 135693
rect 264973 135688 268180 135690
rect 264973 135632 264978 135688
rect 265034 135632 268180 135688
rect 264973 135630 268180 135632
rect 264973 135627 265039 135630
rect 397637 135554 397703 135557
rect 397637 135552 400108 135554
rect 397637 135496 397642 135552
rect 397698 135496 400108 135552
rect 439454 135524 439514 135763
rect 397637 135494 400108 135496
rect 397637 135491 397703 135494
rect 231485 135418 231551 135421
rect 228988 135416 231551 135418
rect 228988 135360 231490 135416
rect 231546 135360 231551 135416
rect 228988 135358 231551 135360
rect 231485 135355 231551 135358
rect 213913 135282 213979 135285
rect 265065 135282 265131 135285
rect 213913 135280 217028 135282
rect 213913 135224 213918 135280
rect 213974 135224 217028 135280
rect 213913 135222 217028 135224
rect 265065 135280 268180 135282
rect 265065 135224 265070 135280
rect 265126 135224 268180 135280
rect 265065 135222 268180 135224
rect 213913 135219 213979 135222
rect 265065 135219 265131 135222
rect 231761 135146 231827 135149
rect 264237 135146 264303 135149
rect 284334 135146 284340 135148
rect 231761 135144 264303 135146
rect 231761 135088 231766 135144
rect 231822 135088 264242 135144
rect 264298 135088 264303 135144
rect 231761 135086 264303 135088
rect 279956 135086 284340 135146
rect 231761 135083 231827 135086
rect 264237 135083 264303 135086
rect 284334 135084 284340 135086
rect 284404 135084 284410 135148
rect 231158 135010 231164 135012
rect 228988 134950 231164 135010
rect 231158 134948 231164 134950
rect 231228 134948 231234 135012
rect 265157 134874 265223 134877
rect 398649 134874 398715 134877
rect 442901 134874 442967 134877
rect 265157 134872 268180 134874
rect 265157 134816 265162 134872
rect 265218 134816 268180 134872
rect 265157 134814 268180 134816
rect 398649 134872 400108 134874
rect 398649 134816 398654 134872
rect 398710 134816 400108 134872
rect 398649 134814 400108 134816
rect 439852 134872 442967 134874
rect 439852 134816 442906 134872
rect 442962 134816 442967 134872
rect 439852 134814 442967 134816
rect 265157 134811 265223 134814
rect 398649 134811 398715 134814
rect 442901 134811 442967 134814
rect 213913 134602 213979 134605
rect 213913 134600 217028 134602
rect 213913 134544 213918 134600
rect 213974 134544 217028 134600
rect 213913 134542 217028 134544
rect 213913 134539 213979 134542
rect 231761 134466 231827 134469
rect 228988 134464 231827 134466
rect 228988 134408 231766 134464
rect 231822 134408 231827 134464
rect 228988 134406 231827 134408
rect 231761 134403 231827 134406
rect 249190 134404 249196 134468
rect 249260 134466 249266 134468
rect 265065 134466 265131 134469
rect 284518 134466 284524 134468
rect 249260 134464 265131 134466
rect 249260 134408 265070 134464
rect 265126 134408 265131 134464
rect 249260 134406 265131 134408
rect 249260 134404 249266 134406
rect 265065 134403 265131 134406
rect 265617 134194 265683 134197
rect 268150 134194 268210 134436
rect 279956 134406 284524 134466
rect 284518 134404 284524 134406
rect 284588 134404 284594 134468
rect 265617 134192 268210 134194
rect 265617 134136 265622 134192
rect 265678 134136 268210 134192
rect 265617 134134 268210 134136
rect 265617 134131 265683 134134
rect 231485 134058 231551 134061
rect 228988 134056 231551 134058
rect 228988 134000 231490 134056
rect 231546 134000 231551 134056
rect 228988 133998 231551 134000
rect 231485 133995 231551 133998
rect 264973 134058 265039 134061
rect 397545 134058 397611 134061
rect 264973 134056 268180 134058
rect 264973 134000 264978 134056
rect 265034 134000 268180 134056
rect 264973 133998 268180 134000
rect 397545 134056 400108 134058
rect 397545 134000 397550 134056
rect 397606 134000 400108 134056
rect 397545 133998 400108 134000
rect 264973 133995 265039 133998
rect 397545 133995 397611 133998
rect 216121 133922 216187 133925
rect 216121 133920 217028 133922
rect 216121 133864 216126 133920
rect 216182 133864 217028 133920
rect 216121 133862 217028 133864
rect 216121 133859 216187 133862
rect 264973 133650 265039 133653
rect 285622 133650 285628 133652
rect 264973 133648 268180 133650
rect 264973 133592 264978 133648
rect 265034 133592 268180 133648
rect 264973 133590 268180 133592
rect 279956 133590 285628 133650
rect 264973 133587 265039 133590
rect 285622 133588 285628 133590
rect 285692 133588 285698 133652
rect 231761 133514 231827 133517
rect 228988 133512 231827 133514
rect 228988 133456 231766 133512
rect 231822 133456 231827 133512
rect 228988 133454 231827 133456
rect 231761 133451 231827 133454
rect 397637 133514 397703 133517
rect 442901 133514 442967 133517
rect 397637 133512 400108 133514
rect 397637 133456 397642 133512
rect 397698 133456 400108 133512
rect 397637 133454 400108 133456
rect 439852 133512 442967 133514
rect 439852 133456 442906 133512
rect 442962 133456 442967 133512
rect 439852 133454 442967 133456
rect 397637 133451 397703 133454
rect 442901 133451 442967 133454
rect 213913 133378 213979 133381
rect 213913 133376 217028 133378
rect 213913 133320 213918 133376
rect 213974 133320 217028 133376
rect 213913 133318 217028 133320
rect 213913 133315 213979 133318
rect 231209 133106 231275 133109
rect 228988 133104 231275 133106
rect 228988 133048 231214 133104
rect 231270 133048 231275 133104
rect 228988 133046 231275 133048
rect 231209 133043 231275 133046
rect 246389 132834 246455 132837
rect 268150 132834 268210 133076
rect 282821 132834 282887 132837
rect 440233 132834 440299 132837
rect 246389 132832 268210 132834
rect 246389 132776 246394 132832
rect 246450 132776 268210 132832
rect 246389 132774 268210 132776
rect 279956 132832 282887 132834
rect 279956 132776 282826 132832
rect 282882 132776 282887 132832
rect 279956 132774 282887 132776
rect 439852 132832 440299 132834
rect 439852 132776 440238 132832
rect 440294 132776 440299 132832
rect 439852 132774 440299 132776
rect 246389 132771 246455 132774
rect 282821 132771 282887 132774
rect 440233 132771 440299 132774
rect 214465 132698 214531 132701
rect 214465 132696 217028 132698
rect 214465 132640 214470 132696
rect 214526 132640 217028 132696
rect 214465 132638 217028 132640
rect 214465 132635 214531 132638
rect 258574 132636 258580 132700
rect 258644 132698 258650 132700
rect 258644 132638 268180 132698
rect 258644 132636 258650 132638
rect 231669 132562 231735 132565
rect 228988 132560 231735 132562
rect 228988 132504 231674 132560
rect 231730 132504 231735 132560
rect 228988 132502 231735 132504
rect 231669 132499 231735 132502
rect 258717 132426 258783 132429
rect 238710 132424 258783 132426
rect 238710 132368 258722 132424
rect 258778 132368 258783 132424
rect 238710 132366 258783 132368
rect 238710 132154 238770 132366
rect 258717 132363 258783 132366
rect 378869 132426 378935 132429
rect 390553 132426 390619 132429
rect 378869 132424 390619 132426
rect 378869 132368 378874 132424
rect 378930 132368 390558 132424
rect 390614 132368 390619 132424
rect 378869 132366 390619 132368
rect 378869 132363 378935 132366
rect 390553 132363 390619 132366
rect 228988 132094 238770 132154
rect 213913 132018 213979 132021
rect 268150 132018 268210 132260
rect 281717 132154 281783 132157
rect 279956 132152 281783 132154
rect 279956 132096 281722 132152
rect 281778 132096 281783 132152
rect 279956 132094 281783 132096
rect 281717 132091 281783 132094
rect 397545 132154 397611 132157
rect 441797 132154 441863 132157
rect 397545 132152 400108 132154
rect 397545 132096 397550 132152
rect 397606 132096 400108 132152
rect 397545 132094 400108 132096
rect 439852 132152 441863 132154
rect 439852 132096 441802 132152
rect 441858 132096 441863 132152
rect 439852 132094 441863 132096
rect 397545 132091 397611 132094
rect 441797 132091 441863 132094
rect 213913 132016 217028 132018
rect 213913 131960 213918 132016
rect 213974 131960 217028 132016
rect 213913 131958 217028 131960
rect 258030 131958 268210 132018
rect 213913 131955 213979 131958
rect 231761 131610 231827 131613
rect 258030 131610 258090 131958
rect 264973 131882 265039 131885
rect 264973 131880 268180 131882
rect 264973 131824 264978 131880
rect 265034 131824 268180 131880
rect 264973 131822 268180 131824
rect 264973 131819 265039 131822
rect 439405 131746 439471 131749
rect 439405 131744 439514 131746
rect 439405 131688 439410 131744
rect 439466 131688 439514 131744
rect 439405 131683 439514 131688
rect 228988 131608 231827 131610
rect 228988 131552 231766 131608
rect 231822 131552 231827 131608
rect 228988 131550 231827 131552
rect 231761 131547 231827 131550
rect 238710 131550 258090 131610
rect 229686 131412 229692 131476
rect 229756 131474 229762 131476
rect 238710 131474 238770 131550
rect 229756 131414 238770 131474
rect 267089 131474 267155 131477
rect 267089 131472 268180 131474
rect 267089 131416 267094 131472
rect 267150 131416 268180 131472
rect 439454 131444 439514 131683
rect 267089 131414 268180 131416
rect 229756 131412 229762 131414
rect 267089 131411 267155 131414
rect 210509 131338 210575 131341
rect 282637 131338 282703 131341
rect 393405 131338 393471 131341
rect 210509 131336 217028 131338
rect 210509 131280 210514 131336
rect 210570 131280 217028 131336
rect 210509 131278 217028 131280
rect 279956 131336 282703 131338
rect 279956 131280 282642 131336
rect 282698 131280 282703 131336
rect 279956 131278 282703 131280
rect 210509 131275 210575 131278
rect 282637 131275 282703 131278
rect 393270 131336 400108 131338
rect 393270 131280 393410 131336
rect 393466 131280 400108 131336
rect 393270 131278 400108 131280
rect 231117 131202 231183 131205
rect 228988 131200 231183 131202
rect 228988 131144 231122 131200
rect 231178 131144 231183 131200
rect 228988 131142 231183 131144
rect 231117 131139 231183 131142
rect 390553 131202 390619 131205
rect 393270 131202 393330 131278
rect 393405 131275 393471 131278
rect 390553 131200 393330 131202
rect 390553 131144 390558 131200
rect 390614 131144 393330 131200
rect 390553 131142 393330 131144
rect 390553 131139 390619 131142
rect 264973 131066 265039 131069
rect 264973 131064 268180 131066
rect 264973 131008 264978 131064
rect 265034 131008 268180 131064
rect 264973 131006 268180 131008
rect 264973 131003 265039 131006
rect 442901 130794 442967 130797
rect 439852 130792 442967 130794
rect 439852 130736 442906 130792
rect 442962 130736 442967 130792
rect 439852 130734 442967 130736
rect 442901 130731 442967 130734
rect 213913 130658 213979 130661
rect 231761 130658 231827 130661
rect 282269 130658 282335 130661
rect 213913 130656 217028 130658
rect 213913 130600 213918 130656
rect 213974 130600 217028 130656
rect 213913 130598 217028 130600
rect 228988 130656 231827 130658
rect 228988 130600 231766 130656
rect 231822 130600 231827 130656
rect 228988 130598 231827 130600
rect 279956 130656 282335 130658
rect 279956 130600 282274 130656
rect 282330 130600 282335 130656
rect 279956 130598 282335 130600
rect 213913 130595 213979 130598
rect 231761 130595 231827 130598
rect 282269 130595 282335 130598
rect 397545 130658 397611 130661
rect 397545 130656 400108 130658
rect 397545 130600 397550 130656
rect 397606 130600 400108 130656
rect 397545 130598 400108 130600
rect 397545 130595 397611 130598
rect 231393 130250 231459 130253
rect 228988 130248 231459 130250
rect 228988 130192 231398 130248
rect 231454 130192 231459 130248
rect 228988 130190 231459 130192
rect 231393 130187 231459 130190
rect 258901 130250 258967 130253
rect 268150 130250 268210 130492
rect 282729 130386 282795 130389
rect 313273 130386 313339 130389
rect 282729 130384 313339 130386
rect 282729 130328 282734 130384
rect 282790 130328 313278 130384
rect 313334 130328 313339 130384
rect 282729 130326 313339 130328
rect 282729 130323 282795 130326
rect 313273 130323 313339 130326
rect 258901 130248 268210 130250
rect 258901 130192 258906 130248
rect 258962 130192 268210 130248
rect 258901 130190 268210 130192
rect 258901 130187 258967 130190
rect 249006 130052 249012 130116
rect 249076 130114 249082 130116
rect 249076 130054 268180 130114
rect 249076 130052 249082 130054
rect 214005 129978 214071 129981
rect 389909 129978 389975 129981
rect 442901 129978 442967 129981
rect 214005 129976 217028 129978
rect 214005 129920 214010 129976
rect 214066 129920 217028 129976
rect 214005 129918 217028 129920
rect 389909 129976 400108 129978
rect 389909 129920 389914 129976
rect 389970 129920 400108 129976
rect 389909 129918 400108 129920
rect 439852 129976 442967 129978
rect 439852 129920 442906 129976
rect 442962 129920 442967 129976
rect 439852 129918 442967 129920
rect 214005 129915 214071 129918
rect 389909 129915 389975 129918
rect 442901 129915 442967 129918
rect 231301 129842 231367 129845
rect 228988 129840 231367 129842
rect 228988 129784 231306 129840
rect 231362 129784 231367 129840
rect 228988 129782 231367 129784
rect 231301 129779 231367 129782
rect 231485 129842 231551 129845
rect 238385 129842 238451 129845
rect 282821 129842 282887 129845
rect 231485 129840 238451 129842
rect 231485 129784 231490 129840
rect 231546 129784 238390 129840
rect 238446 129784 238451 129840
rect 231485 129782 238451 129784
rect 279956 129840 282887 129842
rect 279956 129784 282826 129840
rect 282882 129784 282887 129840
rect 279956 129782 282887 129784
rect 231485 129779 231551 129782
rect 238385 129779 238451 129782
rect 282821 129779 282887 129782
rect 268150 129434 268210 129676
rect 258030 129374 268210 129434
rect 66161 129298 66227 129301
rect 68142 129298 68816 129304
rect 66161 129296 68816 129298
rect 66161 129240 66166 129296
rect 66222 129244 68816 129296
rect 213913 129298 213979 129301
rect 231761 129298 231827 129301
rect 213913 129296 217028 129298
rect 66222 129240 68202 129244
rect 66161 129238 68202 129240
rect 213913 129240 213918 129296
rect 213974 129240 217028 129296
rect 213913 129238 217028 129240
rect 228988 129296 231827 129298
rect 228988 129240 231766 129296
rect 231822 129240 231827 129296
rect 228988 129238 231827 129240
rect 66161 129235 66227 129238
rect 213913 129235 213979 129238
rect 231761 129235 231827 129238
rect 238201 129026 238267 129029
rect 258030 129026 258090 129374
rect 265065 129298 265131 129301
rect 397545 129298 397611 129301
rect 442165 129298 442231 129301
rect 265065 129296 268180 129298
rect 265065 129240 265070 129296
rect 265126 129240 268180 129296
rect 265065 129238 268180 129240
rect 397545 129296 400108 129298
rect 397545 129240 397550 129296
rect 397606 129240 400108 129296
rect 397545 129238 400108 129240
rect 439852 129296 442231 129298
rect 439852 129240 442170 129296
rect 442226 129240 442231 129296
rect 439852 129238 442231 129240
rect 265065 129235 265131 129238
rect 397545 129235 397611 129238
rect 442165 129235 442231 129238
rect 282085 129026 282151 129029
rect 238201 129024 258090 129026
rect 238201 128968 238206 129024
rect 238262 128968 258090 129024
rect 238201 128966 258090 128968
rect 279956 129024 282151 129026
rect 279956 128968 282090 129024
rect 282146 128968 282151 129024
rect 279956 128966 282151 128968
rect 238201 128963 238267 128966
rect 282085 128963 282151 128966
rect 231393 128890 231459 128893
rect 228988 128888 231459 128890
rect 228988 128832 231398 128888
rect 231454 128832 231459 128888
rect 228988 128830 231459 128832
rect 231393 128827 231459 128830
rect 264973 128890 265039 128893
rect 264973 128888 268180 128890
rect 264973 128832 264978 128888
rect 265034 128832 268180 128888
rect 264973 128830 268180 128832
rect 264973 128827 265039 128830
rect 214097 128754 214163 128757
rect 394601 128754 394667 128757
rect 214097 128752 217028 128754
rect 214097 128696 214102 128752
rect 214158 128696 217028 128752
rect 214097 128694 217028 128696
rect 394601 128752 400108 128754
rect 394601 128696 394606 128752
rect 394662 128696 400108 128752
rect 394601 128694 400108 128696
rect 214097 128691 214163 128694
rect 394601 128691 394667 128694
rect 267590 128420 267596 128484
rect 267660 128482 267666 128484
rect 267660 128422 268180 128482
rect 267660 128420 267666 128422
rect 231761 128346 231827 128349
rect 280889 128346 280955 128349
rect 228988 128344 231827 128346
rect 228988 128288 231766 128344
rect 231822 128288 231827 128344
rect 228988 128286 231827 128288
rect 279956 128344 280955 128346
rect 279956 128288 280894 128344
rect 280950 128288 280955 128344
rect 279956 128286 280955 128288
rect 231761 128283 231827 128286
rect 280889 128283 280955 128286
rect 66161 128074 66227 128077
rect 68142 128074 68816 128080
rect 66161 128072 68816 128074
rect 66161 128016 66166 128072
rect 66222 128020 68816 128072
rect 213913 128074 213979 128077
rect 213913 128072 217028 128074
rect 66222 128016 68202 128020
rect 66161 128014 68202 128016
rect 213913 128016 213918 128072
rect 213974 128016 217028 128072
rect 213913 128014 217028 128016
rect 66161 128011 66227 128014
rect 213913 128011 213979 128014
rect 231669 127938 231735 127941
rect 228988 127936 231735 127938
rect 228988 127880 231674 127936
rect 231730 127880 231735 127936
rect 228988 127878 231735 127880
rect 231669 127875 231735 127878
rect 264973 127938 265039 127941
rect 397545 127938 397611 127941
rect 440233 127938 440299 127941
rect 264973 127936 268180 127938
rect 264973 127880 264978 127936
rect 265034 127880 268180 127936
rect 264973 127878 268180 127880
rect 397545 127936 400108 127938
rect 397545 127880 397550 127936
rect 397606 127880 400108 127936
rect 397545 127878 400108 127880
rect 439852 127936 440299 127938
rect 439852 127880 440238 127936
rect 440294 127880 440299 127936
rect 439852 127878 440299 127880
rect 264973 127875 265039 127878
rect 397545 127875 397611 127878
rect 440233 127875 440299 127878
rect 231577 127666 231643 127669
rect 257337 127666 257403 127669
rect 231577 127664 257403 127666
rect 231577 127608 231582 127664
rect 231638 127608 257342 127664
rect 257398 127608 257403 127664
rect 231577 127606 257403 127608
rect 231577 127603 231643 127606
rect 257337 127603 257403 127606
rect 265065 127530 265131 127533
rect 282177 127530 282243 127533
rect 265065 127528 268180 127530
rect 265065 127472 265070 127528
rect 265126 127472 268180 127528
rect 265065 127470 268180 127472
rect 279956 127528 282243 127530
rect 279956 127472 282182 127528
rect 282238 127472 282243 127528
rect 279956 127470 282243 127472
rect 265065 127467 265131 127470
rect 282177 127467 282243 127470
rect 231301 127394 231367 127397
rect 228988 127392 231367 127394
rect 203609 127258 203675 127261
rect 216998 127258 217058 127364
rect 228988 127336 231306 127392
rect 231362 127336 231367 127392
rect 228988 127334 231367 127336
rect 231301 127331 231367 127334
rect 442901 127258 442967 127261
rect 203609 127256 217058 127258
rect 203609 127200 203614 127256
rect 203670 127200 217058 127256
rect 203609 127198 217058 127200
rect 439852 127256 442967 127258
rect 439852 127200 442906 127256
rect 442962 127200 442967 127256
rect 439852 127198 442967 127200
rect 203609 127195 203675 127198
rect 442901 127195 442967 127198
rect 64781 127122 64847 127125
rect 66161 127122 66227 127125
rect 64781 127120 66227 127122
rect 64781 127064 64786 127120
rect 64842 127064 66166 127120
rect 66222 127064 66227 127120
rect 64781 127062 66227 127064
rect 64781 127059 64847 127062
rect 66161 127059 66227 127062
rect 262806 127060 262812 127124
rect 262876 127122 262882 127124
rect 262876 127062 268180 127122
rect 262876 127060 262882 127062
rect 231761 126986 231827 126989
rect 228988 126984 231827 126986
rect 228988 126928 231766 126984
rect 231822 126928 231827 126984
rect 228988 126926 231827 126928
rect 231761 126923 231827 126926
rect 281717 126850 281783 126853
rect 279956 126848 281783 126850
rect 279956 126792 281722 126848
rect 281778 126792 281783 126848
rect 279956 126790 281783 126792
rect 281717 126787 281783 126790
rect 214741 126714 214807 126717
rect 398097 126714 398163 126717
rect 398833 126714 398899 126717
rect 442901 126714 442967 126717
rect 214741 126712 217028 126714
rect 214741 126656 214746 126712
rect 214802 126656 217028 126712
rect 398097 126712 400108 126714
rect 214741 126654 217028 126656
rect 214741 126651 214807 126654
rect 231669 126442 231735 126445
rect 268150 126442 268210 126684
rect 398097 126656 398102 126712
rect 398158 126656 398838 126712
rect 398894 126656 400108 126712
rect 398097 126654 400108 126656
rect 439852 126712 442967 126714
rect 439852 126656 442906 126712
rect 442962 126656 442967 126712
rect 439852 126654 442967 126656
rect 398097 126651 398163 126654
rect 398833 126651 398899 126654
rect 442901 126651 442967 126654
rect 228988 126440 231735 126442
rect 228988 126384 231674 126440
rect 231730 126384 231735 126440
rect 228988 126382 231735 126384
rect 231669 126379 231735 126382
rect 258030 126382 268210 126442
rect 66161 126306 66227 126309
rect 68142 126306 68816 126312
rect 66161 126304 68816 126306
rect 66161 126248 66166 126304
rect 66222 126252 68816 126304
rect 66222 126248 68202 126252
rect 66161 126246 68202 126248
rect 66161 126243 66227 126246
rect 213913 126034 213979 126037
rect 230749 126034 230815 126037
rect 213913 126032 217028 126034
rect 213913 125976 213918 126032
rect 213974 125976 217028 126032
rect 213913 125974 217028 125976
rect 228988 126032 230815 126034
rect 228988 125976 230754 126032
rect 230810 125976 230815 126032
rect 228988 125974 230815 125976
rect 213913 125971 213979 125974
rect 230749 125971 230815 125974
rect 254577 126034 254643 126037
rect 258030 126034 258090 126382
rect 265893 126306 265959 126309
rect 340229 126306 340295 126309
rect 371233 126306 371299 126309
rect 265893 126304 268180 126306
rect 265893 126248 265898 126304
rect 265954 126248 268180 126304
rect 265893 126246 268180 126248
rect 340229 126304 371299 126306
rect 340229 126248 340234 126304
rect 340290 126248 371238 126304
rect 371294 126248 371299 126304
rect 340229 126246 371299 126248
rect 265893 126243 265959 126246
rect 340229 126243 340295 126246
rect 371233 126243 371299 126246
rect 282269 126034 282335 126037
rect 254577 126032 258090 126034
rect 254577 125976 254582 126032
rect 254638 125976 258090 126032
rect 254577 125974 258090 125976
rect 279956 126032 282335 126034
rect 279956 125976 282274 126032
rect 282330 125976 282335 126032
rect 279956 125974 282335 125976
rect 254577 125971 254643 125974
rect 282269 125971 282335 125974
rect 396809 126034 396875 126037
rect 442809 126034 442875 126037
rect 396809 126032 400108 126034
rect 396809 125976 396814 126032
rect 396870 125976 400108 126032
rect 396809 125974 400108 125976
rect 439852 126032 442875 126034
rect 439852 125976 442814 126032
rect 442870 125976 442875 126032
rect 439852 125974 442875 125976
rect 396809 125971 396875 125974
rect 442809 125971 442875 125974
rect 580257 126034 580323 126037
rect 583520 126034 584960 126124
rect 580257 126032 584960 126034
rect 580257 125976 580262 126032
rect 580318 125976 584960 126032
rect 580257 125974 584960 125976
rect 580257 125971 580323 125974
rect 264973 125898 265039 125901
rect 264973 125896 268180 125898
rect 264973 125840 264978 125896
rect 265034 125840 268180 125896
rect 583520 125884 584960 125974
rect 264973 125838 268180 125840
rect 264973 125835 265039 125838
rect 232497 125490 232563 125493
rect 228988 125488 232563 125490
rect 228988 125432 232502 125488
rect 232558 125432 232563 125488
rect 228988 125430 232563 125432
rect 232497 125427 232563 125430
rect 301037 125490 301103 125493
rect 301313 125490 301379 125493
rect 360142 125490 360148 125492
rect 301037 125488 360148 125490
rect 301037 125432 301042 125488
rect 301098 125432 301318 125488
rect 301374 125432 360148 125488
rect 301037 125430 360148 125432
rect 301037 125427 301103 125430
rect 301313 125427 301379 125430
rect 360142 125428 360148 125430
rect 360212 125428 360218 125492
rect 213913 125354 213979 125357
rect 231761 125354 231827 125357
rect 239397 125354 239463 125357
rect 213913 125352 217028 125354
rect 213913 125296 213918 125352
rect 213974 125296 217028 125352
rect 213913 125294 217028 125296
rect 231761 125352 239463 125354
rect 231761 125296 231766 125352
rect 231822 125296 239402 125352
rect 239458 125296 239463 125352
rect 231761 125294 239463 125296
rect 213913 125291 213979 125294
rect 231761 125291 231827 125294
rect 239397 125291 239463 125294
rect 267181 125354 267247 125357
rect 267181 125352 268180 125354
rect 267181 125296 267186 125352
rect 267242 125296 268180 125352
rect 267181 125294 268180 125296
rect 267181 125291 267247 125294
rect 67449 125218 67515 125221
rect 68142 125218 68816 125224
rect 282729 125218 282795 125221
rect 67449 125216 68816 125218
rect 67449 125160 67454 125216
rect 67510 125164 68816 125216
rect 279956 125216 282795 125218
rect 67510 125160 68202 125164
rect 67449 125158 68202 125160
rect 279956 125160 282734 125216
rect 282790 125160 282795 125216
rect 279956 125158 282795 125160
rect 67449 125155 67515 125158
rect 282729 125155 282795 125158
rect 397545 125218 397611 125221
rect 443085 125218 443151 125221
rect 397545 125216 400108 125218
rect 397545 125160 397550 125216
rect 397606 125160 400108 125216
rect 397545 125158 400108 125160
rect 439852 125216 443151 125218
rect 439852 125160 443090 125216
rect 443146 125160 443151 125216
rect 439852 125158 443151 125160
rect 397545 125155 397611 125158
rect 443085 125155 443151 125158
rect 230974 125082 230980 125084
rect 228988 125022 230980 125082
rect 230974 125020 230980 125022
rect 231044 125020 231050 125084
rect 239673 124810 239739 124813
rect 250805 124810 250871 124813
rect 239673 124808 250871 124810
rect 239673 124752 239678 124808
rect 239734 124752 250810 124808
rect 250866 124752 250871 124808
rect 239673 124750 250871 124752
rect 239673 124747 239739 124750
rect 250805 124747 250871 124750
rect 215017 124674 215083 124677
rect 247769 124674 247835 124677
rect 268150 124674 268210 124916
rect 282269 124810 282335 124813
rect 301313 124810 301379 124813
rect 282269 124808 301379 124810
rect 282269 124752 282274 124808
rect 282330 124752 301318 124808
rect 301374 124752 301379 124808
rect 282269 124750 301379 124752
rect 282269 124747 282335 124750
rect 301313 124747 301379 124750
rect 215017 124672 217028 124674
rect 215017 124616 215022 124672
rect 215078 124616 217028 124672
rect 215017 124614 217028 124616
rect 247769 124672 268210 124674
rect 247769 124616 247774 124672
rect 247830 124616 268210 124672
rect 247769 124614 268210 124616
rect 398741 124674 398807 124677
rect 442901 124674 442967 124677
rect 398741 124672 400108 124674
rect 398741 124616 398746 124672
rect 398802 124616 400108 124672
rect 398741 124614 400108 124616
rect 439852 124672 442967 124674
rect 439852 124616 442906 124672
rect 442962 124616 442967 124672
rect 439852 124614 442967 124616
rect 215017 124611 215083 124614
rect 247769 124611 247835 124614
rect 398741 124611 398807 124614
rect 442901 124611 442967 124614
rect 231761 124538 231827 124541
rect 228988 124536 231827 124538
rect 228988 124480 231766 124536
rect 231822 124480 231827 124536
rect 228988 124478 231827 124480
rect 231761 124475 231827 124478
rect 264973 124538 265039 124541
rect 282361 124538 282427 124541
rect 264973 124536 268180 124538
rect 264973 124480 264978 124536
rect 265034 124480 268180 124536
rect 264973 124478 268180 124480
rect 279956 124536 282427 124538
rect 279956 124480 282366 124536
rect 282422 124480 282427 124536
rect 279956 124478 282427 124480
rect 264973 124475 265039 124478
rect 282361 124475 282427 124478
rect 214005 124130 214071 124133
rect 231577 124130 231643 124133
rect 214005 124128 217028 124130
rect 214005 124072 214010 124128
rect 214066 124072 217028 124128
rect 214005 124070 217028 124072
rect 228988 124128 231643 124130
rect 228988 124072 231582 124128
rect 231638 124072 231643 124128
rect 228988 124070 231643 124072
rect 214005 124067 214071 124070
rect 231577 124067 231643 124070
rect 265065 124130 265131 124133
rect 352741 124130 352807 124133
rect 353334 124130 353340 124132
rect 265065 124128 268180 124130
rect 265065 124072 265070 124128
rect 265126 124072 268180 124128
rect 265065 124070 268180 124072
rect 352741 124128 353340 124130
rect 352741 124072 352746 124128
rect 352802 124072 353340 124128
rect 352741 124070 353340 124072
rect 265065 124067 265131 124070
rect 352741 124067 352807 124070
rect 353334 124068 353340 124070
rect 353404 124130 353410 124132
rect 354029 124130 354095 124133
rect 353404 124128 354095 124130
rect 353404 124072 354034 124128
rect 354090 124072 354095 124128
rect 353404 124070 354095 124072
rect 353404 124068 353410 124070
rect 354029 124067 354095 124070
rect 441613 123994 441679 123997
rect 442625 123994 442691 123997
rect 439852 123992 442691 123994
rect 439852 123936 441618 123992
rect 441674 123936 442630 123992
rect 442686 123936 442691 123992
rect 439852 123934 442691 123936
rect 441613 123931 441679 123934
rect 442625 123931 442691 123934
rect 397545 123858 397611 123861
rect 397545 123856 400108 123858
rect -960 123572 480 123812
rect 397545 123800 397550 123856
rect 397606 123800 400108 123856
rect 397545 123798 400108 123800
rect 397545 123795 397611 123798
rect 281993 123722 282059 123725
rect 279956 123720 282059 123722
rect 67357 123586 67423 123589
rect 68142 123586 68816 123592
rect 67357 123584 68816 123586
rect 67357 123528 67362 123584
rect 67418 123532 68816 123584
rect 203517 123586 203583 123589
rect 214097 123586 214163 123589
rect 230565 123586 230631 123589
rect 203517 123584 214163 123586
rect 67418 123528 68202 123532
rect 67357 123526 68202 123528
rect 203517 123528 203522 123584
rect 203578 123528 214102 123584
rect 214158 123528 214163 123584
rect 203517 123526 214163 123528
rect 228988 123584 230631 123586
rect 228988 123528 230570 123584
rect 230626 123528 230631 123584
rect 228988 123526 230631 123528
rect 67357 123523 67423 123526
rect 203517 123523 203583 123526
rect 214097 123523 214163 123526
rect 230565 123523 230631 123526
rect 213913 123450 213979 123453
rect 231209 123450 231275 123453
rect 240869 123450 240935 123453
rect 213913 123448 217028 123450
rect 213913 123392 213918 123448
rect 213974 123392 217028 123448
rect 213913 123390 217028 123392
rect 231209 123448 240935 123450
rect 231209 123392 231214 123448
rect 231270 123392 240874 123448
rect 240930 123392 240935 123448
rect 231209 123390 240935 123392
rect 213913 123387 213979 123390
rect 231209 123387 231275 123390
rect 240869 123387 240935 123390
rect 248413 123450 248479 123453
rect 268150 123450 268210 123692
rect 279956 123664 281998 123720
rect 282054 123664 282059 123720
rect 279956 123662 282059 123664
rect 281993 123659 282059 123662
rect 248413 123448 268210 123450
rect 248413 123392 248418 123448
rect 248474 123392 268210 123448
rect 248413 123390 268210 123392
rect 248413 123387 248479 123390
rect 397637 123314 397703 123317
rect 258030 123254 268180 123314
rect 397637 123312 400108 123314
rect 397637 123256 397642 123312
rect 397698 123256 400108 123312
rect 397637 123254 400108 123256
rect 231761 123178 231827 123181
rect 228988 123176 231827 123178
rect 228988 123120 231766 123176
rect 231822 123120 231827 123176
rect 228988 123118 231827 123120
rect 231761 123115 231827 123118
rect 239397 123178 239463 123181
rect 258030 123178 258090 123254
rect 397637 123251 397703 123254
rect 239397 123176 258090 123178
rect 239397 123120 239402 123176
rect 239458 123120 258090 123176
rect 239397 123118 258090 123120
rect 239397 123115 239463 123118
rect 282821 123042 282887 123045
rect 279956 123040 282887 123042
rect 279956 122984 282826 123040
rect 282882 122984 282887 123040
rect 279956 122982 282887 122984
rect 282821 122979 282887 122982
rect 264973 122906 265039 122909
rect 264973 122904 268180 122906
rect 264973 122848 264978 122904
rect 265034 122848 268180 122904
rect 264973 122846 268180 122848
rect 264973 122843 265039 122846
rect 214005 122770 214071 122773
rect 262857 122770 262923 122773
rect 214005 122768 217028 122770
rect 214005 122712 214010 122768
rect 214066 122712 217028 122768
rect 214005 122710 217028 122712
rect 238710 122768 262923 122770
rect 238710 122712 262862 122768
rect 262918 122712 262923 122768
rect 238710 122710 262923 122712
rect 214005 122707 214071 122710
rect 66069 122634 66135 122637
rect 68142 122634 68816 122640
rect 238710 122634 238770 122710
rect 262857 122707 262923 122710
rect 441889 122634 441955 122637
rect 66069 122632 68816 122634
rect 66069 122576 66074 122632
rect 66130 122580 68816 122632
rect 66130 122576 68202 122580
rect 66069 122574 68202 122576
rect 228988 122574 238770 122634
rect 439852 122632 441955 122634
rect 439852 122576 441894 122632
rect 441950 122576 441955 122632
rect 439852 122574 441955 122576
rect 66069 122571 66135 122574
rect 441889 122571 441955 122574
rect 397545 122498 397611 122501
rect 397545 122496 400108 122498
rect 397545 122440 397550 122496
rect 397606 122440 400108 122496
rect 397545 122438 400108 122440
rect 397545 122435 397611 122438
rect 231761 122226 231827 122229
rect 228988 122224 231827 122226
rect 228988 122168 231766 122224
rect 231822 122168 231827 122224
rect 228988 122166 231827 122168
rect 231761 122163 231827 122166
rect 213913 122090 213979 122093
rect 230013 122090 230079 122093
rect 268150 122090 268210 122332
rect 282821 122226 282887 122229
rect 279956 122224 282887 122226
rect 279956 122168 282826 122224
rect 282882 122168 282887 122224
rect 279956 122166 282887 122168
rect 282821 122163 282887 122166
rect 213913 122088 217028 122090
rect 213913 122032 213918 122088
rect 213974 122032 217028 122088
rect 213913 122030 217028 122032
rect 230013 122088 268210 122090
rect 230013 122032 230018 122088
rect 230074 122032 268210 122088
rect 230013 122030 268210 122032
rect 213913 122027 213979 122030
rect 230013 122027 230079 122030
rect 264973 121954 265039 121957
rect 440325 121954 440391 121957
rect 264973 121952 268180 121954
rect 264973 121896 264978 121952
rect 265034 121896 268180 121952
rect 264973 121894 268180 121896
rect 439852 121952 440391 121954
rect 439852 121896 440330 121952
rect 440386 121896 440391 121952
rect 439852 121894 440391 121896
rect 264973 121891 265039 121894
rect 440325 121891 440391 121894
rect 230933 121682 230999 121685
rect 228988 121680 230999 121682
rect 228988 121624 230938 121680
rect 230994 121624 230999 121680
rect 228988 121622 230999 121624
rect 230933 121619 230999 121622
rect 64689 121546 64755 121549
rect 66069 121546 66135 121549
rect 64689 121544 66135 121546
rect 64689 121488 64694 121544
rect 64750 121488 66074 121544
rect 66130 121488 66135 121544
rect 64689 121486 66135 121488
rect 64689 121483 64755 121486
rect 66069 121483 66135 121486
rect 266997 121546 267063 121549
rect 266997 121544 268180 121546
rect 266997 121488 267002 121544
rect 267058 121488 268180 121544
rect 266997 121486 268180 121488
rect 266997 121483 267063 121486
rect 214005 121410 214071 121413
rect 280429 121410 280495 121413
rect 214005 121408 217028 121410
rect 214005 121352 214010 121408
rect 214066 121352 217028 121408
rect 214005 121350 217028 121352
rect 279956 121408 280495 121410
rect 279956 121352 280434 121408
rect 280490 121352 280495 121408
rect 279956 121350 280495 121352
rect 214005 121347 214071 121350
rect 280429 121347 280495 121350
rect 231761 121274 231827 121277
rect 440182 121274 440188 121276
rect 228988 121272 231827 121274
rect 228988 121216 231766 121272
rect 231822 121216 231827 121272
rect 228988 121214 231827 121216
rect 439852 121214 440188 121274
rect 231761 121211 231827 121214
rect 440182 121212 440188 121214
rect 440252 121212 440258 121276
rect 397729 121138 397795 121141
rect 397729 121136 400108 121138
rect 66069 120866 66135 120869
rect 68142 120866 68816 120872
rect 268150 120866 268210 121108
rect 397729 121080 397734 121136
rect 397790 121080 400108 121136
rect 397729 121078 400108 121080
rect 397729 121075 397795 121078
rect 66069 120864 68816 120866
rect 66069 120808 66074 120864
rect 66130 120812 68816 120864
rect 66130 120808 68202 120812
rect 66069 120806 68202 120808
rect 258030 120806 268210 120866
rect 66069 120803 66135 120806
rect 213913 120730 213979 120733
rect 231669 120730 231735 120733
rect 213913 120728 217028 120730
rect 213913 120672 213918 120728
rect 213974 120672 217028 120728
rect 213913 120670 217028 120672
rect 228988 120728 231735 120730
rect 228988 120672 231674 120728
rect 231730 120672 231735 120728
rect 228988 120670 231735 120672
rect 213913 120667 213979 120670
rect 231669 120667 231735 120670
rect 232497 120458 232563 120461
rect 258030 120458 258090 120806
rect 439262 120804 439268 120868
rect 439332 120866 439338 120868
rect 439405 120866 439471 120869
rect 439332 120864 439471 120866
rect 439332 120808 439410 120864
rect 439466 120808 439471 120864
rect 439332 120806 439471 120808
rect 439332 120804 439338 120806
rect 439405 120803 439471 120806
rect 264973 120730 265039 120733
rect 282821 120730 282887 120733
rect 264973 120728 268180 120730
rect 264973 120672 264978 120728
rect 265034 120672 268180 120728
rect 264973 120670 268180 120672
rect 279956 120728 282887 120730
rect 279956 120672 282826 120728
rect 282882 120672 282887 120728
rect 279956 120670 282887 120672
rect 264973 120667 265039 120670
rect 282821 120667 282887 120670
rect 397637 120594 397703 120597
rect 397637 120592 400108 120594
rect 397637 120536 397642 120592
rect 397698 120536 400108 120592
rect 397637 120534 400108 120536
rect 397637 120531 397703 120534
rect 441613 120458 441679 120461
rect 232497 120456 258090 120458
rect 232497 120400 232502 120456
rect 232558 120400 258090 120456
rect 232497 120398 258090 120400
rect 439852 120456 441679 120458
rect 439852 120400 441618 120456
rect 441674 120400 441679 120456
rect 439852 120398 441679 120400
rect 232497 120395 232563 120398
rect 441613 120395 441679 120398
rect 230657 120322 230723 120325
rect 228988 120320 230723 120322
rect 228988 120264 230662 120320
rect 230718 120264 230723 120320
rect 228988 120262 230723 120264
rect 230657 120259 230723 120262
rect 265065 120322 265131 120325
rect 265065 120320 268180 120322
rect 265065 120264 265070 120320
rect 265126 120264 268180 120320
rect 265065 120262 268180 120264
rect 265065 120259 265131 120262
rect 231117 120186 231183 120189
rect 232865 120186 232931 120189
rect 231117 120184 232931 120186
rect 231117 120128 231122 120184
rect 231178 120128 232870 120184
rect 232926 120128 232931 120184
rect 231117 120126 232931 120128
rect 231117 120123 231183 120126
rect 232865 120123 232931 120126
rect 214005 120050 214071 120053
rect 361573 120050 361639 120053
rect 397729 120050 397795 120053
rect 214005 120048 217028 120050
rect 214005 119992 214010 120048
rect 214066 119992 217028 120048
rect 214005 119990 217028 119992
rect 361573 120048 397795 120050
rect 361573 119992 361578 120048
rect 361634 119992 397734 120048
rect 397790 119992 397795 120048
rect 361573 119990 397795 119992
rect 214005 119987 214071 119990
rect 361573 119987 361639 119990
rect 397729 119987 397795 119990
rect 282821 119914 282887 119917
rect 279956 119912 282887 119914
rect 279956 119856 282826 119912
rect 282882 119856 282887 119912
rect 279956 119854 282887 119856
rect 282821 119851 282887 119854
rect 397637 119914 397703 119917
rect 397637 119912 400108 119914
rect 397637 119856 397642 119912
rect 397698 119856 400108 119912
rect 397637 119854 400108 119856
rect 397637 119851 397703 119854
rect 234153 119778 234219 119781
rect 228988 119776 234219 119778
rect 228988 119720 234158 119776
rect 234214 119720 234219 119776
rect 228988 119718 234219 119720
rect 234153 119715 234219 119718
rect 213913 119506 213979 119509
rect 268150 119506 268210 119748
rect 213913 119504 217028 119506
rect 213913 119448 213918 119504
rect 213974 119448 217028 119504
rect 213913 119446 217028 119448
rect 258030 119446 268210 119506
rect 213913 119443 213979 119446
rect 231301 119370 231367 119373
rect 228988 119368 231367 119370
rect 228988 119312 231306 119368
rect 231362 119312 231367 119368
rect 228988 119310 231367 119312
rect 231301 119307 231367 119310
rect 233969 119098 234035 119101
rect 258030 119098 258090 119446
rect 264973 119370 265039 119373
rect 309777 119370 309843 119373
rect 361573 119370 361639 119373
rect 264973 119368 268180 119370
rect 264973 119312 264978 119368
rect 265034 119312 268180 119368
rect 264973 119310 268180 119312
rect 309777 119368 361639 119370
rect 309777 119312 309782 119368
rect 309838 119312 361578 119368
rect 361634 119312 361639 119368
rect 309777 119310 361639 119312
rect 439822 119370 439882 119748
rect 441654 119370 441660 119372
rect 439822 119310 441660 119370
rect 264973 119307 265039 119310
rect 309777 119307 309843 119310
rect 361573 119307 361639 119310
rect 441654 119308 441660 119310
rect 441724 119370 441730 119372
rect 447225 119370 447291 119373
rect 441724 119368 447291 119370
rect 441724 119312 447230 119368
rect 447286 119312 447291 119368
rect 441724 119310 447291 119312
rect 441724 119308 441730 119310
rect 447225 119307 447291 119310
rect 282729 119234 282795 119237
rect 279956 119232 282795 119234
rect 279956 119176 282734 119232
rect 282790 119176 282795 119232
rect 279956 119174 282795 119176
rect 282729 119171 282795 119174
rect 397545 119234 397611 119237
rect 397545 119232 400108 119234
rect 397545 119176 397550 119232
rect 397606 119176 400108 119232
rect 397545 119174 400108 119176
rect 397545 119171 397611 119174
rect 440417 119098 440483 119101
rect 233969 119096 258090 119098
rect 233969 119040 233974 119096
rect 234030 119040 258090 119096
rect 233969 119038 258090 119040
rect 439852 119096 440483 119098
rect 439852 119040 440422 119096
rect 440478 119040 440483 119096
rect 439852 119038 440483 119040
rect 233969 119035 234035 119038
rect 440417 119035 440483 119038
rect 231761 118962 231827 118965
rect 228988 118960 231827 118962
rect 228988 118904 231766 118960
rect 231822 118904 231827 118960
rect 228988 118902 231827 118904
rect 231761 118899 231827 118902
rect 265065 118962 265131 118965
rect 265065 118960 268180 118962
rect 265065 118904 265070 118960
rect 265126 118904 268180 118960
rect 265065 118902 268180 118904
rect 265065 118899 265131 118902
rect 184381 118826 184447 118829
rect 184381 118824 217028 118826
rect 184381 118768 184386 118824
rect 184442 118768 217028 118824
rect 184381 118766 217028 118768
rect 184381 118763 184447 118766
rect 264973 118554 265039 118557
rect 442901 118554 442967 118557
rect 264973 118552 268180 118554
rect 264973 118496 264978 118552
rect 265034 118496 268180 118552
rect 264973 118494 268180 118496
rect 439852 118552 442967 118554
rect 439852 118496 442906 118552
rect 442962 118496 442967 118552
rect 439852 118494 442967 118496
rect 264973 118491 265039 118494
rect 442901 118491 442967 118494
rect 231761 118418 231827 118421
rect 280153 118418 280219 118421
rect 228988 118416 231827 118418
rect 228988 118360 231766 118416
rect 231822 118360 231827 118416
rect 228988 118358 231827 118360
rect 279956 118416 280219 118418
rect 279956 118360 280158 118416
rect 280214 118360 280219 118416
rect 279956 118358 280219 118360
rect 231761 118355 231827 118358
rect 280153 118355 280219 118358
rect 397637 118418 397703 118421
rect 397637 118416 400108 118418
rect 397637 118360 397642 118416
rect 397698 118360 400108 118416
rect 397637 118358 400108 118360
rect 397637 118355 397703 118358
rect 214005 118146 214071 118149
rect 264329 118146 264395 118149
rect 214005 118144 217028 118146
rect 214005 118088 214010 118144
rect 214066 118088 217028 118144
rect 214005 118086 217028 118088
rect 264329 118144 268180 118146
rect 264329 118088 264334 118144
rect 264390 118088 268180 118144
rect 264329 118086 268180 118088
rect 214005 118083 214071 118086
rect 264329 118083 264395 118086
rect 230933 118010 230999 118013
rect 228988 118008 230999 118010
rect 228988 117952 230938 118008
rect 230994 117952 230999 118008
rect 228988 117950 230999 117952
rect 230933 117947 230999 117950
rect 231577 118010 231643 118013
rect 239581 118010 239647 118013
rect 231577 118008 239647 118010
rect 231577 117952 231582 118008
rect 231638 117952 239586 118008
rect 239642 117952 239647 118008
rect 231577 117950 239647 117952
rect 231577 117947 231643 117950
rect 239581 117947 239647 117950
rect 397545 117874 397611 117877
rect 397545 117872 400108 117874
rect 397545 117816 397550 117872
rect 397606 117816 400108 117872
rect 397545 117814 400108 117816
rect 397545 117811 397611 117814
rect 258030 117678 268180 117738
rect 243629 117602 243695 117605
rect 258030 117602 258090 117678
rect 282545 117602 282611 117605
rect 243629 117600 258090 117602
rect 243629 117544 243634 117600
rect 243690 117544 258090 117600
rect 243629 117542 258090 117544
rect 279956 117600 282611 117602
rect 279956 117544 282550 117600
rect 282606 117544 282611 117600
rect 279956 117542 282611 117544
rect 243629 117539 243695 117542
rect 282545 117539 282611 117542
rect 213913 117466 213979 117469
rect 231025 117466 231091 117469
rect 213913 117464 217028 117466
rect 213913 117408 213918 117464
rect 213974 117408 217028 117464
rect 213913 117406 217028 117408
rect 228988 117464 231091 117466
rect 228988 117408 231030 117464
rect 231086 117408 231091 117464
rect 228988 117406 231091 117408
rect 213913 117403 213979 117406
rect 231025 117403 231091 117406
rect 397545 117194 397611 117197
rect 442901 117194 442967 117197
rect 397545 117192 400108 117194
rect 229829 117058 229895 117061
rect 228988 117056 229895 117058
rect 228988 117000 229834 117056
rect 229890 117000 229895 117056
rect 228988 116998 229895 117000
rect 229829 116995 229895 116998
rect 262857 116922 262923 116925
rect 268150 116922 268210 117164
rect 397545 117136 397550 117192
rect 397606 117136 400108 117192
rect 397545 117134 400108 117136
rect 439852 117192 442967 117194
rect 439852 117136 442906 117192
rect 442962 117136 442967 117192
rect 439852 117134 442967 117136
rect 397545 117131 397611 117134
rect 442901 117131 442967 117134
rect 282269 116922 282335 116925
rect 262857 116920 268210 116922
rect 262857 116864 262862 116920
rect 262918 116864 268210 116920
rect 262857 116862 268210 116864
rect 279956 116920 282335 116922
rect 279956 116864 282274 116920
rect 282330 116864 282335 116920
rect 279956 116862 282335 116864
rect 262857 116859 262923 116862
rect 282269 116859 282335 116862
rect 214005 116786 214071 116789
rect 265157 116786 265223 116789
rect 214005 116784 217028 116786
rect 214005 116728 214010 116784
rect 214066 116728 217028 116784
rect 214005 116726 217028 116728
rect 265157 116784 268180 116786
rect 265157 116728 265162 116784
rect 265218 116728 268180 116784
rect 265157 116726 268180 116728
rect 214005 116723 214071 116726
rect 265157 116723 265223 116726
rect 231485 116514 231551 116517
rect 228988 116512 231551 116514
rect 228988 116456 231490 116512
rect 231546 116456 231551 116512
rect 228988 116454 231551 116456
rect 231485 116451 231551 116454
rect 442901 116378 442967 116381
rect 258030 116318 268180 116378
rect 439852 116376 442967 116378
rect 439852 116320 442906 116376
rect 442962 116320 442967 116376
rect 439852 116318 442967 116320
rect 230974 116180 230980 116244
rect 231044 116242 231050 116244
rect 258030 116242 258090 116318
rect 442901 116315 442967 116318
rect 231044 116182 258090 116242
rect 231044 116180 231050 116182
rect 213913 116106 213979 116109
rect 230749 116106 230815 116109
rect 213913 116104 217028 116106
rect 213913 116048 213918 116104
rect 213974 116048 217028 116104
rect 213913 116046 217028 116048
rect 228988 116104 230815 116106
rect 228988 116048 230754 116104
rect 230810 116048 230815 116104
rect 228988 116046 230815 116048
rect 213913 116043 213979 116046
rect 230749 116043 230815 116046
rect 246246 116044 246252 116108
rect 246316 116106 246322 116108
rect 262857 116106 262923 116109
rect 282821 116106 282887 116109
rect 246316 116104 262923 116106
rect 246316 116048 262862 116104
rect 262918 116048 262923 116104
rect 246316 116046 262923 116048
rect 279956 116104 282887 116106
rect 279956 116048 282826 116104
rect 282882 116048 282887 116104
rect 279956 116046 282887 116048
rect 246316 116044 246322 116046
rect 262857 116043 262923 116046
rect 282821 116043 282887 116046
rect 264973 115970 265039 115973
rect 264973 115968 268180 115970
rect 264973 115912 264978 115968
rect 265034 115912 268180 115968
rect 264973 115910 268180 115912
rect 264973 115907 265039 115910
rect 439262 115908 439268 115972
rect 439332 115970 439338 115972
rect 439405 115970 439471 115973
rect 439332 115968 439471 115970
rect 439332 115912 439410 115968
rect 439466 115912 439471 115968
rect 439332 115910 439471 115912
rect 439332 115908 439338 115910
rect 439405 115907 439471 115910
rect 397545 115834 397611 115837
rect 442901 115834 442967 115837
rect 397545 115832 400108 115834
rect 397545 115776 397550 115832
rect 397606 115776 400108 115832
rect 397545 115774 400108 115776
rect 439852 115832 442967 115834
rect 439852 115776 442906 115832
rect 442962 115776 442967 115832
rect 439852 115774 442967 115776
rect 397545 115771 397611 115774
rect 442901 115771 442967 115774
rect 246297 115562 246363 115565
rect 228988 115560 246363 115562
rect 228988 115504 246302 115560
rect 246358 115504 246363 115560
rect 228988 115502 246363 115504
rect 246297 115499 246363 115502
rect 214005 115426 214071 115429
rect 214005 115424 217028 115426
rect 214005 115368 214010 115424
rect 214066 115368 217028 115424
rect 214005 115366 217028 115368
rect 214005 115363 214071 115366
rect 268150 115290 268210 115532
rect 282177 115426 282243 115429
rect 279956 115424 282243 115426
rect 279956 115368 282182 115424
rect 282238 115368 282243 115424
rect 279956 115366 282243 115368
rect 282177 115363 282243 115366
rect 258030 115230 268210 115290
rect 197261 115154 197327 115157
rect 209221 115154 209287 115157
rect 231485 115154 231551 115157
rect 197261 115152 209287 115154
rect 197261 115096 197266 115152
rect 197322 115096 209226 115152
rect 209282 115096 209287 115152
rect 197261 115094 209287 115096
rect 228988 115152 231551 115154
rect 228988 115096 231490 115152
rect 231546 115096 231551 115152
rect 228988 115094 231551 115096
rect 197261 115091 197327 115094
rect 209221 115091 209287 115094
rect 231485 115091 231551 115094
rect 213913 114882 213979 114885
rect 229829 114882 229895 114885
rect 258030 114882 258090 115230
rect 265065 115154 265131 115157
rect 397637 115154 397703 115157
rect 265065 115152 268180 115154
rect 265065 115096 265070 115152
rect 265126 115096 268180 115152
rect 265065 115094 268180 115096
rect 397637 115152 400108 115154
rect 397637 115096 397642 115152
rect 397698 115096 400108 115152
rect 397637 115094 400108 115096
rect 265065 115091 265131 115094
rect 397637 115091 397703 115094
rect 440325 115018 440391 115021
rect 439852 115016 440391 115018
rect 439852 114960 440330 115016
rect 440386 114960 440391 115016
rect 439852 114958 440391 114960
rect 440325 114955 440391 114958
rect 213913 114880 217028 114882
rect 213913 114824 213918 114880
rect 213974 114824 217028 114880
rect 213913 114822 217028 114824
rect 229829 114880 258090 114882
rect 229829 114824 229834 114880
rect 229890 114824 258090 114880
rect 229829 114822 258090 114824
rect 213913 114819 213979 114822
rect 229829 114819 229895 114822
rect 230657 114610 230723 114613
rect 228988 114608 230723 114610
rect 228988 114552 230662 114608
rect 230718 114552 230723 114608
rect 228988 114550 230723 114552
rect 230657 114547 230723 114550
rect 264973 114610 265039 114613
rect 282453 114610 282519 114613
rect 264973 114608 268180 114610
rect 264973 114552 264978 114608
rect 265034 114552 268180 114608
rect 264973 114550 268180 114552
rect 279956 114608 282519 114610
rect 279956 114552 282458 114608
rect 282514 114552 282519 114608
rect 279956 114550 282519 114552
rect 264973 114547 265039 114550
rect 282453 114547 282519 114550
rect 397545 114474 397611 114477
rect 440877 114474 440943 114477
rect 397545 114472 400108 114474
rect 397545 114416 397550 114472
rect 397606 114416 400108 114472
rect 397545 114414 400108 114416
rect 439852 114472 440943 114474
rect 439852 114416 440882 114472
rect 440938 114416 440943 114472
rect 439852 114414 440943 114416
rect 397545 114411 397611 114414
rect 440877 114411 440943 114414
rect 213913 114202 213979 114205
rect 231761 114202 231827 114205
rect 213913 114200 217028 114202
rect 213913 114144 213918 114200
rect 213974 114144 217028 114200
rect 213913 114142 217028 114144
rect 228988 114200 231827 114202
rect 228988 114144 231766 114200
rect 231822 114144 231827 114200
rect 228988 114142 231827 114144
rect 213913 114139 213979 114142
rect 231761 114139 231827 114142
rect 264973 114202 265039 114205
rect 264973 114200 268180 114202
rect 264973 114144 264978 114200
rect 265034 114144 268180 114200
rect 264973 114142 268180 114144
rect 264973 114139 265039 114142
rect 242433 113930 242499 113933
rect 265157 113930 265223 113933
rect 242433 113928 265223 113930
rect 242433 113872 242438 113928
rect 242494 113872 265162 113928
rect 265218 113872 265223 113928
rect 242433 113870 265223 113872
rect 242433 113867 242499 113870
rect 265157 113867 265223 113870
rect 231393 113794 231459 113797
rect 264605 113794 264671 113797
rect 231393 113792 264671 113794
rect 231393 113736 231398 113792
rect 231454 113736 264610 113792
rect 264666 113736 264671 113792
rect 231393 113734 264671 113736
rect 231393 113731 231459 113734
rect 264605 113731 264671 113734
rect 267774 113732 267780 113796
rect 267844 113794 267850 113796
rect 282821 113794 282887 113797
rect 267844 113734 268180 113794
rect 279956 113792 282887 113794
rect 279956 113736 282826 113792
rect 282882 113736 282887 113792
rect 279956 113734 282887 113736
rect 267844 113732 267850 113734
rect 282821 113731 282887 113734
rect 397637 113794 397703 113797
rect 397637 113792 400108 113794
rect 397637 113736 397642 113792
rect 397698 113736 400108 113792
rect 397637 113734 400108 113736
rect 397637 113731 397703 113734
rect 231669 113658 231735 113661
rect 442901 113658 442967 113661
rect 228988 113656 231735 113658
rect 228988 113600 231674 113656
rect 231730 113600 231735 113656
rect 228988 113598 231735 113600
rect 439852 113656 442967 113658
rect 439852 113600 442906 113656
rect 442962 113600 442967 113656
rect 439852 113598 442967 113600
rect 231669 113595 231735 113598
rect 442901 113595 442967 113598
rect 199377 113386 199443 113389
rect 216998 113386 217058 113492
rect 199377 113384 217058 113386
rect 199377 113328 199382 113384
rect 199438 113328 217058 113384
rect 199377 113326 217058 113328
rect 199377 113323 199443 113326
rect 266854 113324 266860 113388
rect 266924 113386 266930 113388
rect 266924 113326 268180 113386
rect 266924 113324 266930 113326
rect 229921 113250 229987 113253
rect 228988 113248 229987 113250
rect 228988 113192 229926 113248
rect 229982 113192 229987 113248
rect 228988 113190 229987 113192
rect 229921 113187 229987 113190
rect 281809 113114 281875 113117
rect 442901 113114 442967 113117
rect 279956 113112 281875 113114
rect 279956 113056 281814 113112
rect 281870 113056 281875 113112
rect 279956 113054 281875 113056
rect 439852 113112 442967 113114
rect 439852 113056 442906 113112
rect 442962 113056 442967 113112
rect 439852 113054 442967 113056
rect 281809 113051 281875 113054
rect 442901 113051 442967 113054
rect 398741 112978 398807 112981
rect 398741 112976 400108 112978
rect 214005 112842 214071 112845
rect 214005 112840 217028 112842
rect 214005 112784 214010 112840
rect 214066 112784 217028 112840
rect 214005 112782 217028 112784
rect 214005 112779 214071 112782
rect 230933 112706 230999 112709
rect 268150 112706 268210 112948
rect 398741 112920 398746 112976
rect 398802 112920 400108 112976
rect 398741 112918 400108 112920
rect 398741 112915 398807 112918
rect 583017 112842 583083 112845
rect 583520 112842 584960 112932
rect 583017 112840 584960 112842
rect 583017 112784 583022 112840
rect 583078 112784 584960 112840
rect 583017 112782 584960 112784
rect 583017 112779 583083 112782
rect 228988 112704 230999 112706
rect 228988 112648 230938 112704
rect 230994 112648 230999 112704
rect 228988 112646 230999 112648
rect 230933 112643 230999 112646
rect 258030 112646 268210 112706
rect 583520 112692 584960 112782
rect 170254 112372 170260 112436
rect 170324 112434 170330 112436
rect 202137 112434 202203 112437
rect 170324 112432 202203 112434
rect 170324 112376 202142 112432
rect 202198 112376 202203 112432
rect 170324 112374 202203 112376
rect 170324 112372 170330 112374
rect 202137 112371 202203 112374
rect 231761 112298 231827 112301
rect 228988 112296 231827 112298
rect 228988 112240 231766 112296
rect 231822 112240 231827 112296
rect 228988 112238 231827 112240
rect 231761 112235 231827 112238
rect 213913 112162 213979 112165
rect 232681 112162 232747 112165
rect 258030 112162 258090 112646
rect 264973 112570 265039 112573
rect 264973 112568 268180 112570
rect 264973 112512 264978 112568
rect 265034 112512 268180 112568
rect 264973 112510 268180 112512
rect 264973 112507 265039 112510
rect 397545 112434 397611 112437
rect 397545 112432 400108 112434
rect 397545 112376 397550 112432
rect 397606 112376 400108 112432
rect 397545 112374 400108 112376
rect 397545 112371 397611 112374
rect 282821 112298 282887 112301
rect 279956 112296 282887 112298
rect 279956 112240 282826 112296
rect 282882 112240 282887 112296
rect 279956 112238 282887 112240
rect 282821 112235 282887 112238
rect 213913 112160 217028 112162
rect 213913 112104 213918 112160
rect 213974 112104 217028 112160
rect 213913 112102 217028 112104
rect 232681 112160 258090 112162
rect 232681 112104 232686 112160
rect 232742 112104 258090 112160
rect 232681 112102 258090 112104
rect 213913 112099 213979 112102
rect 232681 112099 232747 112102
rect 264237 112026 264303 112029
rect 264237 112024 268180 112026
rect 264237 111968 264242 112024
rect 264298 111968 268180 112024
rect 264237 111966 268180 111968
rect 264237 111963 264303 111966
rect 439313 111890 439379 111893
rect 439270 111888 439379 111890
rect 439270 111832 439318 111888
rect 439374 111832 439379 111888
rect 439270 111827 439379 111832
rect 164724 111754 165354 111760
rect 167637 111754 167703 111757
rect 231577 111754 231643 111757
rect 164724 111752 167703 111754
rect 164724 111700 167642 111752
rect 165294 111696 167642 111700
rect 167698 111696 167703 111752
rect 165294 111694 167703 111696
rect 228988 111752 231643 111754
rect 228988 111696 231582 111752
rect 231638 111696 231643 111752
rect 228988 111694 231643 111696
rect 167637 111691 167703 111694
rect 231577 111691 231643 111694
rect 397453 111754 397519 111757
rect 397453 111752 400108 111754
rect 397453 111696 397458 111752
rect 397514 111696 400108 111752
rect 439270 111724 439330 111827
rect 397453 111694 400108 111696
rect 397453 111691 397519 111694
rect 265065 111618 265131 111621
rect 282821 111618 282887 111621
rect 265065 111616 268180 111618
rect 265065 111560 265070 111616
rect 265126 111560 268180 111616
rect 265065 111558 268180 111560
rect 279956 111616 282887 111618
rect 279956 111560 282826 111616
rect 282882 111560 282887 111616
rect 279956 111558 282887 111560
rect 265065 111555 265131 111558
rect 282821 111555 282887 111558
rect 214005 111482 214071 111485
rect 214005 111480 217028 111482
rect 214005 111424 214010 111480
rect 214066 111424 217028 111480
rect 214005 111422 217028 111424
rect 214005 111419 214071 111422
rect 231761 111346 231827 111349
rect 228988 111344 231827 111346
rect 228988 111288 231766 111344
rect 231822 111288 231827 111344
rect 228988 111286 231827 111288
rect 231761 111283 231827 111286
rect 439262 111284 439268 111348
rect 439332 111284 439338 111348
rect 264973 111210 265039 111213
rect 264973 111208 268180 111210
rect 264973 111152 264978 111208
rect 265034 111152 268180 111208
rect 264973 111150 268180 111152
rect 264973 111147 265039 111150
rect 231485 111074 231551 111077
rect 242249 111074 242315 111077
rect 231485 111072 242315 111074
rect 231485 111016 231490 111072
rect 231546 111016 242254 111072
rect 242310 111016 242315 111072
rect 231485 111014 242315 111016
rect 231485 111011 231551 111014
rect 242249 111011 242315 111014
rect 302734 111012 302740 111076
rect 302804 111074 302810 111076
rect 398189 111074 398255 111077
rect 302804 111072 398255 111074
rect 302804 111016 398194 111072
rect 398250 111016 398255 111072
rect 439270 111044 439330 111284
rect 302804 111014 398255 111016
rect 302804 111012 302810 111014
rect 398189 111011 398255 111014
rect 213913 110802 213979 110805
rect 230749 110802 230815 110805
rect 213913 110800 217028 110802
rect -960 110666 480 110756
rect 213913 110744 213918 110800
rect 213974 110744 217028 110800
rect 213913 110742 217028 110744
rect 228988 110800 230815 110802
rect 228988 110744 230754 110800
rect 230810 110744 230815 110800
rect 228988 110742 230815 110744
rect 213913 110739 213979 110742
rect 230749 110739 230815 110742
rect 238293 110802 238359 110805
rect 281533 110802 281599 110805
rect 238293 110800 268180 110802
rect 238293 110744 238298 110800
rect 238354 110744 268180 110800
rect 238293 110742 268180 110744
rect 279956 110800 281599 110802
rect 279956 110744 281538 110800
rect 281594 110744 281599 110800
rect 279956 110742 281599 110744
rect 238293 110739 238359 110742
rect 281533 110739 281599 110742
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 193949 110530 194015 110533
rect 198181 110530 198247 110533
rect 193949 110528 198247 110530
rect 193949 110472 193954 110528
rect 194010 110472 198186 110528
rect 198242 110472 198247 110528
rect 193949 110470 198247 110472
rect 193949 110467 194015 110470
rect 198181 110467 198247 110470
rect 247953 110394 248019 110397
rect 228988 110392 248019 110394
rect 228988 110336 247958 110392
rect 248014 110336 248019 110392
rect 228988 110334 248019 110336
rect 247953 110331 248019 110334
rect 265065 110394 265131 110397
rect 265065 110392 268180 110394
rect 265065 110336 265070 110392
rect 265126 110336 268180 110392
rect 265065 110334 268180 110336
rect 265065 110331 265131 110334
rect 214005 110258 214071 110261
rect 397545 110258 397611 110261
rect 214005 110256 217028 110258
rect 214005 110200 214010 110256
rect 214066 110200 217028 110256
rect 214005 110198 217028 110200
rect 397545 110256 400108 110258
rect 397545 110200 397550 110256
rect 397606 110200 400108 110256
rect 397545 110198 400108 110200
rect 214005 110195 214071 110198
rect 397545 110195 397611 110198
rect 164724 110122 165354 110128
rect 167729 110122 167795 110125
rect 164724 110120 167795 110122
rect 164724 110068 167734 110120
rect 165294 110064 167734 110068
rect 167790 110064 167795 110120
rect 165294 110062 167795 110064
rect 167729 110059 167795 110062
rect 283782 109986 283788 109988
rect 231669 109850 231735 109853
rect 228988 109848 231735 109850
rect 228988 109792 231674 109848
rect 231730 109792 231735 109848
rect 228988 109790 231735 109792
rect 231669 109787 231735 109790
rect 258073 109714 258139 109717
rect 268150 109714 268210 109956
rect 279956 109926 283788 109986
rect 283782 109924 283788 109926
rect 283852 109924 283858 109988
rect 439822 109850 439882 110228
rect 446029 109850 446095 109853
rect 449985 109850 450051 109853
rect 439822 109848 450051 109850
rect 439822 109792 446034 109848
rect 446090 109792 449990 109848
rect 450046 109792 450051 109848
rect 439822 109790 450051 109792
rect 446029 109787 446095 109790
rect 449985 109787 450051 109790
rect 258073 109712 268210 109714
rect 258073 109656 258078 109712
rect 258134 109656 268210 109712
rect 258073 109654 268210 109656
rect 258073 109651 258139 109654
rect 213913 109578 213979 109581
rect 442165 109578 442231 109581
rect 213913 109576 217028 109578
rect 213913 109520 213918 109576
rect 213974 109520 217028 109576
rect 213913 109518 217028 109520
rect 258030 109518 268180 109578
rect 439852 109576 442231 109578
rect 213913 109515 213979 109518
rect 231761 109442 231827 109445
rect 228988 109440 231827 109442
rect 228988 109384 231766 109440
rect 231822 109384 231827 109440
rect 228988 109382 231827 109384
rect 231761 109379 231827 109382
rect 241053 109442 241119 109445
rect 258030 109442 258090 109518
rect 241053 109440 258090 109442
rect 241053 109384 241058 109440
rect 241114 109384 258090 109440
rect 241053 109382 258090 109384
rect 241053 109379 241119 109382
rect 250621 109306 250687 109309
rect 258073 109306 258139 109309
rect 282821 109306 282887 109309
rect 400078 109306 400138 109548
rect 439852 109520 442170 109576
rect 442226 109520 442231 109576
rect 439852 109518 442231 109520
rect 442165 109515 442231 109518
rect 250621 109304 258139 109306
rect 250621 109248 250626 109304
rect 250682 109248 258078 109304
rect 258134 109248 258139 109304
rect 250621 109246 258139 109248
rect 279956 109304 282887 109306
rect 279956 109248 282826 109304
rect 282882 109248 282887 109304
rect 279956 109246 282887 109248
rect 250621 109243 250687 109246
rect 258073 109243 258139 109246
rect 282821 109243 282887 109246
rect 287010 109246 400138 109306
rect 282126 109108 282132 109172
rect 282196 109170 282202 109172
rect 287010 109170 287070 109246
rect 282196 109110 287070 109170
rect 282196 109108 282202 109110
rect 253381 109034 253447 109037
rect 238710 109032 253447 109034
rect 238710 108976 253386 109032
rect 253442 108976 253447 109032
rect 238710 108974 253447 108976
rect 214005 108898 214071 108901
rect 238710 108898 238770 108974
rect 253381 108971 253447 108974
rect 264973 109034 265039 109037
rect 397453 109034 397519 109037
rect 442441 109034 442507 109037
rect 264973 109032 268180 109034
rect 264973 108976 264978 109032
rect 265034 108976 268180 109032
rect 264973 108974 268180 108976
rect 397453 109032 400108 109034
rect 397453 108976 397458 109032
rect 397514 108976 400108 109032
rect 397453 108974 400108 108976
rect 439852 109032 442507 109034
rect 439852 108976 442446 109032
rect 442502 108976 442507 109032
rect 439852 108974 442507 108976
rect 264973 108971 265039 108974
rect 397453 108971 397519 108974
rect 442441 108971 442507 108974
rect 214005 108896 217028 108898
rect 214005 108840 214010 108896
rect 214066 108840 217028 108896
rect 214005 108838 217028 108840
rect 228988 108838 238770 108898
rect 214005 108835 214071 108838
rect 164724 108762 165354 108768
rect 167545 108762 167611 108765
rect 164724 108760 167611 108762
rect 164724 108708 167550 108760
rect 165294 108704 167550 108708
rect 167606 108704 167611 108760
rect 165294 108702 167611 108704
rect 167545 108699 167611 108702
rect 264421 108626 264487 108629
rect 264421 108624 268180 108626
rect 264421 108568 264426 108624
rect 264482 108568 268180 108624
rect 264421 108566 268180 108568
rect 264421 108563 264487 108566
rect 231761 108490 231827 108493
rect 282269 108490 282335 108493
rect 228988 108488 231827 108490
rect 228988 108432 231766 108488
rect 231822 108432 231827 108488
rect 228988 108430 231827 108432
rect 279956 108488 282335 108490
rect 279956 108432 282274 108488
rect 282330 108432 282335 108488
rect 279956 108430 282335 108432
rect 231761 108427 231827 108430
rect 282269 108427 282335 108430
rect 324957 108354 325023 108357
rect 397494 108354 397500 108356
rect 324957 108352 397500 108354
rect 324957 108296 324962 108352
rect 325018 108296 397500 108352
rect 324957 108294 397500 108296
rect 324957 108291 325023 108294
rect 397494 108292 397500 108294
rect 397564 108292 397570 108356
rect 397637 108354 397703 108357
rect 397637 108352 400108 108354
rect 397637 108296 397642 108352
rect 397698 108296 400108 108352
rect 397637 108294 400108 108296
rect 397637 108291 397703 108294
rect 213913 108218 213979 108221
rect 441705 108218 441771 108221
rect 213913 108216 217028 108218
rect 213913 108160 213918 108216
rect 213974 108160 217028 108216
rect 213913 108158 217028 108160
rect 258030 108158 268180 108218
rect 439852 108216 441771 108218
rect 439852 108160 441710 108216
rect 441766 108160 441771 108216
rect 439852 108158 441771 108160
rect 213913 108155 213979 108158
rect 247953 108082 248019 108085
rect 258030 108082 258090 108158
rect 441705 108155 441771 108158
rect 247953 108080 258090 108082
rect 247953 108024 247958 108080
rect 248014 108024 258090 108080
rect 247953 108022 258090 108024
rect 247953 108019 248019 108022
rect 231301 107946 231367 107949
rect 228988 107944 231367 107946
rect 228988 107888 231306 107944
rect 231362 107888 231367 107944
rect 228988 107886 231367 107888
rect 231301 107883 231367 107886
rect 282361 107810 282427 107813
rect 258030 107750 268180 107810
rect 279956 107808 282427 107810
rect 279956 107752 282366 107808
rect 282422 107752 282427 107808
rect 279956 107750 282427 107752
rect 242249 107674 242315 107677
rect 258030 107674 258090 107750
rect 282361 107747 282427 107750
rect 242249 107672 258090 107674
rect 242249 107616 242254 107672
rect 242310 107616 258090 107672
rect 242249 107614 258090 107616
rect 242249 107611 242315 107614
rect 214005 107538 214071 107541
rect 264094 107538 264100 107540
rect 214005 107536 217028 107538
rect 214005 107480 214010 107536
rect 214066 107480 217028 107536
rect 214005 107478 217028 107480
rect 228988 107478 264100 107538
rect 214005 107475 214071 107478
rect 264094 107476 264100 107478
rect 264164 107476 264170 107540
rect 397453 107538 397519 107541
rect 442901 107538 442967 107541
rect 397453 107536 400108 107538
rect 397453 107480 397458 107536
rect 397514 107480 400108 107536
rect 397453 107478 400108 107480
rect 439852 107536 442967 107538
rect 439852 107480 442906 107536
rect 442962 107480 442967 107536
rect 439852 107478 442967 107480
rect 397453 107475 397519 107478
rect 442901 107475 442967 107478
rect 231761 107130 231827 107133
rect 228988 107128 231827 107130
rect 228988 107072 231766 107128
rect 231822 107072 231827 107128
rect 228988 107070 231827 107072
rect 231761 107067 231827 107070
rect 258901 107130 258967 107133
rect 268150 107130 268210 107372
rect 258901 107128 268210 107130
rect 258901 107072 258906 107128
rect 258962 107072 268210 107128
rect 258901 107070 268210 107072
rect 258901 107067 258967 107070
rect 265249 106994 265315 106997
rect 282821 106994 282887 106997
rect 265249 106992 268180 106994
rect 265249 106936 265254 106992
rect 265310 106936 268180 106992
rect 265249 106934 268180 106936
rect 279956 106992 282887 106994
rect 279956 106936 282826 106992
rect 282882 106936 282887 106992
rect 279956 106934 282887 106936
rect 265249 106931 265315 106934
rect 282821 106931 282887 106934
rect 213913 106858 213979 106861
rect 397545 106858 397611 106861
rect 213913 106856 217028 106858
rect 213913 106800 213918 106856
rect 213974 106800 217028 106856
rect 213913 106798 217028 106800
rect 397545 106856 400108 106858
rect 397545 106800 397550 106856
rect 397606 106800 400108 106856
rect 397545 106798 400108 106800
rect 213913 106795 213979 106798
rect 397545 106795 397611 106798
rect 231669 106586 231735 106589
rect 228988 106584 231735 106586
rect 228988 106528 231674 106584
rect 231730 106528 231735 106584
rect 228988 106526 231735 106528
rect 231669 106523 231735 106526
rect 267273 106450 267339 106453
rect 267273 106448 268180 106450
rect 267273 106392 267278 106448
rect 267334 106392 268180 106448
rect 267273 106390 268180 106392
rect 267273 106387 267339 106390
rect 214005 106178 214071 106181
rect 231577 106178 231643 106181
rect 214005 106176 217028 106178
rect 214005 106120 214010 106176
rect 214066 106120 217028 106176
rect 214005 106118 217028 106120
rect 228988 106176 231643 106178
rect 228988 106120 231582 106176
rect 231638 106120 231643 106176
rect 397453 106178 397519 106181
rect 442349 106178 442415 106181
rect 397453 106176 400108 106178
rect 228988 106118 231643 106120
rect 214005 106115 214071 106118
rect 231577 106115 231643 106118
rect 264973 106042 265039 106045
rect 264973 106040 268180 106042
rect 264973 105984 264978 106040
rect 265034 105984 268180 106040
rect 264973 105982 268180 105984
rect 264973 105979 265039 105982
rect 279374 105773 279434 106148
rect 397453 106120 397458 106176
rect 397514 106120 400108 106176
rect 397453 106118 400108 106120
rect 439852 106176 442415 106178
rect 439852 106120 442354 106176
rect 442410 106120 442415 106176
rect 439852 106118 442415 106120
rect 397453 106115 397519 106118
rect 442349 106115 442415 106118
rect 279325 105768 279434 105773
rect 279325 105712 279330 105768
rect 279386 105712 279434 105768
rect 279325 105710 279434 105712
rect 279325 105707 279391 105710
rect 213913 105634 213979 105637
rect 231301 105634 231367 105637
rect 213913 105632 217028 105634
rect 213913 105576 213918 105632
rect 213974 105576 217028 105632
rect 213913 105574 217028 105576
rect 228988 105632 231367 105634
rect 228988 105576 231306 105632
rect 231362 105576 231367 105632
rect 228988 105574 231367 105576
rect 213913 105571 213979 105574
rect 231301 105571 231367 105574
rect 265157 105634 265223 105637
rect 442717 105634 442783 105637
rect 265157 105632 268180 105634
rect 265157 105576 265162 105632
rect 265218 105576 268180 105632
rect 265157 105574 268180 105576
rect 439852 105632 442783 105634
rect 439852 105576 442722 105632
rect 442778 105576 442783 105632
rect 439852 105574 442783 105576
rect 265157 105571 265223 105574
rect 442717 105571 442783 105574
rect 280245 105498 280311 105501
rect 279956 105496 280311 105498
rect 279956 105440 280250 105496
rect 280306 105440 280311 105496
rect 279956 105438 280311 105440
rect 280245 105435 280311 105438
rect 231209 105226 231275 105229
rect 228988 105224 231275 105226
rect 228988 105168 231214 105224
rect 231270 105168 231275 105224
rect 228988 105166 231275 105168
rect 231209 105163 231275 105166
rect 233877 105226 233943 105229
rect 233877 105224 268180 105226
rect 233877 105168 233882 105224
rect 233938 105168 268180 105224
rect 233877 105166 268180 105168
rect 233877 105163 233943 105166
rect 214741 104954 214807 104957
rect 279417 104954 279483 104957
rect 214741 104952 217028 104954
rect 214741 104896 214746 104952
rect 214802 104896 217028 104952
rect 214741 104894 217028 104896
rect 279374 104952 279483 104954
rect 279374 104896 279422 104952
rect 279478 104896 279483 104952
rect 214741 104891 214807 104894
rect 279374 104891 279483 104896
rect 265065 104818 265131 104821
rect 265065 104816 268180 104818
rect 265065 104760 265070 104816
rect 265126 104760 268180 104816
rect 265065 104758 268180 104760
rect 265065 104755 265131 104758
rect 231669 104682 231735 104685
rect 228988 104680 231735 104682
rect 228988 104624 231674 104680
rect 231730 104624 231735 104680
rect 279374 104652 279434 104891
rect 397453 104818 397519 104821
rect 397453 104816 400108 104818
rect 397453 104760 397458 104816
rect 397514 104760 400108 104816
rect 397453 104758 400108 104760
rect 397453 104755 397519 104758
rect 228988 104622 231735 104624
rect 231669 104619 231735 104622
rect 439270 104413 439330 104788
rect 264973 104410 265039 104413
rect 264973 104408 268180 104410
rect 264973 104352 264978 104408
rect 265034 104352 268180 104408
rect 264973 104350 268180 104352
rect 439270 104408 439379 104413
rect 439270 104352 439318 104408
rect 439374 104352 439379 104408
rect 439270 104350 439379 104352
rect 264973 104347 265039 104350
rect 439313 104347 439379 104350
rect 232446 104274 232452 104276
rect 181529 103866 181595 103869
rect 216998 103866 217058 104244
rect 228988 104214 232452 104274
rect 232446 104212 232452 104214
rect 232516 104212 232522 104276
rect 397545 104274 397611 104277
rect 397545 104272 400108 104274
rect 397545 104216 397550 104272
rect 397606 104216 400108 104272
rect 397545 104214 400108 104216
rect 397545 104211 397611 104214
rect 380157 104138 380223 104141
rect 398649 104138 398715 104141
rect 380157 104136 398715 104138
rect 380157 104080 380162 104136
rect 380218 104080 398654 104136
rect 398710 104080 398715 104136
rect 380157 104078 398715 104080
rect 380157 104075 380223 104078
rect 398649 104075 398715 104078
rect 281533 104002 281599 104005
rect 279956 104000 281599 104002
rect 279956 103944 281538 104000
rect 281594 103944 281599 104000
rect 279956 103942 281599 103944
rect 281533 103939 281599 103942
rect 439454 103869 439514 104108
rect 181529 103864 217058 103866
rect 181529 103808 181534 103864
rect 181590 103808 217058 103864
rect 181529 103806 217058 103808
rect 264513 103866 264579 103869
rect 264513 103864 268180 103866
rect 264513 103808 264518 103864
rect 264574 103808 268180 103864
rect 264513 103806 268180 103808
rect 439405 103864 439514 103869
rect 439405 103808 439410 103864
rect 439466 103808 439514 103864
rect 439405 103806 439514 103808
rect 181529 103803 181595 103806
rect 264513 103803 264579 103806
rect 439405 103803 439471 103806
rect 231761 103730 231827 103733
rect 228988 103728 231827 103730
rect 228988 103672 231766 103728
rect 231822 103672 231827 103728
rect 228988 103670 231827 103672
rect 231761 103667 231827 103670
rect 213269 103594 213335 103597
rect 213269 103592 217028 103594
rect 213269 103536 213274 103592
rect 213330 103536 217028 103592
rect 213269 103534 217028 103536
rect 213269 103531 213335 103534
rect 264973 103458 265039 103461
rect 397453 103458 397519 103461
rect 443177 103458 443243 103461
rect 264973 103456 268180 103458
rect 264973 103400 264978 103456
rect 265034 103400 268180 103456
rect 264973 103398 268180 103400
rect 397453 103456 400108 103458
rect 397453 103400 397458 103456
rect 397514 103400 400108 103456
rect 397453 103398 400108 103400
rect 439852 103456 443243 103458
rect 439852 103400 443182 103456
rect 443238 103400 443243 103456
rect 439852 103398 443243 103400
rect 264973 103395 265039 103398
rect 397453 103395 397519 103398
rect 443177 103395 443243 103398
rect 231117 103322 231183 103325
rect 228988 103320 231183 103322
rect 228988 103264 231122 103320
rect 231178 103264 231183 103320
rect 228988 103262 231183 103264
rect 231117 103259 231183 103262
rect 281625 103186 281691 103189
rect 279956 103184 281691 103186
rect 279956 103128 281630 103184
rect 281686 103128 281691 103184
rect 279956 103126 281691 103128
rect 281625 103123 281691 103126
rect 370497 103186 370563 103189
rect 399886 103186 399892 103188
rect 370497 103184 399892 103186
rect 370497 103128 370502 103184
rect 370558 103128 399892 103184
rect 370497 103126 399892 103128
rect 370497 103123 370563 103126
rect 399886 103124 399892 103126
rect 399956 103124 399962 103188
rect 258030 102990 268180 103050
rect 239581 102914 239647 102917
rect 258030 102914 258090 102990
rect 239581 102912 258090 102914
rect 170254 102444 170260 102508
rect 170324 102506 170330 102508
rect 216998 102506 217058 102884
rect 239581 102856 239586 102912
rect 239642 102856 258090 102912
rect 239581 102854 258090 102856
rect 239581 102851 239647 102854
rect 231301 102778 231367 102781
rect 228988 102776 231367 102778
rect 228988 102720 231306 102776
rect 231362 102720 231367 102776
rect 228988 102718 231367 102720
rect 231301 102715 231367 102718
rect 381629 102778 381695 102781
rect 397494 102778 397500 102780
rect 381629 102776 397500 102778
rect 381629 102720 381634 102776
rect 381690 102720 397500 102776
rect 381629 102718 397500 102720
rect 381629 102715 381695 102718
rect 397494 102716 397500 102718
rect 397564 102778 397570 102780
rect 397564 102718 400108 102778
rect 397564 102716 397570 102718
rect 265065 102642 265131 102645
rect 265065 102640 268180 102642
rect 265065 102584 265070 102640
rect 265126 102584 268180 102640
rect 265065 102582 268180 102584
rect 265065 102579 265131 102582
rect 170324 102446 217058 102506
rect 170324 102444 170330 102446
rect 67633 102370 67699 102373
rect 68142 102370 68816 102376
rect 439454 102373 439514 102748
rect 230749 102370 230815 102373
rect 67633 102368 68816 102370
rect 67633 102312 67638 102368
rect 67694 102316 68816 102368
rect 228988 102368 230815 102370
rect 67694 102312 68202 102316
rect 67633 102310 68202 102312
rect 228988 102312 230754 102368
rect 230810 102312 230815 102368
rect 228988 102310 230815 102312
rect 67633 102307 67699 102310
rect 230749 102307 230815 102310
rect 258758 102308 258764 102372
rect 258828 102370 258834 102372
rect 258828 102310 268210 102370
rect 279956 102310 287070 102370
rect 439454 102368 439563 102373
rect 439454 102312 439502 102368
rect 439558 102312 439563 102368
rect 439454 102310 439563 102312
rect 258828 102308 258834 102310
rect 213913 102234 213979 102237
rect 231301 102234 231367 102237
rect 237966 102234 237972 102236
rect 213913 102232 217028 102234
rect 213913 102176 213918 102232
rect 213974 102176 217028 102232
rect 213913 102174 217028 102176
rect 231301 102232 237972 102234
rect 231301 102176 231306 102232
rect 231362 102176 237972 102232
rect 231301 102174 237972 102176
rect 213913 102171 213979 102174
rect 231301 102171 231367 102174
rect 237966 102172 237972 102174
rect 238036 102172 238042 102236
rect 255957 102234 256023 102237
rect 257337 102234 257403 102237
rect 255957 102232 257403 102234
rect 255957 102176 255962 102232
rect 256018 102176 257342 102232
rect 257398 102176 257403 102232
rect 268150 102204 268210 102310
rect 287010 102234 287070 102310
rect 439497 102307 439563 102310
rect 290590 102234 290596 102236
rect 255957 102174 257403 102176
rect 287010 102174 290596 102234
rect 255957 102171 256023 102174
rect 257337 102171 257403 102174
rect 290590 102172 290596 102174
rect 290660 102172 290666 102236
rect 398189 102098 398255 102101
rect 398189 102096 400108 102098
rect 398189 102040 398194 102096
rect 398250 102040 400108 102096
rect 398189 102038 400108 102040
rect 398189 102035 398255 102038
rect 230565 101826 230631 101829
rect 228988 101824 230631 101826
rect 228988 101768 230570 101824
rect 230626 101768 230631 101824
rect 228988 101766 230631 101768
rect 230565 101763 230631 101766
rect 264094 101764 264100 101828
rect 264164 101826 264170 101828
rect 264164 101766 268180 101826
rect 264164 101764 264170 101766
rect 439270 101693 439330 102068
rect 439270 101688 439379 101693
rect 214005 101554 214071 101557
rect 231485 101554 231551 101557
rect 261661 101554 261727 101557
rect 214005 101552 217028 101554
rect 214005 101496 214010 101552
rect 214066 101496 217028 101552
rect 214005 101494 217028 101496
rect 231485 101552 261727 101554
rect 231485 101496 231490 101552
rect 231546 101496 261666 101552
rect 261722 101496 261727 101552
rect 231485 101494 261727 101496
rect 214005 101491 214071 101494
rect 231485 101491 231551 101494
rect 261661 101491 261727 101494
rect 231393 101418 231459 101421
rect 228988 101416 231459 101418
rect 228988 101360 231398 101416
rect 231454 101360 231459 101416
rect 228988 101358 231459 101360
rect 231393 101355 231459 101358
rect 264973 101282 265039 101285
rect 264973 101280 268180 101282
rect 264973 101224 264978 101280
rect 265034 101224 268180 101280
rect 264973 101222 268180 101224
rect 264973 101219 265039 101222
rect 213913 101010 213979 101013
rect 279926 101010 279986 101660
rect 439270 101632 439318 101688
rect 439374 101632 439379 101688
rect 439270 101630 439379 101632
rect 439313 101627 439379 101630
rect 293217 101418 293283 101421
rect 293217 101416 296730 101418
rect 293217 101360 293222 101416
rect 293278 101360 296730 101416
rect 293217 101358 296730 101360
rect 293217 101355 293283 101358
rect 296670 101146 296730 101358
rect 400078 101146 400138 101388
rect 296670 101086 400138 101146
rect 287094 101010 287100 101012
rect 213913 101008 217028 101010
rect 213913 100952 213918 101008
rect 213974 100952 217028 101008
rect 213913 100950 217028 100952
rect 279926 100950 287100 101010
rect 213913 100947 213979 100950
rect 287094 100948 287100 100950
rect 287164 100948 287170 101012
rect 231577 100874 231643 100877
rect 228988 100872 231643 100874
rect 228988 100816 231582 100872
rect 231638 100816 231643 100872
rect 228988 100814 231643 100816
rect 231577 100811 231643 100814
rect 265157 100874 265223 100877
rect 280521 100874 280587 100877
rect 265157 100872 268180 100874
rect 265157 100816 265162 100872
rect 265218 100816 268180 100872
rect 265157 100814 268180 100816
rect 279956 100872 280587 100874
rect 279956 100816 280526 100872
rect 280582 100816 280587 100872
rect 279956 100814 280587 100816
rect 265157 100811 265223 100814
rect 280521 100811 280587 100814
rect 292573 100874 292639 100877
rect 293217 100874 293283 100877
rect 292573 100872 293283 100874
rect 292573 100816 292578 100872
rect 292634 100816 293222 100872
rect 293278 100816 293283 100872
rect 292573 100814 293283 100816
rect 292573 100811 292639 100814
rect 293217 100811 293283 100814
rect 397453 100874 397519 100877
rect 442165 100874 442231 100877
rect 397453 100872 400108 100874
rect 397453 100816 397458 100872
rect 397514 100816 400108 100872
rect 397453 100814 400108 100816
rect 439852 100872 442231 100874
rect 439852 100816 442170 100872
rect 442226 100816 442231 100872
rect 439852 100814 442231 100816
rect 397453 100811 397519 100814
rect 442165 100811 442231 100814
rect 67541 100738 67607 100741
rect 68142 100738 68816 100744
rect 67541 100736 68816 100738
rect 67541 100680 67546 100736
rect 67602 100684 68816 100736
rect 230933 100738 230999 100741
rect 244222 100738 244228 100740
rect 230933 100736 244228 100738
rect 67602 100680 68202 100684
rect 67541 100678 68202 100680
rect 230933 100680 230938 100736
rect 230994 100680 244228 100736
rect 230933 100678 244228 100680
rect 67541 100675 67607 100678
rect 230933 100675 230999 100678
rect 244222 100676 244228 100678
rect 244292 100676 244298 100740
rect 231761 100466 231827 100469
rect 228988 100464 231827 100466
rect 228988 100408 231766 100464
rect 231822 100408 231827 100464
rect 228988 100406 231827 100408
rect 231761 100403 231827 100406
rect 214925 100330 214991 100333
rect 214925 100328 217028 100330
rect 214925 100272 214930 100328
rect 214986 100272 217028 100328
rect 214925 100270 217028 100272
rect 214925 100267 214991 100270
rect 260230 100132 260236 100196
rect 260300 100194 260306 100196
rect 268150 100194 268210 100436
rect 442901 100194 442967 100197
rect 260300 100134 268210 100194
rect 439852 100192 442967 100194
rect 260300 100132 260306 100134
rect 197997 100058 198063 100061
rect 216305 100058 216371 100061
rect 197997 100056 216371 100058
rect 197997 100000 198002 100056
rect 198058 100000 216310 100056
rect 216366 100000 216371 100056
rect 197997 99998 216371 100000
rect 197997 99995 198063 99998
rect 216305 99995 216371 99998
rect 264973 100058 265039 100061
rect 264973 100056 268180 100058
rect 264973 100000 264978 100056
rect 265034 100000 268180 100056
rect 264973 99998 268180 100000
rect 264973 99995 265039 99998
rect 231669 99922 231735 99925
rect 228988 99920 231735 99922
rect 228988 99864 231674 99920
rect 231730 99864 231735 99920
rect 228988 99862 231735 99864
rect 231669 99859 231735 99862
rect 279374 99653 279434 100164
rect 439852 100136 442906 100192
rect 442962 100136 442967 100192
rect 439852 100134 442967 100136
rect 442901 100131 442967 100134
rect 412398 99860 412404 99924
rect 412468 99922 412474 99924
rect 413553 99922 413619 99925
rect 412468 99920 413619 99922
rect 412468 99864 413558 99920
rect 413614 99864 413619 99920
rect 412468 99862 413619 99864
rect 412468 99860 412474 99862
rect 413553 99859 413619 99862
rect 414238 99860 414244 99924
rect 414308 99922 414314 99924
rect 414841 99922 414907 99925
rect 414308 99920 414907 99922
rect 414308 99864 414846 99920
rect 414902 99864 414907 99920
rect 414308 99862 414907 99864
rect 414308 99860 414314 99862
rect 414841 99859 414907 99862
rect 433374 99860 433380 99924
rect 433444 99922 433450 99924
rect 433517 99922 433583 99925
rect 433444 99920 433583 99922
rect 433444 99864 433522 99920
rect 433578 99864 433583 99920
rect 433444 99862 433583 99864
rect 433444 99860 433450 99862
rect 433517 99859 433583 99862
rect 434805 99922 434871 99925
rect 435030 99922 435036 99924
rect 434805 99920 435036 99922
rect 434805 99864 434810 99920
rect 434866 99864 435036 99920
rect 434805 99862 435036 99864
rect 434805 99859 434871 99862
rect 435030 99860 435036 99862
rect 435100 99860 435106 99924
rect 213913 99650 213979 99653
rect 213913 99648 217028 99650
rect 213913 99592 213918 99648
rect 213974 99592 217028 99648
rect 213913 99590 217028 99592
rect 258030 99590 268180 99650
rect 279374 99648 279483 99653
rect 279374 99592 279422 99648
rect 279478 99592 279483 99648
rect 279374 99590 279483 99592
rect 213913 99587 213979 99590
rect 230933 99514 230999 99517
rect 228988 99512 230999 99514
rect 228988 99456 230938 99512
rect 230994 99456 230999 99512
rect 228988 99454 230999 99456
rect 230933 99451 230999 99454
rect 245009 99514 245075 99517
rect 258030 99514 258090 99590
rect 279417 99587 279483 99590
rect 245009 99512 258090 99514
rect 245009 99456 245014 99512
rect 245070 99456 258090 99512
rect 245009 99454 258090 99456
rect 245009 99451 245075 99454
rect 279366 99452 279372 99516
rect 279436 99452 279442 99516
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 279374 99348 279434 99452
rect 580165 99451 580231 99454
rect 376017 99378 376083 99381
rect 404537 99378 404603 99381
rect 376017 99376 404603 99378
rect 376017 99320 376022 99376
rect 376078 99320 404542 99376
rect 404598 99320 404603 99376
rect 583520 99364 584960 99454
rect 376017 99318 404603 99320
rect 376017 99315 376083 99318
rect 404537 99315 404603 99318
rect 214005 98970 214071 98973
rect 231761 98970 231827 98973
rect 265065 98970 265131 98973
rect 214005 98968 217028 98970
rect 214005 98912 214010 98968
rect 214066 98912 217028 98968
rect 214005 98910 217028 98912
rect 228988 98968 231827 98970
rect 228988 98912 231766 98968
rect 231822 98912 231827 98968
rect 228988 98910 231827 98912
rect 214005 98907 214071 98910
rect 231761 98907 231827 98910
rect 258030 98968 265131 98970
rect 258030 98912 265070 98968
rect 265126 98912 265131 98968
rect 258030 98910 265131 98912
rect 187049 98698 187115 98701
rect 216673 98698 216739 98701
rect 187049 98696 216739 98698
rect 187049 98640 187054 98696
rect 187110 98640 216678 98696
rect 216734 98640 216739 98696
rect 187049 98638 216739 98640
rect 187049 98635 187115 98638
rect 216673 98635 216739 98638
rect 231117 98698 231183 98701
rect 258030 98698 258090 98910
rect 265065 98907 265131 98910
rect 268150 98834 268210 99212
rect 400254 99180 400260 99244
rect 400324 99242 400330 99244
rect 421925 99242 421991 99245
rect 400324 99240 421991 99242
rect 400324 99184 421930 99240
rect 421986 99184 421991 99240
rect 400324 99182 421991 99184
rect 400324 99180 400330 99182
rect 421925 99179 421991 99182
rect 419993 99106 420059 99109
rect 583661 99106 583727 99109
rect 419993 99104 583727 99106
rect 419993 99048 419998 99104
rect 420054 99048 583666 99104
rect 583722 99048 583727 99104
rect 419993 99046 583727 99048
rect 419993 99043 420059 99046
rect 583661 99043 583727 99046
rect 231117 98696 258090 98698
rect 231117 98640 231122 98696
rect 231178 98640 258090 98696
rect 231117 98638 258090 98640
rect 262814 98774 268210 98834
rect 231117 98635 231183 98638
rect 231301 98562 231367 98565
rect 228988 98560 231367 98562
rect 228988 98504 231306 98560
rect 231362 98504 231367 98560
rect 228988 98502 231367 98504
rect 231301 98499 231367 98502
rect 250437 98426 250503 98429
rect 262814 98426 262874 98774
rect 264973 98698 265039 98701
rect 264973 98696 268180 98698
rect 264973 98640 264978 98696
rect 265034 98640 268180 98696
rect 264973 98638 268180 98640
rect 264973 98635 265039 98638
rect 280153 98562 280219 98565
rect 279956 98560 280219 98562
rect 279956 98504 280158 98560
rect 280214 98504 280219 98560
rect 279956 98502 280219 98504
rect 280153 98499 280219 98502
rect 250437 98424 262874 98426
rect 250437 98368 250442 98424
rect 250498 98368 262874 98424
rect 250437 98366 262874 98368
rect 250437 98363 250503 98366
rect 213913 98290 213979 98293
rect 265709 98290 265775 98293
rect 213913 98288 217028 98290
rect 213913 98232 213918 98288
rect 213974 98232 217028 98288
rect 213913 98230 217028 98232
rect 265709 98288 268180 98290
rect 265709 98232 265714 98288
rect 265770 98232 268180 98288
rect 265709 98230 268180 98232
rect 213913 98227 213979 98230
rect 265709 98227 265775 98230
rect 231669 98018 231735 98021
rect 228988 98016 231735 98018
rect 228988 97960 231674 98016
rect 231730 97960 231735 98016
rect 228988 97958 231735 97960
rect 231669 97955 231735 97958
rect 264973 97882 265039 97885
rect 281993 97882 282059 97885
rect 264973 97880 268180 97882
rect 264973 97824 264978 97880
rect 265034 97824 268180 97880
rect 264973 97822 268180 97824
rect 279956 97880 282059 97882
rect 279956 97824 281998 97880
rect 282054 97824 282059 97880
rect 279956 97822 282059 97824
rect 264973 97819 265039 97822
rect 281993 97819 282059 97822
rect 291193 97882 291259 97885
rect 291694 97882 291700 97884
rect 291193 97880 291700 97882
rect 291193 97824 291198 97880
rect 291254 97824 291700 97880
rect 291193 97822 291700 97824
rect 291193 97819 291259 97822
rect 291694 97820 291700 97822
rect 291764 97882 291770 97884
rect 400029 97882 400095 97885
rect 434805 97884 434871 97885
rect 434805 97882 434852 97884
rect 291764 97880 400095 97882
rect 291764 97824 400034 97880
rect 400090 97824 400095 97880
rect 291764 97822 400095 97824
rect 434760 97880 434852 97882
rect 434760 97824 434810 97880
rect 434760 97822 434852 97824
rect 291764 97820 291770 97822
rect 400029 97819 400095 97822
rect 434805 97820 434852 97822
rect 434916 97820 434922 97884
rect 437381 97882 437447 97885
rect 448605 97882 448671 97885
rect 437381 97880 448671 97882
rect 437381 97824 437386 97880
rect 437442 97824 448610 97880
rect 448666 97824 448671 97880
rect 437381 97822 448671 97824
rect 434805 97819 434871 97820
rect 437381 97819 437447 97822
rect 448605 97819 448671 97822
rect 381537 97746 381603 97749
rect 431585 97746 431651 97749
rect 381537 97744 431970 97746
rect -960 97610 480 97700
rect 381537 97688 381542 97744
rect 381598 97688 431590 97744
rect 431646 97688 431970 97744
rect 381537 97686 431970 97688
rect 381537 97683 381603 97686
rect 431585 97683 431651 97686
rect 3509 97610 3575 97613
rect 231485 97610 231551 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect 228988 97608 231551 97610
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 174721 97066 174787 97069
rect 216998 97066 217058 97580
rect 228988 97552 231490 97608
rect 231546 97552 231551 97608
rect 228988 97550 231551 97552
rect 231485 97547 231551 97550
rect 264513 97474 264579 97477
rect 264513 97472 268180 97474
rect 264513 97416 264518 97472
rect 264574 97416 268180 97472
rect 264513 97414 268180 97416
rect 264513 97411 264579 97414
rect 414657 97202 414723 97205
rect 423857 97202 423923 97205
rect 414657 97200 423923 97202
rect 414657 97144 414662 97200
rect 414718 97144 423862 97200
rect 423918 97144 423923 97200
rect 414657 97142 423923 97144
rect 431910 97202 431970 97686
rect 582465 97202 582531 97205
rect 431910 97200 582531 97202
rect 431910 97144 582470 97200
rect 582526 97144 582531 97200
rect 431910 97142 582531 97144
rect 414657 97139 414723 97142
rect 423857 97139 423923 97142
rect 582465 97139 582531 97142
rect 229134 97066 229140 97068
rect 174721 97064 217058 97066
rect 174721 97008 174726 97064
rect 174782 97008 217058 97064
rect 174721 97006 217058 97008
rect 228988 97006 229140 97066
rect 174721 97003 174787 97006
rect 229134 97004 229140 97006
rect 229204 97066 229210 97068
rect 231761 97066 231827 97069
rect 425697 97066 425763 97069
rect 427721 97066 427787 97069
rect 229204 97064 231827 97066
rect 229204 97008 231766 97064
rect 231822 97008 231827 97064
rect 229204 97006 231827 97008
rect 229204 97004 229210 97006
rect 231761 97003 231827 97006
rect 258030 97006 268180 97066
rect 425697 97064 427787 97066
rect 213913 96930 213979 96933
rect 258030 96930 258090 97006
rect 213913 96928 217028 96930
rect 213913 96872 213918 96928
rect 213974 96872 217028 96928
rect 213913 96870 217028 96872
rect 238710 96870 258090 96930
rect 213913 96867 213979 96870
rect 229134 96732 229140 96796
rect 229204 96794 229210 96796
rect 238710 96794 238770 96870
rect 229204 96734 238770 96794
rect 229204 96732 229210 96734
rect 279374 96661 279434 97036
rect 425697 97008 425702 97064
rect 425758 97008 427726 97064
rect 427782 97008 427787 97064
rect 425697 97006 427787 97008
rect 425697 97003 425763 97006
rect 427721 97003 427787 97006
rect 400857 96930 400923 96933
rect 402605 96930 402671 96933
rect 400857 96928 402671 96930
rect 400857 96872 400862 96928
rect 400918 96872 402610 96928
rect 402666 96872 402671 96928
rect 400857 96870 402671 96872
rect 400857 96867 400923 96870
rect 402605 96867 402671 96870
rect 427077 96930 427143 96933
rect 427905 96930 427971 96933
rect 427077 96928 427971 96930
rect 427077 96872 427082 96928
rect 427138 96872 427910 96928
rect 427966 96872 427971 96928
rect 427077 96870 427971 96872
rect 427077 96867 427143 96870
rect 427905 96867 427971 96870
rect 230565 96658 230631 96661
rect 231669 96658 231735 96661
rect 228988 96656 231735 96658
rect 228988 96600 230570 96656
rect 230626 96600 231674 96656
rect 231730 96600 231735 96656
rect 228988 96598 231735 96600
rect 230565 96595 230631 96598
rect 231669 96595 231735 96598
rect 267825 96658 267891 96661
rect 267825 96656 268180 96658
rect 267825 96600 267830 96656
rect 267886 96600 268180 96656
rect 267825 96598 268180 96600
rect 279325 96656 279434 96661
rect 279325 96600 279330 96656
rect 279386 96600 279434 96656
rect 279325 96598 279434 96600
rect 267825 96595 267891 96598
rect 279325 96595 279391 96598
rect 231761 96522 231827 96525
rect 255262 96522 255268 96524
rect 231761 96520 255268 96522
rect 231761 96464 231766 96520
rect 231822 96464 255268 96520
rect 231761 96462 255268 96464
rect 231761 96459 231827 96462
rect 255262 96460 255268 96462
rect 255332 96522 255338 96524
rect 298001 96522 298067 96525
rect 418705 96522 418771 96525
rect 255332 96462 258090 96522
rect 255332 96460 255338 96462
rect 214833 96386 214899 96389
rect 214833 96384 217028 96386
rect 214833 96328 214838 96384
rect 214894 96328 217028 96384
rect 214833 96326 217028 96328
rect 214833 96323 214899 96326
rect 230473 96250 230539 96253
rect 228988 96248 230539 96250
rect 228988 96192 230478 96248
rect 230534 96192 230539 96248
rect 228988 96190 230539 96192
rect 230473 96187 230539 96190
rect 219157 95980 219223 95981
rect 219157 95978 219204 95980
rect 219112 95976 219204 95978
rect 219112 95920 219162 95976
rect 219112 95918 219204 95920
rect 219157 95916 219204 95918
rect 219268 95916 219274 95980
rect 219157 95915 219223 95916
rect 166390 95780 166396 95844
rect 166460 95842 166466 95844
rect 203609 95842 203675 95845
rect 166460 95840 203675 95842
rect 166460 95784 203614 95840
rect 203670 95784 203675 95840
rect 166460 95782 203675 95784
rect 166460 95780 166466 95782
rect 203609 95779 203675 95782
rect 204897 95842 204963 95845
rect 216029 95842 216095 95845
rect 204897 95840 216095 95842
rect 204897 95784 204902 95840
rect 204958 95784 216034 95840
rect 216090 95784 216095 95840
rect 204897 95782 216095 95784
rect 258030 95842 258090 96462
rect 298001 96520 418771 96522
rect 298001 96464 298006 96520
rect 298062 96464 418710 96520
rect 418766 96464 418771 96520
rect 298001 96462 418771 96464
rect 298001 96459 298067 96462
rect 418705 96459 418771 96462
rect 397913 96386 397979 96389
rect 405733 96386 405799 96389
rect 406469 96386 406535 96389
rect 397913 96384 406535 96386
rect 267733 95842 267799 95845
rect 258030 95840 267799 95842
rect 258030 95784 267738 95840
rect 267794 95784 267799 95840
rect 258030 95782 267799 95784
rect 204897 95779 204963 95782
rect 216029 95779 216095 95782
rect 267733 95779 267799 95782
rect 224902 95508 224908 95572
rect 224972 95570 224978 95572
rect 228950 95570 228956 95572
rect 224972 95510 228956 95570
rect 224972 95508 224978 95510
rect 228950 95508 228956 95510
rect 229020 95508 229026 95572
rect 228449 95298 228515 95301
rect 268150 95298 268210 96220
rect 279926 95842 279986 96356
rect 397913 96328 397918 96384
rect 397974 96328 405738 96384
rect 405794 96328 406474 96384
rect 406530 96328 406535 96384
rect 397913 96326 406535 96328
rect 397913 96323 397979 96326
rect 405733 96323 405799 96326
rect 406469 96323 406535 96326
rect 280061 95842 280127 95845
rect 279926 95840 280127 95842
rect 279926 95784 280066 95840
rect 280122 95784 280127 95840
rect 279926 95782 280127 95784
rect 280061 95779 280127 95782
rect 228449 95296 268210 95298
rect 228449 95240 228454 95296
rect 228510 95240 268210 95296
rect 228449 95238 268210 95240
rect 228449 95235 228515 95238
rect 205398 95100 205404 95164
rect 205468 95162 205474 95164
rect 280153 95162 280219 95165
rect 205468 95160 280219 95162
rect 205468 95104 280158 95160
rect 280214 95104 280219 95160
rect 205468 95102 280219 95104
rect 205468 95100 205474 95102
rect 280153 95099 280219 95102
rect 396901 95162 396967 95165
rect 438669 95162 438735 95165
rect 396901 95160 438735 95162
rect 396901 95104 396906 95160
rect 396962 95104 438674 95160
rect 438730 95104 438735 95160
rect 396901 95102 438735 95104
rect 396901 95099 396967 95102
rect 438669 95099 438735 95102
rect 260046 94964 260052 95028
rect 260116 95026 260122 95028
rect 279325 95026 279391 95029
rect 260116 95024 279391 95026
rect 260116 94968 279330 95024
rect 279386 94968 279391 95024
rect 260116 94966 279391 94968
rect 260116 94964 260122 94966
rect 279325 94963 279391 94966
rect 100661 94756 100727 94757
rect 120625 94756 120691 94757
rect 100624 94692 100630 94756
rect 100694 94754 100727 94756
rect 100694 94752 100786 94754
rect 100722 94696 100786 94752
rect 100694 94694 100786 94696
rect 100694 94692 100727 94694
rect 120616 94692 120622 94756
rect 120686 94754 120692 94756
rect 120686 94694 120778 94754
rect 120686 94692 120692 94694
rect 151486 94692 151492 94756
rect 151556 94754 151562 94756
rect 151760 94754 151766 94756
rect 151556 94694 151766 94754
rect 151556 94692 151562 94694
rect 151760 94692 151766 94694
rect 151830 94692 151836 94756
rect 100661 94691 100727 94692
rect 120625 94691 120691 94692
rect 66161 94482 66227 94485
rect 106917 94482 106983 94485
rect 66161 94480 106983 94482
rect 66161 94424 66166 94480
rect 66222 94424 106922 94480
rect 106978 94424 106983 94480
rect 66161 94422 106983 94424
rect 66161 94419 66227 94422
rect 106917 94419 106983 94422
rect 160737 94482 160803 94485
rect 170397 94482 170463 94485
rect 160737 94480 170463 94482
rect 160737 94424 160742 94480
rect 160798 94424 170402 94480
rect 170458 94424 170463 94480
rect 160737 94422 170463 94424
rect 160737 94419 160803 94422
rect 170397 94419 170463 94422
rect 191097 94482 191163 94485
rect 231209 94482 231275 94485
rect 191097 94480 231275 94482
rect 191097 94424 191102 94480
rect 191158 94424 231214 94480
rect 231270 94424 231275 94480
rect 191097 94422 231275 94424
rect 191097 94419 191163 94422
rect 231209 94419 231275 94422
rect 267590 94420 267596 94484
rect 267660 94482 267666 94484
rect 273345 94482 273411 94485
rect 267660 94480 273411 94482
rect 267660 94424 273350 94480
rect 273406 94424 273411 94480
rect 267660 94422 273411 94424
rect 267660 94420 267666 94422
rect 273345 94419 273411 94422
rect 122046 94012 122052 94076
rect 122116 94074 122122 94076
rect 174537 94074 174603 94077
rect 122116 94072 174603 94074
rect 122116 94016 174542 94072
rect 174598 94016 174603 94072
rect 122116 94014 174603 94016
rect 122116 94012 122122 94014
rect 174537 94011 174603 94014
rect 114318 93876 114324 93940
rect 114388 93938 114394 93940
rect 215937 93938 216003 93941
rect 114388 93936 216003 93938
rect 114388 93880 215942 93936
rect 215998 93880 216003 93936
rect 114388 93878 216003 93880
rect 114388 93876 114394 93878
rect 215937 93875 216003 93878
rect 224309 93938 224375 93941
rect 229686 93938 229692 93940
rect 224309 93936 229692 93938
rect 224309 93880 224314 93936
rect 224370 93880 229692 93936
rect 224309 93878 229692 93880
rect 224309 93875 224375 93878
rect 229686 93876 229692 93878
rect 229756 93876 229762 93940
rect 94998 93740 95004 93804
rect 95068 93802 95074 93804
rect 170765 93802 170831 93805
rect 95068 93800 170831 93802
rect 95068 93744 170770 93800
rect 170826 93744 170831 93800
rect 95068 93742 170831 93744
rect 95068 93740 95074 93742
rect 170765 93739 170831 93742
rect 201125 93802 201191 93805
rect 280061 93802 280127 93805
rect 201125 93800 280127 93802
rect 201125 93744 201130 93800
rect 201186 93744 280066 93800
rect 280122 93744 280127 93800
rect 201125 93742 280127 93744
rect 201125 93739 201191 93742
rect 280061 93739 280127 93742
rect 378869 93802 378935 93805
rect 409689 93802 409755 93805
rect 378869 93800 409755 93802
rect 378869 93744 378874 93800
rect 378930 93744 409694 93800
rect 409750 93744 409755 93800
rect 378869 93742 409755 93744
rect 378869 93739 378935 93742
rect 409689 93739 409755 93742
rect 118233 93532 118299 93533
rect 124121 93532 124187 93533
rect 118182 93530 118188 93532
rect 118142 93470 118188 93530
rect 118252 93528 118299 93532
rect 124070 93530 124076 93532
rect 118294 93472 118299 93528
rect 118182 93468 118188 93470
rect 118252 93468 118299 93472
rect 124030 93470 124076 93530
rect 124140 93528 124187 93532
rect 124182 93472 124187 93528
rect 124070 93468 124076 93470
rect 124140 93468 124187 93472
rect 118233 93467 118299 93468
rect 124121 93467 124187 93468
rect 162485 93394 162551 93397
rect 185577 93394 185643 93397
rect 162485 93392 185643 93394
rect 162485 93336 162490 93392
rect 162546 93336 185582 93392
rect 185638 93336 185643 93392
rect 162485 93334 185643 93336
rect 162485 93331 162551 93334
rect 185577 93331 185643 93334
rect 103278 93196 103284 93260
rect 103348 93258 103354 93260
rect 103421 93258 103487 93261
rect 110137 93260 110203 93261
rect 110086 93258 110092 93260
rect 103348 93256 103487 93258
rect 103348 93200 103426 93256
rect 103482 93200 103487 93256
rect 103348 93198 103487 93200
rect 110046 93198 110092 93258
rect 110156 93256 110203 93260
rect 110198 93200 110203 93256
rect 103348 93196 103354 93198
rect 103421 93195 103487 93198
rect 110086 93196 110092 93198
rect 110156 93196 110203 93200
rect 110137 93195 110203 93196
rect 162117 93258 162183 93261
rect 214925 93258 214991 93261
rect 162117 93256 214991 93258
rect 162117 93200 162122 93256
rect 162178 93200 214930 93256
rect 214986 93200 214991 93256
rect 162117 93198 214991 93200
rect 162117 93195 162183 93198
rect 214925 93195 214991 93198
rect 115790 93060 115796 93124
rect 115860 93122 115866 93124
rect 166349 93122 166415 93125
rect 115860 93120 166415 93122
rect 115860 93064 166354 93120
rect 166410 93064 166415 93120
rect 115860 93062 166415 93064
rect 115860 93060 115866 93062
rect 166349 93059 166415 93062
rect 181437 93122 181503 93125
rect 258758 93122 258764 93124
rect 181437 93120 258764 93122
rect 181437 93064 181442 93120
rect 181498 93064 258764 93120
rect 181437 93062 258764 93064
rect 181437 93059 181503 93062
rect 258758 93060 258764 93062
rect 258828 93060 258834 93124
rect 286174 93060 286180 93124
rect 286244 93122 286250 93124
rect 289813 93122 289879 93125
rect 286244 93120 289879 93122
rect 286244 93064 289818 93120
rect 289874 93064 289879 93120
rect 286244 93062 289879 93064
rect 286244 93060 286250 93062
rect 289813 93059 289879 93062
rect 412265 93122 412331 93125
rect 583109 93122 583175 93125
rect 412265 93120 583175 93122
rect 412265 93064 412270 93120
rect 412326 93064 583114 93120
rect 583170 93064 583175 93120
rect 412265 93062 583175 93064
rect 412265 93059 412331 93062
rect 583109 93059 583175 93062
rect 408493 92578 408559 92581
rect 409689 92578 409755 92581
rect 408493 92576 409755 92578
rect 408493 92520 408498 92576
rect 408554 92520 409694 92576
rect 409750 92520 409755 92576
rect 408493 92518 409755 92520
rect 408493 92515 408559 92518
rect 409689 92515 409755 92518
rect 84326 92380 84332 92444
rect 84396 92442 84402 92444
rect 85113 92442 85179 92445
rect 108113 92444 108179 92445
rect 108062 92442 108068 92444
rect 84396 92440 85179 92442
rect 84396 92384 85118 92440
rect 85174 92384 85179 92440
rect 84396 92382 85179 92384
rect 108022 92382 108068 92442
rect 108132 92440 108179 92444
rect 108174 92384 108179 92440
rect 84396 92380 84402 92382
rect 85113 92379 85179 92382
rect 108062 92380 108068 92382
rect 108132 92380 108179 92384
rect 110638 92380 110644 92444
rect 110708 92442 110714 92444
rect 111241 92442 111307 92445
rect 110708 92440 111307 92442
rect 110708 92384 111246 92440
rect 111302 92384 111307 92440
rect 110708 92382 111307 92384
rect 110708 92380 110714 92382
rect 108113 92379 108179 92380
rect 111241 92379 111307 92382
rect 114870 92380 114876 92444
rect 114940 92442 114946 92444
rect 115749 92442 115815 92445
rect 116761 92444 116827 92445
rect 125777 92444 125843 92445
rect 133137 92444 133203 92445
rect 116710 92442 116716 92444
rect 114940 92440 115815 92442
rect 114940 92384 115754 92440
rect 115810 92384 115815 92440
rect 114940 92382 115815 92384
rect 116670 92382 116716 92442
rect 116780 92440 116827 92444
rect 125726 92442 125732 92444
rect 116822 92384 116827 92440
rect 114940 92380 114946 92382
rect 115749 92379 115815 92382
rect 116710 92380 116716 92382
rect 116780 92380 116827 92384
rect 125686 92382 125732 92442
rect 125796 92440 125843 92444
rect 133086 92442 133092 92444
rect 125838 92384 125843 92440
rect 125726 92380 125732 92382
rect 125796 92380 125843 92384
rect 133046 92382 133092 92442
rect 133156 92440 133203 92444
rect 133198 92384 133203 92440
rect 133086 92380 133092 92382
rect 133156 92380 133203 92384
rect 116761 92379 116827 92380
rect 125777 92379 125843 92380
rect 133137 92379 133203 92380
rect 120206 92244 120212 92308
rect 120276 92306 120282 92308
rect 173341 92306 173407 92309
rect 120276 92304 173407 92306
rect 120276 92248 173346 92304
rect 173402 92248 173407 92304
rect 120276 92246 173407 92248
rect 120276 92244 120282 92246
rect 173341 92243 173407 92246
rect 115473 92172 115539 92173
rect 115422 92170 115428 92172
rect 115382 92110 115428 92170
rect 115492 92168 115539 92172
rect 115534 92112 115539 92168
rect 115422 92108 115428 92110
rect 115492 92108 115539 92112
rect 127566 92108 127572 92172
rect 127636 92170 127642 92172
rect 165061 92170 165127 92173
rect 127636 92168 165127 92170
rect 127636 92112 165066 92168
rect 165122 92112 165127 92168
rect 127636 92110 165127 92112
rect 127636 92108 127642 92110
rect 115473 92107 115539 92108
rect 165061 92107 165127 92110
rect 104566 91972 104572 92036
rect 104636 92034 104642 92036
rect 104636 91974 113190 92034
rect 104636 91972 104642 91974
rect 111190 91836 111196 91900
rect 111260 91898 111266 91900
rect 111333 91898 111399 91901
rect 111260 91896 111399 91898
rect 111260 91840 111338 91896
rect 111394 91840 111399 91896
rect 111260 91838 111399 91840
rect 113130 91898 113190 91974
rect 116577 91898 116643 91901
rect 120717 91898 120783 91901
rect 113130 91896 116643 91898
rect 113130 91840 116582 91896
rect 116638 91840 116643 91896
rect 113130 91838 116643 91840
rect 111260 91836 111266 91838
rect 111333 91835 111399 91838
rect 116577 91835 116643 91838
rect 116902 91896 120783 91898
rect 116902 91840 120722 91896
rect 120778 91840 120783 91896
rect 116902 91838 120783 91840
rect 100886 91700 100892 91764
rect 100956 91762 100962 91764
rect 116902 91762 116962 91838
rect 120717 91835 120783 91838
rect 206461 91898 206527 91901
rect 276013 91898 276079 91901
rect 206461 91896 276079 91898
rect 206461 91840 206466 91896
rect 206522 91840 276018 91896
rect 276074 91840 276079 91896
rect 206461 91838 276079 91840
rect 206461 91835 206527 91838
rect 276013 91835 276079 91838
rect 100956 91702 116962 91762
rect 100956 91700 100962 91702
rect 119654 91700 119660 91764
rect 119724 91762 119730 91764
rect 119889 91762 119955 91765
rect 130745 91764 130811 91765
rect 130694 91762 130700 91764
rect 119724 91760 119955 91762
rect 119724 91704 119894 91760
rect 119950 91704 119955 91760
rect 119724 91702 119955 91704
rect 130654 91702 130700 91762
rect 130764 91760 130811 91764
rect 130806 91704 130811 91760
rect 119724 91700 119730 91702
rect 119889 91699 119955 91702
rect 130694 91700 130700 91702
rect 130764 91700 130811 91704
rect 151302 91700 151308 91764
rect 151372 91762 151378 91764
rect 151629 91762 151695 91765
rect 151372 91760 151695 91762
rect 151372 91704 151634 91760
rect 151690 91704 151695 91760
rect 151372 91702 151695 91704
rect 151372 91700 151378 91702
rect 130745 91699 130811 91700
rect 151629 91699 151695 91702
rect 170397 91762 170463 91765
rect 265801 91762 265867 91765
rect 170397 91760 265867 91762
rect 170397 91704 170402 91760
rect 170458 91704 265806 91760
rect 265862 91704 265867 91760
rect 170397 91702 265867 91704
rect 170397 91699 170463 91702
rect 265801 91699 265867 91702
rect 286317 91762 286383 91765
rect 418061 91762 418127 91765
rect 286317 91760 418127 91762
rect 286317 91704 286322 91760
rect 286378 91704 418066 91760
rect 418122 91704 418127 91760
rect 286317 91702 418127 91704
rect 286317 91699 286383 91702
rect 418061 91699 418127 91702
rect 113214 91564 113220 91628
rect 113284 91626 113290 91628
rect 177481 91626 177547 91629
rect 113284 91624 177547 91626
rect 113284 91568 177486 91624
rect 177542 91568 177547 91624
rect 113284 91566 177547 91568
rect 113284 91564 113290 91566
rect 177481 91563 177547 91566
rect 99046 91428 99052 91492
rect 99116 91490 99122 91492
rect 104157 91490 104223 91493
rect 99116 91488 104223 91490
rect 99116 91432 104162 91488
rect 104218 91432 104223 91488
rect 99116 91430 104223 91432
rect 99116 91428 99122 91430
rect 104157 91427 104223 91430
rect 122782 91428 122788 91492
rect 122852 91490 122858 91492
rect 124029 91490 124095 91493
rect 122852 91488 124095 91490
rect 122852 91432 124034 91488
rect 124090 91432 124095 91488
rect 122852 91430 124095 91432
rect 122852 91428 122858 91430
rect 124029 91427 124095 91430
rect 85798 91292 85804 91356
rect 85868 91354 85874 91356
rect 86861 91354 86927 91357
rect 85868 91352 86927 91354
rect 85868 91296 86866 91352
rect 86922 91296 86927 91352
rect 85868 91294 86927 91296
rect 85868 91292 85874 91294
rect 86861 91291 86927 91294
rect 96654 91292 96660 91356
rect 96724 91354 96730 91356
rect 97809 91354 97875 91357
rect 96724 91352 97875 91354
rect 96724 91296 97814 91352
rect 97870 91296 97875 91352
rect 96724 91294 97875 91296
rect 96724 91292 96730 91294
rect 97809 91291 97875 91294
rect 101806 91292 101812 91356
rect 101876 91354 101882 91356
rect 101949 91354 102015 91357
rect 101876 91352 102015 91354
rect 101876 91296 101954 91352
rect 102010 91296 102015 91352
rect 101876 91294 102015 91296
rect 101876 91292 101882 91294
rect 101949 91291 102015 91294
rect 105486 91292 105492 91356
rect 105556 91354 105562 91356
rect 106181 91354 106247 91357
rect 105556 91352 106247 91354
rect 105556 91296 106186 91352
rect 106242 91296 106247 91352
rect 105556 91294 106247 91296
rect 105556 91292 105562 91294
rect 106181 91291 106247 91294
rect 106406 91292 106412 91356
rect 106476 91354 106482 91356
rect 107561 91354 107627 91357
rect 106476 91352 107627 91354
rect 106476 91296 107566 91352
rect 107622 91296 107627 91352
rect 106476 91294 107627 91296
rect 106476 91292 106482 91294
rect 107561 91291 107627 91294
rect 126462 91292 126468 91356
rect 126532 91354 126538 91356
rect 126789 91354 126855 91357
rect 151537 91356 151603 91357
rect 151486 91354 151492 91356
rect 126532 91352 126855 91354
rect 126532 91296 126794 91352
rect 126850 91296 126855 91352
rect 126532 91294 126855 91296
rect 151446 91294 151492 91354
rect 151556 91352 151603 91356
rect 151598 91296 151603 91352
rect 126532 91292 126538 91294
rect 126789 91291 126855 91294
rect 151486 91292 151492 91294
rect 151556 91292 151603 91296
rect 151537 91291 151603 91292
rect 74758 91156 74764 91220
rect 74828 91218 74834 91220
rect 75269 91218 75335 91221
rect 86769 91220 86835 91221
rect 88057 91220 88123 91221
rect 86718 91218 86724 91220
rect 74828 91216 75335 91218
rect 74828 91160 75274 91216
rect 75330 91160 75335 91216
rect 74828 91158 75335 91160
rect 86678 91158 86724 91218
rect 86788 91216 86835 91220
rect 88006 91218 88012 91220
rect 86830 91160 86835 91216
rect 74828 91156 74834 91158
rect 75269 91155 75335 91158
rect 86718 91156 86724 91158
rect 86788 91156 86835 91160
rect 87966 91158 88012 91218
rect 88076 91216 88123 91220
rect 88118 91160 88123 91216
rect 88006 91156 88012 91158
rect 88076 91156 88123 91160
rect 88926 91156 88932 91220
rect 88996 91218 89002 91220
rect 89621 91218 89687 91221
rect 88996 91216 89687 91218
rect 88996 91160 89626 91216
rect 89682 91160 89687 91216
rect 88996 91158 89687 91160
rect 88996 91156 89002 91158
rect 86769 91155 86835 91156
rect 88057 91155 88123 91156
rect 89621 91155 89687 91158
rect 90214 91156 90220 91220
rect 90284 91218 90290 91220
rect 90725 91218 90791 91221
rect 90284 91216 90791 91218
rect 90284 91160 90730 91216
rect 90786 91160 90791 91216
rect 90284 91158 90791 91160
rect 90284 91156 90290 91158
rect 90725 91155 90791 91158
rect 91318 91156 91324 91220
rect 91388 91218 91394 91220
rect 91921 91218 91987 91221
rect 91388 91216 91987 91218
rect 91388 91160 91926 91216
rect 91982 91160 91987 91216
rect 91388 91158 91987 91160
rect 91388 91156 91394 91158
rect 91921 91155 91987 91158
rect 92606 91156 92612 91220
rect 92676 91218 92682 91220
rect 93025 91218 93091 91221
rect 92676 91216 93091 91218
rect 92676 91160 93030 91216
rect 93086 91160 93091 91216
rect 92676 91158 93091 91160
rect 92676 91156 92682 91158
rect 93025 91155 93091 91158
rect 93894 91156 93900 91220
rect 93964 91218 93970 91220
rect 95141 91218 95207 91221
rect 96337 91220 96403 91221
rect 96286 91218 96292 91220
rect 93964 91216 95207 91218
rect 93964 91160 95146 91216
rect 95202 91160 95207 91216
rect 93964 91158 95207 91160
rect 96246 91158 96292 91218
rect 96356 91216 96403 91220
rect 96398 91160 96403 91216
rect 93964 91156 93970 91158
rect 95141 91155 95207 91158
rect 96286 91156 96292 91158
rect 96356 91156 96403 91160
rect 97206 91156 97212 91220
rect 97276 91218 97282 91220
rect 97901 91218 97967 91221
rect 97276 91216 97967 91218
rect 97276 91160 97906 91216
rect 97962 91160 97967 91216
rect 97276 91158 97967 91160
rect 97276 91156 97282 91158
rect 96337 91155 96403 91156
rect 97901 91155 97967 91158
rect 98126 91156 98132 91220
rect 98196 91218 98202 91220
rect 99189 91218 99255 91221
rect 98196 91216 99255 91218
rect 98196 91160 99194 91216
rect 99250 91160 99255 91216
rect 98196 91158 99255 91160
rect 98196 91156 98202 91158
rect 99189 91155 99255 91158
rect 99966 91156 99972 91220
rect 100036 91218 100042 91220
rect 100661 91218 100727 91221
rect 102041 91220 102107 91221
rect 101990 91218 101996 91220
rect 100036 91216 100727 91218
rect 100036 91160 100666 91216
rect 100722 91160 100727 91216
rect 100036 91158 100727 91160
rect 101950 91158 101996 91218
rect 102060 91216 102107 91220
rect 102102 91160 102107 91216
rect 100036 91156 100042 91158
rect 100661 91155 100727 91158
rect 101990 91156 101996 91158
rect 102060 91156 102107 91160
rect 102726 91156 102732 91220
rect 102796 91218 102802 91220
rect 103329 91218 103395 91221
rect 102796 91216 103395 91218
rect 102796 91160 103334 91216
rect 103390 91160 103395 91216
rect 102796 91158 103395 91160
rect 102796 91156 102802 91158
rect 102041 91155 102107 91156
rect 103329 91155 103395 91158
rect 104198 91156 104204 91220
rect 104268 91218 104274 91220
rect 104433 91218 104499 91221
rect 104268 91216 104499 91218
rect 104268 91160 104438 91216
rect 104494 91160 104499 91216
rect 104268 91158 104499 91160
rect 104268 91156 104274 91158
rect 104433 91155 104499 91158
rect 105670 91156 105676 91220
rect 105740 91218 105746 91220
rect 106089 91218 106155 91221
rect 105740 91216 106155 91218
rect 105740 91160 106094 91216
rect 106150 91160 106155 91216
rect 105740 91158 106155 91160
rect 105740 91156 105746 91158
rect 106089 91155 106155 91158
rect 106774 91156 106780 91220
rect 106844 91218 106850 91220
rect 107469 91218 107535 91221
rect 106844 91216 107535 91218
rect 106844 91160 107474 91216
rect 107530 91160 107535 91216
rect 106844 91158 107535 91160
rect 106844 91156 106850 91158
rect 107469 91155 107535 91158
rect 107694 91156 107700 91220
rect 107764 91218 107770 91220
rect 108665 91218 108731 91221
rect 109217 91220 109283 91221
rect 109166 91218 109172 91220
rect 107764 91216 108731 91218
rect 107764 91160 108670 91216
rect 108726 91160 108731 91216
rect 107764 91158 108731 91160
rect 109126 91158 109172 91218
rect 109236 91216 109283 91220
rect 109278 91160 109283 91216
rect 107764 91156 107770 91158
rect 108665 91155 108731 91158
rect 109166 91156 109172 91158
rect 109236 91156 109283 91160
rect 109534 91156 109540 91220
rect 109604 91218 109610 91220
rect 110137 91218 110203 91221
rect 109604 91216 110203 91218
rect 109604 91160 110142 91216
rect 110198 91160 110203 91216
rect 109604 91158 110203 91160
rect 109604 91156 109610 91158
rect 109217 91155 109283 91156
rect 110137 91155 110203 91158
rect 111926 91156 111932 91220
rect 111996 91218 112002 91220
rect 112161 91218 112227 91221
rect 111996 91216 112227 91218
rect 111996 91160 112166 91216
rect 112222 91160 112227 91216
rect 111996 91158 112227 91160
rect 111996 91156 112002 91158
rect 112161 91155 112227 91158
rect 112294 91156 112300 91220
rect 112364 91218 112370 91220
rect 113081 91218 113147 91221
rect 114369 91220 114435 91221
rect 117129 91220 117195 91221
rect 118049 91220 118115 91221
rect 114318 91218 114324 91220
rect 112364 91216 113147 91218
rect 112364 91160 113086 91216
rect 113142 91160 113147 91216
rect 112364 91158 113147 91160
rect 114278 91158 114324 91218
rect 114388 91216 114435 91220
rect 117078 91218 117084 91220
rect 114430 91160 114435 91216
rect 112364 91156 112370 91158
rect 113081 91155 113147 91158
rect 114318 91156 114324 91158
rect 114388 91156 114435 91160
rect 117038 91158 117084 91218
rect 117148 91216 117195 91220
rect 117998 91218 118004 91220
rect 117190 91160 117195 91216
rect 117078 91156 117084 91158
rect 117148 91156 117195 91160
rect 117958 91158 118004 91218
rect 118068 91216 118115 91220
rect 118110 91160 118115 91216
rect 117998 91156 118004 91158
rect 118068 91156 118115 91160
rect 119286 91156 119292 91220
rect 119356 91218 119362 91220
rect 119981 91218 120047 91221
rect 119356 91216 120047 91218
rect 119356 91160 119986 91216
rect 120042 91160 120047 91216
rect 119356 91158 120047 91160
rect 119356 91156 119362 91158
rect 114369 91155 114435 91156
rect 117129 91155 117195 91156
rect 118049 91155 118115 91156
rect 119981 91155 120047 91158
rect 121678 91156 121684 91220
rect 121748 91218 121754 91220
rect 122281 91218 122347 91221
rect 121748 91216 122347 91218
rect 121748 91160 122286 91216
rect 122342 91160 122347 91216
rect 121748 91158 122347 91160
rect 121748 91156 121754 91158
rect 122281 91155 122347 91158
rect 123150 91156 123156 91220
rect 123220 91218 123226 91220
rect 124121 91218 124187 91221
rect 125409 91220 125475 91221
rect 125358 91218 125364 91220
rect 123220 91216 124187 91218
rect 123220 91160 124126 91216
rect 124182 91160 124187 91216
rect 123220 91158 124187 91160
rect 125318 91158 125364 91218
rect 125428 91216 125475 91220
rect 125470 91160 125475 91216
rect 123220 91156 123226 91158
rect 124121 91155 124187 91158
rect 125358 91156 125364 91158
rect 125428 91156 125475 91160
rect 126646 91156 126652 91220
rect 126716 91218 126722 91220
rect 126881 91218 126947 91221
rect 126716 91216 126947 91218
rect 126716 91160 126886 91216
rect 126942 91160 126947 91216
rect 126716 91158 126947 91160
rect 126716 91156 126722 91158
rect 125409 91155 125475 91156
rect 126881 91155 126947 91158
rect 129406 91156 129412 91220
rect 129476 91218 129482 91220
rect 129641 91218 129707 91221
rect 132401 91220 132467 91221
rect 132350 91218 132356 91220
rect 129476 91216 129707 91218
rect 129476 91160 129646 91216
rect 129702 91160 129707 91216
rect 129476 91158 129707 91160
rect 132310 91158 132356 91218
rect 132420 91216 132467 91220
rect 132462 91160 132467 91216
rect 129476 91156 129482 91158
rect 129641 91155 129707 91158
rect 132350 91156 132356 91158
rect 132420 91156 132467 91160
rect 134374 91156 134380 91220
rect 134444 91218 134450 91220
rect 135161 91218 135227 91221
rect 134444 91216 135227 91218
rect 134444 91160 135166 91216
rect 135222 91160 135227 91216
rect 134444 91158 135227 91160
rect 134444 91156 134450 91158
rect 132401 91155 132467 91156
rect 135161 91155 135227 91158
rect 136030 91156 136036 91220
rect 136100 91218 136106 91220
rect 136541 91218 136607 91221
rect 151721 91220 151787 91221
rect 151670 91218 151676 91220
rect 136100 91216 136607 91218
rect 136100 91160 136546 91216
rect 136602 91160 136607 91216
rect 136100 91158 136607 91160
rect 151630 91158 151676 91218
rect 151740 91216 151787 91220
rect 151782 91160 151787 91216
rect 136100 91156 136106 91158
rect 136541 91155 136607 91158
rect 151670 91156 151676 91158
rect 151740 91156 151787 91160
rect 152038 91156 152044 91220
rect 152108 91218 152114 91220
rect 153101 91218 153167 91221
rect 152108 91216 153167 91218
rect 152108 91160 153106 91216
rect 153162 91160 153167 91216
rect 152108 91158 153167 91160
rect 152108 91156 152114 91158
rect 151721 91155 151787 91156
rect 153101 91155 153167 91158
rect 98494 91020 98500 91084
rect 98564 91082 98570 91084
rect 181621 91082 181687 91085
rect 98564 91080 181687 91082
rect 98564 91024 181626 91080
rect 181682 91024 181687 91080
rect 98564 91022 181687 91024
rect 98564 91020 98570 91022
rect 181621 91019 181687 91022
rect 209221 91082 209287 91085
rect 421281 91082 421347 91085
rect 209221 91080 421347 91082
rect 209221 91024 209226 91080
rect 209282 91024 421286 91080
rect 421342 91024 421347 91080
rect 209221 91022 421347 91024
rect 209221 91019 209287 91022
rect 421281 91019 421347 91022
rect 124438 90884 124444 90948
rect 124508 90946 124514 90948
rect 191281 90946 191347 90949
rect 124508 90944 191347 90946
rect 124508 90888 191286 90944
rect 191342 90888 191347 90944
rect 124508 90886 191347 90888
rect 124508 90884 124514 90886
rect 191281 90883 191347 90886
rect 115473 90402 115539 90405
rect 168373 90402 168439 90405
rect 115473 90400 168439 90402
rect 115473 90344 115478 90400
rect 115534 90344 168378 90400
rect 168434 90344 168439 90400
rect 115473 90342 168439 90344
rect 115473 90339 115539 90342
rect 168373 90339 168439 90342
rect 215937 90402 216003 90405
rect 249190 90402 249196 90404
rect 215937 90400 249196 90402
rect 215937 90344 215942 90400
rect 215998 90344 249196 90400
rect 215937 90342 249196 90344
rect 215937 90339 216003 90342
rect 249190 90340 249196 90342
rect 249260 90340 249266 90404
rect 352557 90402 352623 90405
rect 442022 90402 442028 90404
rect 352557 90400 442028 90402
rect 352557 90344 352562 90400
rect 352618 90344 442028 90400
rect 352557 90342 442028 90344
rect 352557 90339 352623 90342
rect 442022 90340 442028 90342
rect 442092 90340 442098 90404
rect 111333 89722 111399 89725
rect 194041 89722 194107 89725
rect 111333 89720 194107 89722
rect 111333 89664 111338 89720
rect 111394 89664 194046 89720
rect 194102 89664 194107 89720
rect 111333 89662 194107 89664
rect 111333 89659 111399 89662
rect 194041 89659 194107 89662
rect 215886 89660 215892 89724
rect 215956 89722 215962 89724
rect 410977 89722 411043 89725
rect 215956 89720 411043 89722
rect 215956 89664 410982 89720
rect 411038 89664 411043 89720
rect 215956 89662 411043 89664
rect 215956 89660 215962 89662
rect 410977 89659 411043 89662
rect 130745 89586 130811 89589
rect 167729 89586 167795 89589
rect 130745 89584 167795 89586
rect 130745 89528 130750 89584
rect 130806 89528 167734 89584
rect 167790 89528 167795 89584
rect 130745 89526 167795 89528
rect 130745 89523 130811 89526
rect 167729 89523 167795 89526
rect 162209 89042 162275 89045
rect 175917 89042 175983 89045
rect 162209 89040 175983 89042
rect 162209 88984 162214 89040
rect 162270 88984 175922 89040
rect 175978 88984 175983 89040
rect 162209 88982 175983 88984
rect 162209 88979 162275 88982
rect 175917 88979 175983 88982
rect 202229 89042 202295 89045
rect 230013 89042 230079 89045
rect 202229 89040 230079 89042
rect 202229 88984 202234 89040
rect 202290 88984 230018 89040
rect 230074 88984 230079 89040
rect 202229 88982 230079 88984
rect 202229 88979 202295 88982
rect 230013 88979 230079 88982
rect 304206 88980 304212 89044
rect 304276 89042 304282 89044
rect 326337 89042 326403 89045
rect 304276 89040 326403 89042
rect 304276 88984 326342 89040
rect 326398 88984 326403 89040
rect 304276 88982 326403 88984
rect 304276 88980 304282 88982
rect 326337 88979 326403 88982
rect 90725 88226 90791 88229
rect 178677 88226 178743 88229
rect 90725 88224 178743 88226
rect 90725 88168 90730 88224
rect 90786 88168 178682 88224
rect 178738 88168 178743 88224
rect 90725 88166 178743 88168
rect 90725 88163 90791 88166
rect 178677 88163 178743 88166
rect 217174 88164 217180 88228
rect 217244 88226 217250 88228
rect 282126 88226 282132 88228
rect 217244 88166 282132 88226
rect 217244 88164 217250 88166
rect 282126 88164 282132 88166
rect 282196 88164 282202 88228
rect 96337 88090 96403 88093
rect 167637 88090 167703 88093
rect 96337 88088 167703 88090
rect 96337 88032 96342 88088
rect 96398 88032 167642 88088
rect 167698 88032 167703 88088
rect 96337 88030 167703 88032
rect 96337 88027 96403 88030
rect 167637 88027 167703 88030
rect 112161 87954 112227 87957
rect 182909 87954 182975 87957
rect 112161 87952 182975 87954
rect 112161 87896 112166 87952
rect 112222 87896 182914 87952
rect 182970 87896 182975 87952
rect 112161 87894 182975 87896
rect 112161 87891 112227 87894
rect 182909 87891 182975 87894
rect 199469 87546 199535 87549
rect 228357 87546 228423 87549
rect 199469 87544 228423 87546
rect 199469 87488 199474 87544
rect 199530 87488 228362 87544
rect 228418 87488 228423 87544
rect 199469 87486 228423 87488
rect 199469 87483 199535 87486
rect 228357 87483 228423 87486
rect 91921 86866 91987 86869
rect 185761 86866 185827 86869
rect 91921 86864 185827 86866
rect 91921 86808 91926 86864
rect 91982 86808 185766 86864
rect 185822 86808 185827 86864
rect 91921 86806 185827 86808
rect 91921 86803 91987 86806
rect 185761 86803 185827 86806
rect 132861 86730 132927 86733
rect 178033 86730 178099 86733
rect 132861 86728 178099 86730
rect 132861 86672 132866 86728
rect 132922 86672 178038 86728
rect 178094 86672 178099 86728
rect 132861 86670 178099 86672
rect 132861 86667 132927 86670
rect 178033 86667 178099 86670
rect 206277 86322 206343 86325
rect 247033 86322 247099 86325
rect 299657 86324 299723 86325
rect 206277 86320 247099 86322
rect 206277 86264 206282 86320
rect 206338 86264 247038 86320
rect 247094 86264 247099 86320
rect 206277 86262 247099 86264
rect 206277 86259 206343 86262
rect 247033 86259 247099 86262
rect 299606 86260 299612 86324
rect 299676 86322 299723 86324
rect 299676 86320 299768 86322
rect 299718 86264 299768 86320
rect 299676 86262 299768 86264
rect 299676 86260 299723 86262
rect 299657 86259 299723 86260
rect 178677 86186 178743 86189
rect 257521 86186 257587 86189
rect 178677 86184 257587 86186
rect 178677 86128 178682 86184
rect 178738 86128 257526 86184
rect 257582 86128 257587 86184
rect 178677 86126 257587 86128
rect 178677 86123 178743 86126
rect 257521 86123 257587 86126
rect 582741 86186 582807 86189
rect 583520 86186 584960 86276
rect 582741 86184 584960 86186
rect 582741 86128 582746 86184
rect 582802 86128 584960 86184
rect 582741 86126 584960 86128
rect 582741 86123 582807 86126
rect 583520 86036 584960 86126
rect 104433 85506 104499 85509
rect 207749 85506 207815 85509
rect 104433 85504 207815 85506
rect 104433 85448 104438 85504
rect 104494 85448 207754 85504
rect 207810 85448 207815 85504
rect 104433 85446 207815 85448
rect 104433 85443 104499 85446
rect 207749 85443 207815 85446
rect 93025 85370 93091 85373
rect 166441 85370 166507 85373
rect 93025 85368 166507 85370
rect 93025 85312 93030 85368
rect 93086 85312 166446 85368
rect 166502 85312 166507 85368
rect 93025 85310 166507 85312
rect 93025 85307 93091 85310
rect 166441 85307 166507 85310
rect 118049 85234 118115 85237
rect 162485 85234 162551 85237
rect 118049 85232 162551 85234
rect 118049 85176 118054 85232
rect 118110 85176 162490 85232
rect 162546 85176 162551 85232
rect 118049 85174 162551 85176
rect 118049 85171 118115 85174
rect 162485 85171 162551 85174
rect 204989 84826 205055 84829
rect 309133 84826 309199 84829
rect 441613 84826 441679 84829
rect 204989 84824 441679 84826
rect -960 84690 480 84780
rect 204989 84768 204994 84824
rect 205050 84768 309138 84824
rect 309194 84768 441618 84824
rect 441674 84768 441679 84824
rect 204989 84766 441679 84768
rect 204989 84763 205055 84766
rect 309133 84763 309199 84766
rect 441613 84763 441679 84766
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 106917 84146 106983 84149
rect 181529 84146 181595 84149
rect 106917 84144 181595 84146
rect 106917 84088 106922 84144
rect 106978 84088 181534 84144
rect 181590 84088 181595 84144
rect 106917 84086 181595 84088
rect 106917 84083 106983 84086
rect 181529 84083 181595 84086
rect 219198 84084 219204 84148
rect 219268 84146 219274 84148
rect 279049 84146 279115 84149
rect 219268 84144 279115 84146
rect 219268 84088 279054 84144
rect 279110 84088 279115 84144
rect 219268 84086 279115 84088
rect 219268 84084 219274 84086
rect 279049 84083 279115 84086
rect 117221 83602 117287 83605
rect 267181 83602 267247 83605
rect 117221 83600 267247 83602
rect 117221 83544 117226 83600
rect 117282 83544 267186 83600
rect 267242 83544 267247 83600
rect 117221 83542 267247 83544
rect 117221 83539 117287 83542
rect 267181 83539 267247 83542
rect 34421 83466 34487 83469
rect 264094 83466 264100 83468
rect 34421 83464 264100 83466
rect 34421 83408 34426 83464
rect 34482 83408 264100 83464
rect 34421 83406 264100 83408
rect 34421 83403 34487 83406
rect 264094 83404 264100 83406
rect 264164 83404 264170 83468
rect 120717 82786 120783 82789
rect 210601 82786 210667 82789
rect 120717 82784 210667 82786
rect 120717 82728 120722 82784
rect 120778 82728 210606 82784
rect 210662 82728 210667 82784
rect 120717 82726 210667 82728
rect 120717 82723 120783 82726
rect 210601 82723 210667 82726
rect 105537 82650 105603 82653
rect 169293 82650 169359 82653
rect 105537 82648 169359 82650
rect 105537 82592 105542 82648
rect 105598 82592 169298 82648
rect 169354 82592 169359 82648
rect 105537 82590 169359 82592
rect 105537 82587 105603 82590
rect 169293 82587 169359 82590
rect 119981 82514 120047 82517
rect 162209 82514 162275 82517
rect 119981 82512 162275 82514
rect 119981 82456 119986 82512
rect 120042 82456 162214 82512
rect 162270 82456 162275 82512
rect 119981 82454 162275 82456
rect 119981 82451 120047 82454
rect 162209 82451 162275 82454
rect 197997 82242 198063 82245
rect 232681 82242 232747 82245
rect 197997 82240 232747 82242
rect 197997 82184 198002 82240
rect 198058 82184 232686 82240
rect 232742 82184 232747 82240
rect 197997 82182 232747 82184
rect 197997 82179 198063 82182
rect 232681 82179 232747 82182
rect 223021 82106 223087 82109
rect 278037 82106 278103 82109
rect 223021 82104 278103 82106
rect 223021 82048 223026 82104
rect 223082 82048 278042 82104
rect 278098 82048 278103 82104
rect 223021 82046 278103 82048
rect 223021 82043 223087 82046
rect 278037 82043 278103 82046
rect 95141 81426 95207 81429
rect 203701 81426 203767 81429
rect 95141 81424 203767 81426
rect 95141 81368 95146 81424
rect 95202 81368 203706 81424
rect 203762 81368 203767 81424
rect 95141 81366 203767 81368
rect 95141 81363 95207 81366
rect 203701 81363 203767 81366
rect 97257 81290 97323 81293
rect 170254 81290 170260 81292
rect 97257 81288 170260 81290
rect 97257 81232 97262 81288
rect 97318 81232 170260 81288
rect 97257 81230 170260 81232
rect 97257 81227 97323 81230
rect 170254 81228 170260 81230
rect 170324 81228 170330 81292
rect 12341 80746 12407 80749
rect 264513 80746 264579 80749
rect 12341 80744 264579 80746
rect 12341 80688 12346 80744
rect 12402 80688 264518 80744
rect 264574 80688 264579 80744
rect 12341 80686 264579 80688
rect 12341 80683 12407 80686
rect 264513 80683 264579 80686
rect 5441 79522 5507 79525
rect 228449 79522 228515 79525
rect 5441 79520 228515 79522
rect 5441 79464 5446 79520
rect 5502 79464 228454 79520
rect 228510 79464 228515 79520
rect 5441 79462 228515 79464
rect 5441 79459 5507 79462
rect 228449 79459 228515 79462
rect 26141 79386 26207 79389
rect 261661 79386 261727 79389
rect 26141 79384 261727 79386
rect 26141 79328 26146 79384
rect 26202 79328 261666 79384
rect 261722 79328 261727 79384
rect 26141 79326 261727 79328
rect 26141 79323 26207 79326
rect 261661 79323 261727 79326
rect 132401 78570 132467 78573
rect 166206 78570 166212 78572
rect 132401 78568 166212 78570
rect 132401 78512 132406 78568
rect 132462 78512 166212 78568
rect 132401 78510 166212 78512
rect 132401 78507 132467 78510
rect 166206 78508 166212 78510
rect 166276 78508 166282 78572
rect 95141 78026 95207 78029
rect 252093 78026 252159 78029
rect 95141 78024 252159 78026
rect 95141 77968 95146 78024
rect 95202 77968 252098 78024
rect 252154 77968 252159 78024
rect 95141 77966 252159 77968
rect 95141 77963 95207 77966
rect 252093 77963 252159 77966
rect 13721 77890 13787 77893
rect 266854 77890 266860 77892
rect 13721 77888 266860 77890
rect 13721 77832 13726 77888
rect 13782 77832 266860 77888
rect 13721 77830 266860 77832
rect 13721 77827 13787 77830
rect 266854 77828 266860 77830
rect 266924 77828 266930 77892
rect 280797 77890 280863 77893
rect 426382 77890 426388 77892
rect 280797 77888 426388 77890
rect 280797 77832 280802 77888
rect 280858 77832 426388 77888
rect 280797 77830 426388 77832
rect 280797 77827 280863 77830
rect 426382 77828 426388 77830
rect 426452 77828 426458 77892
rect 111701 76802 111767 76805
rect 256233 76802 256299 76805
rect 111701 76800 256299 76802
rect 111701 76744 111706 76800
rect 111762 76744 256238 76800
rect 256294 76744 256299 76800
rect 111701 76742 256299 76744
rect 111701 76739 111767 76742
rect 256233 76739 256299 76742
rect 70301 76666 70367 76669
rect 233969 76666 234035 76669
rect 70301 76664 234035 76666
rect 70301 76608 70306 76664
rect 70362 76608 233974 76664
rect 234030 76608 234035 76664
rect 70301 76606 234035 76608
rect 70301 76603 70367 76606
rect 233969 76603 234035 76606
rect 15101 76530 15167 76533
rect 262806 76530 262812 76532
rect 15101 76528 262812 76530
rect 15101 76472 15106 76528
rect 15162 76472 262812 76528
rect 15101 76470 262812 76472
rect 15101 76467 15167 76470
rect 262806 76468 262812 76470
rect 262876 76468 262882 76532
rect 97901 75306 97967 75309
rect 241053 75306 241119 75309
rect 97901 75304 241119 75306
rect 97901 75248 97906 75304
rect 97962 75248 241058 75304
rect 241114 75248 241119 75304
rect 97901 75246 241119 75248
rect 97901 75243 97967 75246
rect 241053 75243 241119 75246
rect 53741 75170 53807 75173
rect 249149 75170 249215 75173
rect 53741 75168 249215 75170
rect 53741 75112 53746 75168
rect 53802 75112 249154 75168
rect 249210 75112 249215 75168
rect 53741 75110 249215 75112
rect 53741 75107 53807 75110
rect 249149 75107 249215 75110
rect 111057 74490 111123 74493
rect 198181 74490 198247 74493
rect 111057 74488 198247 74490
rect 111057 74432 111062 74488
rect 111118 74432 198186 74488
rect 198242 74432 198247 74488
rect 111057 74430 198247 74432
rect 111057 74427 111123 74430
rect 198181 74427 198247 74430
rect 119981 73946 120047 73949
rect 257429 73946 257495 73949
rect 119981 73944 257495 73946
rect 119981 73888 119986 73944
rect 120042 73888 257434 73944
rect 257490 73888 257495 73944
rect 119981 73886 257495 73888
rect 119981 73883 120047 73886
rect 257429 73883 257495 73886
rect 73061 73810 73127 73813
rect 267273 73810 267339 73813
rect 73061 73808 267339 73810
rect 73061 73752 73066 73808
rect 73122 73752 267278 73808
rect 267334 73752 267339 73808
rect 73061 73750 267339 73752
rect 73061 73747 73127 73750
rect 267273 73747 267339 73750
rect 97809 73130 97875 73133
rect 166390 73130 166396 73132
rect 97809 73128 166396 73130
rect 97809 73072 97814 73128
rect 97870 73072 166396 73128
rect 97809 73070 166396 73072
rect 97809 73067 97875 73070
rect 166390 73068 166396 73070
rect 166460 73068 166466 73132
rect 582465 72994 582531 72997
rect 583520 72994 584960 73084
rect 582465 72992 584960 72994
rect 582465 72936 582470 72992
rect 582526 72936 584960 72992
rect 582465 72934 584960 72936
rect 582465 72931 582531 72934
rect 583520 72844 584960 72934
rect 30281 72450 30347 72453
rect 255957 72450 256023 72453
rect 30281 72448 256023 72450
rect 30281 72392 30286 72448
rect 30342 72392 255962 72448
rect 256018 72392 256023 72448
rect 30281 72390 256023 72392
rect 30281 72387 30347 72390
rect 255957 72387 256023 72390
rect 35157 71906 35223 71909
rect 35157 71904 35266 71906
rect 35157 71848 35162 71904
rect 35218 71848 35266 71904
rect 35157 71843 35266 71848
rect 35206 71770 35266 71843
rect 443085 71770 443151 71773
rect 6870 71768 443151 71770
rect -960 71634 480 71724
rect 6870 71712 443090 71768
rect 443146 71712 443151 71768
rect 6870 71710 443151 71712
rect 6870 71634 6930 71710
rect 443085 71707 443151 71710
rect -960 71574 6930 71634
rect -960 71484 480 71574
rect 68921 71090 68987 71093
rect 246389 71090 246455 71093
rect 68921 71088 246455 71090
rect 68921 71032 68926 71088
rect 68982 71032 246394 71088
rect 246450 71032 246455 71088
rect 68921 71030 246455 71032
rect 68921 71027 68987 71030
rect 246389 71027 246455 71030
rect 126881 69730 126947 69733
rect 191046 69730 191052 69732
rect 126881 69728 191052 69730
rect 126881 69672 126886 69728
rect 126942 69672 191052 69728
rect 126881 69670 191052 69672
rect 126881 69667 126947 69670
rect 191046 69668 191052 69670
rect 191116 69668 191122 69732
rect 75821 69594 75887 69597
rect 260189 69594 260255 69597
rect 75821 69592 260255 69594
rect 75821 69536 75826 69592
rect 75882 69536 260194 69592
rect 260250 69536 260255 69592
rect 75821 69534 260255 69536
rect 75821 69531 75887 69534
rect 260189 69531 260255 69534
rect 70209 68370 70275 68373
rect 245193 68370 245259 68373
rect 70209 68368 245259 68370
rect 70209 68312 70214 68368
rect 70270 68312 245198 68368
rect 245254 68312 245259 68368
rect 70209 68310 245259 68312
rect 70209 68307 70275 68310
rect 245193 68307 245259 68310
rect 53741 68234 53807 68237
rect 267089 68234 267155 68237
rect 53741 68232 267155 68234
rect 53741 68176 53746 68232
rect 53802 68176 267094 68232
rect 267150 68176 267155 68232
rect 53741 68174 267155 68176
rect 53741 68171 53807 68174
rect 267089 68171 267155 68174
rect 329097 68234 329163 68237
rect 430614 68234 430620 68236
rect 329097 68232 430620 68234
rect 329097 68176 329102 68232
rect 329158 68176 430620 68232
rect 329097 68174 430620 68176
rect 329097 68171 329163 68174
rect 430614 68172 430620 68174
rect 430684 68172 430690 68236
rect 77201 67010 77267 67013
rect 262949 67010 263015 67013
rect 77201 67008 263015 67010
rect 77201 66952 77206 67008
rect 77262 66952 262954 67008
rect 263010 66952 263015 67008
rect 77201 66950 263015 66952
rect 77201 66947 77267 66950
rect 262949 66947 263015 66950
rect 50889 66874 50955 66877
rect 256049 66874 256115 66877
rect 50889 66872 256115 66874
rect 50889 66816 50894 66872
rect 50950 66816 256054 66872
rect 256110 66816 256115 66872
rect 50889 66814 256115 66816
rect 50889 66811 50955 66814
rect 256049 66811 256115 66814
rect 273161 66874 273227 66877
rect 298134 66874 298140 66876
rect 273161 66872 298140 66874
rect 273161 66816 273166 66872
rect 273222 66816 298140 66872
rect 273161 66814 298140 66816
rect 273161 66811 273227 66814
rect 298134 66812 298140 66814
rect 298204 66812 298210 66876
rect 291142 66132 291148 66196
rect 291212 66194 291218 66196
rect 292481 66194 292547 66197
rect 291212 66192 292547 66194
rect 291212 66136 292486 66192
rect 292542 66136 292547 66192
rect 291212 66134 292547 66136
rect 291212 66132 291218 66134
rect 292481 66131 292547 66134
rect 79961 65650 80027 65653
rect 258901 65650 258967 65653
rect 79961 65648 258967 65650
rect 79961 65592 79966 65648
rect 80022 65592 258906 65648
rect 258962 65592 258967 65648
rect 79961 65590 258967 65592
rect 79961 65587 80027 65590
rect 258901 65587 258967 65590
rect 38561 65514 38627 65517
rect 253289 65514 253355 65517
rect 38561 65512 253355 65514
rect 38561 65456 38566 65512
rect 38622 65456 253294 65512
rect 253350 65456 253355 65512
rect 38561 65454 253355 65456
rect 38561 65451 38627 65454
rect 253289 65451 253355 65454
rect 147029 64290 147095 64293
rect 181437 64290 181503 64293
rect 147029 64288 181503 64290
rect 147029 64232 147034 64288
rect 147090 64232 181442 64288
rect 181498 64232 181503 64288
rect 147029 64230 181503 64232
rect 147029 64227 147095 64230
rect 181437 64227 181503 64230
rect 186814 64228 186820 64292
rect 186884 64290 186890 64292
rect 283557 64290 283623 64293
rect 186884 64288 283623 64290
rect 186884 64232 283562 64288
rect 283618 64232 283623 64288
rect 186884 64230 283623 64232
rect 186884 64228 186890 64230
rect 283557 64227 283623 64230
rect 23381 64154 23447 64157
rect 245101 64154 245167 64157
rect 23381 64152 245167 64154
rect 23381 64096 23386 64152
rect 23442 64096 245106 64152
rect 245162 64096 245167 64152
rect 23381 64094 245167 64096
rect 23381 64091 23447 64094
rect 245101 64091 245167 64094
rect 102041 62930 102107 62933
rect 250621 62930 250687 62933
rect 102041 62928 250687 62930
rect 102041 62872 102046 62928
rect 102102 62872 250626 62928
rect 250682 62872 250687 62928
rect 102041 62870 250687 62872
rect 102041 62867 102107 62870
rect 250621 62867 250687 62870
rect 19241 62794 19307 62797
rect 267774 62794 267780 62796
rect 19241 62792 267780 62794
rect 19241 62736 19246 62792
rect 19302 62736 267780 62792
rect 19241 62734 267780 62736
rect 19241 62731 19307 62734
rect 267774 62732 267780 62734
rect 267844 62732 267850 62796
rect 87597 61434 87663 61437
rect 265617 61434 265683 61437
rect 87597 61432 265683 61434
rect 87597 61376 87602 61432
rect 87658 61376 265622 61432
rect 265678 61376 265683 61432
rect 87597 61374 265683 61376
rect 87597 61371 87663 61374
rect 265617 61371 265683 61374
rect 310513 60618 310579 60621
rect 311157 60618 311223 60621
rect 424174 60618 424180 60620
rect 310513 60616 424180 60618
rect 310513 60560 310518 60616
rect 310574 60560 311162 60616
rect 311218 60560 424180 60616
rect 310513 60558 424180 60560
rect 310513 60555 310579 60558
rect 311157 60555 311223 60558
rect 424174 60556 424180 60558
rect 424244 60556 424250 60620
rect 57789 59938 57855 59941
rect 252001 59938 252067 59941
rect 57789 59936 252067 59938
rect 57789 59880 57794 59936
rect 57850 59880 252006 59936
rect 252062 59880 252067 59936
rect 57789 59878 252067 59880
rect 57789 59875 57855 59878
rect 252001 59875 252067 59878
rect 582649 59666 582715 59669
rect 583520 59666 584960 59756
rect 582649 59664 584960 59666
rect 582649 59608 582654 59664
rect 582710 59608 584960 59664
rect 582649 59606 584960 59608
rect 582649 59603 582715 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 31661 58578 31727 58581
rect 250529 58578 250595 58581
rect 31661 58576 250595 58578
rect 31661 58520 31666 58576
rect 31722 58520 250534 58576
rect 250590 58520 250595 58576
rect 31661 58518 250595 58520
rect 31661 58515 31727 58518
rect 250529 58515 250595 58518
rect 35801 57218 35867 57221
rect 229829 57218 229895 57221
rect 35801 57216 229895 57218
rect 35801 57160 35806 57216
rect 35862 57160 229834 57216
rect 229890 57160 229895 57216
rect 35801 57158 229895 57160
rect 35801 57155 35867 57158
rect 229829 57155 229895 57158
rect 10961 55858 11027 55861
rect 254577 55858 254643 55861
rect 10961 55856 254643 55858
rect 10961 55800 10966 55856
rect 11022 55800 254582 55856
rect 254638 55800 254643 55856
rect 10961 55798 254643 55800
rect 10961 55795 11027 55798
rect 254577 55795 254643 55798
rect 282177 55858 282243 55861
rect 436686 55858 436692 55860
rect 282177 55856 436692 55858
rect 282177 55800 282182 55856
rect 282238 55800 436692 55856
rect 282177 55798 436692 55800
rect 282177 55795 282243 55798
rect 436686 55796 436692 55798
rect 436756 55796 436762 55860
rect 48221 54498 48287 54501
rect 308397 54498 308463 54501
rect 48221 54496 308463 54498
rect 48221 54440 48226 54496
rect 48282 54440 308402 54496
rect 308458 54440 308463 54496
rect 48221 54438 308463 54440
rect 48221 54435 48287 54438
rect 308397 54435 308463 54438
rect 22001 53138 22067 53141
rect 260230 53138 260236 53140
rect 22001 53136 260236 53138
rect 22001 53080 22006 53136
rect 22062 53080 260236 53136
rect 22001 53078 260236 53080
rect 22001 53075 22067 53078
rect 260230 53076 260236 53078
rect 260300 53076 260306 53140
rect 93761 51778 93827 51781
rect 233734 51778 233740 51780
rect 93761 51776 233740 51778
rect 93761 51720 93766 51776
rect 93822 51720 233740 51776
rect 93761 51718 233740 51720
rect 93761 51715 93827 51718
rect 233734 51716 233740 51718
rect 233804 51716 233810 51780
rect 53649 50282 53715 50285
rect 243629 50282 243695 50285
rect 53649 50280 243695 50282
rect 53649 50224 53654 50280
rect 53710 50224 243634 50280
rect 243690 50224 243695 50280
rect 53649 50222 243695 50224
rect 53649 50219 53715 50222
rect 243629 50219 243695 50222
rect 66161 48922 66227 48925
rect 256141 48922 256207 48925
rect 66161 48920 256207 48922
rect 66161 48864 66166 48920
rect 66222 48864 256146 48920
rect 256202 48864 256207 48920
rect 66161 48862 256207 48864
rect 66161 48859 66227 48862
rect 256141 48859 256207 48862
rect 33041 47562 33107 47565
rect 251909 47562 251975 47565
rect 33041 47560 251975 47562
rect 33041 47504 33046 47560
rect 33102 47504 251914 47560
rect 251970 47504 251975 47560
rect 33041 47502 251975 47504
rect 33041 47499 33107 47502
rect 251909 47499 251975 47502
rect 583017 46338 583083 46341
rect 583520 46338 584960 46428
rect 583017 46336 584960 46338
rect 583017 46280 583022 46336
rect 583078 46280 584960 46336
rect 583017 46278 584960 46280
rect 583017 46275 583083 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 64781 44842 64847 44845
rect 258574 44842 258580 44844
rect 64781 44840 258580 44842
rect 64781 44784 64786 44840
rect 64842 44784 258580 44840
rect 64781 44782 258580 44784
rect 64781 44779 64847 44782
rect 258574 44780 258580 44782
rect 258644 44780 258650 44844
rect 44081 43482 44147 43485
rect 249006 43482 249012 43484
rect 44081 43480 249012 43482
rect 44081 43424 44086 43480
rect 44142 43424 249012 43480
rect 44081 43422 249012 43424
rect 44081 43419 44147 43422
rect 249006 43420 249012 43422
rect 249076 43420 249082 43484
rect 144821 40626 144887 40629
rect 388437 40626 388503 40629
rect 144821 40624 388503 40626
rect 144821 40568 144826 40624
rect 144882 40568 388442 40624
rect 388498 40568 388503 40624
rect 144821 40566 388503 40568
rect 144821 40563 144887 40566
rect 388437 40563 388503 40566
rect 49601 39402 49667 39405
rect 246246 39402 246252 39404
rect 49601 39400 246252 39402
rect 49601 39344 49606 39400
rect 49662 39344 246252 39400
rect 49601 39342 246252 39344
rect 49601 39339 49667 39342
rect 246246 39340 246252 39342
rect 246316 39340 246322 39404
rect 6821 39266 6887 39269
rect 224902 39266 224908 39268
rect 6821 39264 224908 39266
rect 6821 39208 6826 39264
rect 6882 39208 224908 39264
rect 6821 39206 224908 39208
rect 6821 39203 6887 39206
rect 224902 39204 224908 39206
rect 224972 39204 224978 39268
rect 169518 37980 169524 38044
rect 169588 38042 169594 38044
rect 273897 38042 273963 38045
rect 169588 38040 273963 38042
rect 169588 37984 273902 38040
rect 273958 37984 273963 38040
rect 169588 37982 273963 37984
rect 169588 37980 169594 37982
rect 273897 37979 273963 37982
rect 65926 37844 65932 37908
rect 65996 37906 66002 37908
rect 325049 37906 325115 37909
rect 65996 37904 325115 37906
rect 65996 37848 325054 37904
rect 325110 37848 325115 37904
rect 65996 37846 325115 37848
rect 65996 37844 66002 37846
rect 325049 37843 325115 37846
rect 4061 36546 4127 36549
rect 242014 36546 242020 36548
rect 4061 36544 242020 36546
rect 4061 36488 4066 36544
rect 4122 36488 242020 36544
rect 4061 36486 242020 36488
rect 4061 36483 4127 36486
rect 242014 36484 242020 36486
rect 242084 36484 242090 36548
rect 28901 35186 28967 35189
rect 273345 35186 273411 35189
rect 28901 35184 273411 35186
rect 28901 35128 28906 35184
rect 28962 35128 273350 35184
rect 273406 35128 273411 35184
rect 28901 35126 273411 35128
rect 28901 35123 28967 35126
rect 273345 35123 273411 35126
rect 313917 34506 313983 34509
rect 314561 34506 314627 34509
rect 439078 34506 439084 34508
rect 313917 34504 439084 34506
rect 313917 34448 313922 34504
rect 313978 34448 314566 34504
rect 314622 34448 439084 34504
rect 313917 34446 439084 34448
rect 313917 34443 313983 34446
rect 314561 34443 314627 34446
rect 439078 34444 439084 34446
rect 439148 34444 439154 34508
rect 582833 33146 582899 33149
rect 583520 33146 584960 33236
rect 582833 33144 584960 33146
rect 582833 33088 582838 33144
rect 582894 33088 584960 33144
rect 582833 33086 584960 33088
rect 582833 33083 582899 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 302969 30970 303035 30973
rect 434846 30970 434852 30972
rect 302969 30968 434852 30970
rect 302969 30912 302974 30968
rect 303030 30912 434852 30968
rect 302969 30910 434852 30912
rect 302969 30907 303035 30910
rect 434846 30908 434852 30910
rect 434916 30908 434922 30972
rect 202137 30290 202203 30293
rect 252553 30290 252619 30293
rect 202137 30288 252619 30290
rect 202137 30232 202142 30288
rect 202198 30232 252558 30288
rect 252614 30232 252619 30288
rect 202137 30230 252619 30232
rect 202137 30227 202203 30230
rect 252553 30227 252619 30230
rect 269113 29610 269179 29613
rect 281574 29610 281580 29612
rect 269113 29608 281580 29610
rect 269113 29552 269118 29608
rect 269174 29552 281580 29608
rect 269113 29550 281580 29552
rect 269113 29547 269179 29550
rect 281574 29548 281580 29550
rect 281644 29548 281650 29612
rect 141417 28250 141483 28253
rect 189717 28250 189783 28253
rect 141417 28248 189783 28250
rect 141417 28192 141422 28248
rect 141478 28192 189722 28248
rect 189778 28192 189783 28248
rect 141417 28190 189783 28192
rect 141417 28187 141483 28190
rect 189717 28187 189783 28190
rect 184289 26890 184355 26893
rect 280889 26890 280955 26893
rect 184289 26888 280955 26890
rect 184289 26832 184294 26888
rect 184350 26832 280894 26888
rect 280950 26832 280955 26888
rect 184289 26830 280955 26832
rect 184289 26827 184355 26830
rect 280889 26827 280955 26830
rect 52269 26210 52335 26213
rect 324405 26210 324471 26213
rect 324957 26210 325023 26213
rect 52269 26208 325023 26210
rect 52269 26152 52274 26208
rect 52330 26152 324410 26208
rect 324466 26152 324962 26208
rect 325018 26152 325023 26208
rect 52269 26150 325023 26152
rect 52269 26147 52335 26150
rect 324405 26147 324471 26150
rect 324957 26147 325023 26150
rect 67766 24788 67772 24852
rect 67836 24850 67842 24852
rect 284937 24850 285003 24853
rect 67836 24848 285003 24850
rect 67836 24792 284942 24848
rect 284998 24792 285003 24848
rect 67836 24790 285003 24792
rect 67836 24788 67842 24790
rect 284937 24787 285003 24790
rect 284293 23490 284359 23493
rect 284937 23490 285003 23493
rect 284293 23488 285003 23490
rect 284293 23432 284298 23488
rect 284354 23432 284942 23488
rect 284998 23432 285003 23488
rect 284293 23430 285003 23432
rect 284293 23427 284359 23430
rect 284937 23427 285003 23430
rect 287646 21388 287652 21452
rect 287716 21450 287722 21452
rect 288750 21450 288756 21452
rect 287716 21390 288756 21450
rect 287716 21388 287722 21390
rect 288750 21388 288756 21390
rect 288820 21388 288826 21452
rect 130377 19954 130443 19957
rect 172462 19954 172468 19956
rect 130377 19952 172468 19954
rect 130377 19896 130382 19952
rect 130438 19896 172468 19952
rect 130377 19894 172468 19896
rect 130377 19891 130443 19894
rect 172462 19892 172468 19894
rect 172532 19892 172538 19956
rect 582557 19818 582623 19821
rect 583520 19818 584960 19908
rect 582557 19816 584960 19818
rect 582557 19760 582562 19816
rect 582618 19760 584960 19816
rect 582557 19758 584960 19760
rect 582557 19755 582623 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 253054 19348 253060 19412
rect 253124 19410 253130 19412
rect 259545 19410 259611 19413
rect 260097 19410 260163 19413
rect 253124 19408 260163 19410
rect 253124 19352 259550 19408
rect 259606 19352 260102 19408
rect 260158 19352 260163 19408
rect 253124 19350 260163 19352
rect 253124 19348 253130 19350
rect 259545 19347 259611 19350
rect 260097 19347 260163 19350
rect 55070 19212 55076 19276
rect 55140 19274 55146 19276
rect 262213 19274 262279 19277
rect 262949 19274 263015 19277
rect 55140 19272 263015 19274
rect 55140 19216 262218 19272
rect 262274 19216 262954 19272
rect 263010 19216 263015 19272
rect 55140 19214 263015 19216
rect 55140 19212 55146 19214
rect 262213 19211 262279 19214
rect 262949 19211 263015 19214
rect 59118 15132 59124 15196
rect 59188 15194 59194 15196
rect 249977 15194 250043 15197
rect 59188 15192 250043 15194
rect 59188 15136 249982 15192
rect 250038 15136 250043 15192
rect 59188 15134 250043 15136
rect 59188 15132 59194 15134
rect 249977 15131 250043 15134
rect 316677 14514 316743 14517
rect 425462 14514 425468 14516
rect 316677 14512 425468 14514
rect 316677 14456 316682 14512
rect 316738 14456 425468 14512
rect 316677 14454 425468 14456
rect 316677 14451 316743 14454
rect 425462 14452 425468 14454
rect 425532 14452 425538 14516
rect 273897 12338 273963 12341
rect 274541 12338 274607 12341
rect 376109 12338 376175 12341
rect 273897 12336 376175 12338
rect 273897 12280 273902 12336
rect 273958 12280 274546 12336
rect 274602 12280 376114 12336
rect 376170 12280 376175 12336
rect 273897 12278 376175 12280
rect 273897 12275 273963 12278
rect 274541 12275 274607 12278
rect 376109 12275 376175 12278
rect 288341 12202 288407 12205
rect 288750 12202 288756 12204
rect 288341 12200 288756 12202
rect 288341 12144 288346 12200
rect 288402 12144 288756 12200
rect 288341 12142 288756 12144
rect 288341 12139 288407 12142
rect 288750 12140 288756 12142
rect 288820 12140 288826 12204
rect 299606 11732 299612 11796
rect 299676 11794 299682 11796
rect 300761 11794 300827 11797
rect 299676 11792 300827 11794
rect 299676 11736 300766 11792
rect 300822 11736 300827 11792
rect 299676 11734 300827 11736
rect 299676 11732 299682 11734
rect 300761 11731 300827 11734
rect 42701 11658 42767 11661
rect 230974 11658 230980 11660
rect 42701 11656 230980 11658
rect 42701 11600 42706 11656
rect 42762 11600 230980 11656
rect 42701 11598 230980 11600
rect 42701 11595 42767 11598
rect 230974 11596 230980 11598
rect 231044 11596 231050 11660
rect 175181 10298 175247 10301
rect 261753 10298 261819 10301
rect 175181 10296 261819 10298
rect 175181 10240 175186 10296
rect 175242 10240 261758 10296
rect 261814 10240 261819 10296
rect 175181 10238 261819 10240
rect 175181 10235 175247 10238
rect 261753 10235 261819 10238
rect 377397 9618 377463 9621
rect 258030 9616 377463 9618
rect 258030 9560 377402 9616
rect 377458 9560 377463 9616
rect 258030 9558 377463 9560
rect 251909 9482 251975 9485
rect 258030 9482 258090 9558
rect 377397 9555 377463 9558
rect 251909 9480 258090 9482
rect 251909 9424 251914 9480
rect 251970 9424 258090 9480
rect 251909 9422 258090 9424
rect 251909 9419 251975 9422
rect 288566 8196 288572 8260
rect 288636 8258 288642 8260
rect 288985 8258 289051 8261
rect 288636 8256 289051 8258
rect 288636 8200 288990 8256
rect 289046 8200 289051 8256
rect 288636 8198 289051 8200
rect 288636 8196 288642 8198
rect 288985 8195 289051 8198
rect 184197 7578 184263 7581
rect 292573 7578 292639 7581
rect 184197 7576 292639 7578
rect 184197 7520 184202 7576
rect 184258 7520 292578 7576
rect 292634 7520 292639 7576
rect 184197 7518 292639 7520
rect 184197 7515 184263 7518
rect 292573 7515 292639 7518
rect 300669 7578 300735 7581
rect 420862 7578 420868 7580
rect 300669 7576 420868 7578
rect 300669 7520 300674 7576
rect 300730 7520 420868 7576
rect 300669 7518 420868 7520
rect 300669 7515 300735 7518
rect 420862 7516 420868 7518
rect 420932 7516 420938 7580
rect 182817 6898 182883 6901
rect 268377 6898 268443 6901
rect 182817 6896 268443 6898
rect 182817 6840 182822 6896
rect 182878 6840 268382 6896
rect 268438 6840 268443 6896
rect 182817 6838 268443 6840
rect 182817 6835 182883 6838
rect 268377 6835 268443 6838
rect 13 6762 79 6765
rect 13 6760 122 6762
rect 13 6704 18 6760
rect 74 6704 122 6760
rect 13 6699 122 6704
rect 62 6626 122 6699
rect 583109 6626 583175 6629
rect 583520 6626 584960 6716
rect 62 6580 674 6626
rect -960 6566 674 6580
rect -960 6490 480 6566
rect 614 6490 674 6566
rect 583109 6624 584960 6626
rect 583109 6568 583114 6624
rect 583170 6568 584960 6624
rect 583109 6566 584960 6568
rect 583109 6563 583175 6566
rect -960 6430 674 6490
rect 583520 6476 584960 6566
rect -960 6340 480 6430
rect 132953 6218 133019 6221
rect 166993 6218 167059 6221
rect 132953 6216 167059 6218
rect 132953 6160 132958 6216
rect 133014 6160 166998 6216
rect 167054 6160 167059 6216
rect 132953 6158 167059 6160
rect 132953 6155 133019 6158
rect 166993 6155 167059 6158
rect 188838 4932 188844 4996
rect 188908 4994 188914 4996
rect 244089 4994 244155 4997
rect 188908 4992 244155 4994
rect 188908 4936 244094 4992
rect 244150 4936 244155 4992
rect 188908 4934 244155 4936
rect 188908 4932 188914 4934
rect 244089 4931 244155 4934
rect 1669 4858 1735 4861
rect 227662 4858 227668 4860
rect 1669 4856 227668 4858
rect 1669 4800 1674 4856
rect 1730 4800 227668 4856
rect 1669 4798 227668 4800
rect 1669 4795 1735 4798
rect 227662 4796 227668 4798
rect 227732 4796 227738 4860
rect 177297 4042 177363 4045
rect 282269 4042 282335 4045
rect 177297 4040 282335 4042
rect 177297 3984 177302 4040
rect 177358 3984 282274 4040
rect 282330 3984 282335 4040
rect 177297 3982 282335 3984
rect 177297 3979 177363 3982
rect 282269 3979 282335 3982
rect 298686 3980 298692 4044
rect 298756 4042 298762 4044
rect 299657 4042 299723 4045
rect 300669 4042 300735 4045
rect 298756 4040 300735 4042
rect 298756 3984 299662 4040
rect 299718 3984 300674 4040
rect 300730 3984 300735 4040
rect 298756 3982 300735 3984
rect 298756 3980 298762 3982
rect 299657 3979 299723 3982
rect 300669 3979 300735 3982
rect 308397 4042 308463 4045
rect 309041 4042 309107 4045
rect 382917 4042 382983 4045
rect 308397 4040 309107 4042
rect 308397 3984 308402 4040
rect 308458 3984 309046 4040
rect 309102 3984 309107 4040
rect 308397 3982 309107 3984
rect 308397 3979 308463 3982
rect 309041 3979 309107 3982
rect 354630 4040 382983 4042
rect 354630 3984 382922 4040
rect 382978 3984 382983 4040
rect 354630 3982 382983 3984
rect 240726 3844 240732 3908
rect 240796 3906 240802 3908
rect 245653 3906 245719 3909
rect 280797 3906 280863 3909
rect 240796 3904 245719 3906
rect 240796 3848 245658 3904
rect 245714 3848 245719 3904
rect 240796 3846 245719 3848
rect 240796 3844 240802 3846
rect 245653 3843 245719 3846
rect 258030 3904 280863 3906
rect 258030 3848 280802 3904
rect 280858 3848 280863 3904
rect 258030 3846 280863 3848
rect 251817 3634 251883 3637
rect 252369 3634 252435 3637
rect 258030 3634 258090 3846
rect 280797 3843 280863 3846
rect 351637 3906 351703 3909
rect 354630 3906 354690 3982
rect 382917 3979 382983 3982
rect 351637 3904 354690 3906
rect 351637 3848 351642 3904
rect 351698 3848 354690 3904
rect 351637 3846 354690 3848
rect 351637 3843 351703 3846
rect 292573 3770 292639 3773
rect 322289 3770 322355 3773
rect 292573 3768 322355 3770
rect 292573 3712 292578 3768
rect 292634 3712 322294 3768
rect 322350 3712 322355 3768
rect 292573 3710 322355 3712
rect 292573 3707 292639 3710
rect 322289 3707 322355 3710
rect 251817 3632 258090 3634
rect 251817 3576 251822 3632
rect 251878 3576 252374 3632
rect 252430 3576 258090 3632
rect 251817 3574 258090 3576
rect 251817 3571 251883 3574
rect 252369 3571 252435 3574
rect 121085 3498 121151 3501
rect 170397 3498 170463 3501
rect 121085 3496 170463 3498
rect 121085 3440 121090 3496
rect 121146 3440 170402 3496
rect 170458 3440 170463 3496
rect 121085 3438 170463 3440
rect 121085 3435 121151 3438
rect 170397 3435 170463 3438
rect 260097 3498 260163 3501
rect 260649 3498 260715 3501
rect 260097 3496 260715 3498
rect 260097 3440 260102 3496
rect 260158 3440 260654 3496
rect 260710 3440 260715 3496
rect 260097 3438 260715 3440
rect 260097 3435 260163 3438
rect 260649 3435 260715 3438
rect 268326 3436 268332 3500
rect 268396 3498 268402 3500
rect 276105 3498 276171 3501
rect 268396 3496 276171 3498
rect 268396 3440 276110 3496
rect 276166 3440 276171 3496
rect 268396 3438 276171 3440
rect 268396 3436 268402 3438
rect 276105 3435 276171 3438
rect 287789 3498 287855 3501
rect 288341 3498 288407 3501
rect 287789 3496 288407 3498
rect 287789 3440 287794 3496
rect 287850 3440 288346 3496
rect 288402 3440 288407 3496
rect 287789 3438 288407 3440
rect 287789 3435 287855 3438
rect 288341 3435 288407 3438
rect 350441 3498 350507 3501
rect 352557 3498 352623 3501
rect 350441 3496 352623 3498
rect 350441 3440 350446 3496
rect 350502 3440 352562 3496
rect 352618 3440 352623 3496
rect 350441 3438 352623 3440
rect 350441 3435 350507 3438
rect 352557 3435 352623 3438
rect 85665 3362 85731 3365
rect 189717 3362 189783 3365
rect 85665 3360 189783 3362
rect 85665 3304 85670 3360
rect 85726 3304 189722 3360
rect 189778 3304 189783 3360
rect 85665 3302 189783 3304
rect 85665 3299 85731 3302
rect 189717 3299 189783 3302
rect 209037 3362 209103 3365
rect 247585 3362 247651 3365
rect 247769 3362 247835 3365
rect 209037 3360 247835 3362
rect 209037 3304 209042 3360
rect 209098 3304 247590 3360
rect 247646 3304 247774 3360
rect 247830 3304 247835 3360
rect 209037 3302 247835 3304
rect 209037 3299 209103 3302
rect 247585 3299 247651 3302
rect 247769 3299 247835 3302
rect 342161 3362 342227 3365
rect 358077 3362 358143 3365
rect 342161 3360 358143 3362
rect 342161 3304 342166 3360
rect 342222 3304 358082 3360
rect 358138 3304 358143 3360
rect 342161 3302 358143 3304
rect 342161 3299 342227 3302
rect 358077 3299 358143 3302
rect 82077 2002 82143 2005
rect 177389 2002 177455 2005
rect 82077 2000 177455 2002
rect 82077 1944 82082 2000
rect 82138 1944 177394 2000
rect 177450 1944 177455 2000
rect 82077 1942 177455 1944
rect 82077 1939 82143 1942
rect 177389 1939 177455 1942
<< via3 >>
rect 69612 702476 69676 702540
rect 88196 588508 88260 588572
rect 88196 585652 88260 585716
rect 69428 582252 69492 582316
rect 119476 579668 119540 579732
rect 67772 578852 67836 578916
rect 120028 578308 120092 578372
rect 166212 557500 166276 557564
rect 66668 556820 66732 556884
rect 115060 553420 115124 553484
rect 160692 547844 160756 547908
rect 353340 546620 353404 546684
rect 91508 546484 91572 546548
rect 191052 545260 191116 545324
rect 200804 545124 200868 545188
rect 352052 544036 352116 544100
rect 181300 543900 181364 543964
rect 68692 542948 68756 543012
rect 161244 542404 161308 542468
rect 356100 542464 356164 542468
rect 356100 542408 356114 542464
rect 356114 542408 356164 542464
rect 356100 542404 356164 542408
rect 88196 541452 88260 541516
rect 91508 541180 91572 541244
rect 197860 541180 197924 541244
rect 352236 541180 352300 541244
rect 159220 539684 159284 539748
rect 99972 538868 100036 538932
rect 106412 538732 106476 538796
rect 195100 538460 195164 538524
rect 88196 536692 88260 536756
rect 69612 535528 69676 535532
rect 69612 535472 69626 535528
rect 69626 535472 69676 535528
rect 69612 535468 69676 535472
rect 199332 535468 199396 535532
rect 67772 535332 67836 535396
rect 199884 535196 199948 535260
rect 199332 527716 199396 527780
rect 175780 526356 175844 526420
rect 197860 526356 197924 526420
rect 163452 518876 163516 518940
rect 161980 514796 162044 514860
rect 360148 514932 360212 514996
rect 198596 512484 198660 512548
rect 356284 499836 356348 499900
rect 168972 496844 169036 496908
rect 356284 480116 356348 480180
rect 104940 471140 105004 471204
rect 89668 469780 89732 469844
rect 118004 469780 118068 469844
rect 100708 468420 100772 468484
rect 115980 468420 116044 468484
rect 108988 467060 109052 467124
rect 96660 465700 96724 465764
rect 107700 465700 107764 465764
rect 156644 465216 156708 465220
rect 156644 465160 156658 465216
rect 156658 465160 156708 465216
rect 156644 465156 156708 465160
rect 102180 462844 102244 462908
rect 91140 458900 91204 458964
rect 198780 458356 198844 458420
rect 98132 457540 98196 457604
rect 111748 457404 111812 457468
rect 72004 456044 72068 456108
rect 92612 456044 92676 456108
rect 69060 452508 69124 452572
rect 69060 451828 69124 451892
rect 184796 449924 184860 449988
rect 93900 449108 93964 449172
rect 122604 449108 122668 449172
rect 95188 447748 95252 447812
rect 187004 447068 187068 447132
rect 71820 446388 71884 446452
rect 72004 445844 72068 445908
rect 72740 445844 72804 445908
rect 93716 445844 93780 445908
rect 100524 445768 100588 445772
rect 100524 445712 100538 445768
rect 100538 445712 100588 445768
rect 100524 445708 100588 445712
rect 114324 445768 114388 445772
rect 114324 445712 114374 445768
rect 114374 445712 114388 445768
rect 114324 445708 114388 445712
rect 118556 445768 118620 445772
rect 118556 445712 118570 445768
rect 118570 445712 118620 445768
rect 118556 445708 118620 445712
rect 94452 444816 94516 444820
rect 94452 444760 94502 444816
rect 94502 444760 94516 444816
rect 94452 444756 94516 444760
rect 109540 444892 109604 444956
rect 111564 444892 111628 444956
rect 154068 442308 154132 442372
rect 196572 438908 196636 438972
rect 357572 438908 357636 438972
rect 120212 430578 120276 430642
rect 177804 430612 177868 430676
rect 120396 428708 120460 428772
rect 121684 426260 121748 426324
rect 122604 426260 122668 426324
rect 66668 419596 66732 419660
rect 67772 419596 67836 419660
rect 121500 419596 121564 419660
rect 69060 409940 69124 410004
rect 358860 409396 358924 409460
rect 173020 401644 173084 401708
rect 173204 396068 173268 396132
rect 360332 396884 360396 396948
rect 122788 394708 122852 394772
rect 65932 393212 65996 393276
rect 119476 392124 119540 392188
rect 80468 391308 80532 391372
rect 104940 391036 105004 391100
rect 80468 390900 80532 390964
rect 121500 390628 121564 390692
rect 71820 390552 71884 390556
rect 71820 390496 71870 390552
rect 71870 390496 71884 390552
rect 71820 390492 71884 390496
rect 108988 390492 109052 390556
rect 69612 390356 69676 390420
rect 89668 390356 89732 390420
rect 91140 390356 91204 390420
rect 92612 390356 92676 390420
rect 93900 390356 93964 390420
rect 95372 390356 95436 390420
rect 96660 390356 96724 390420
rect 98132 390356 98196 390420
rect 100708 390416 100772 390420
rect 100708 390360 100722 390416
rect 100722 390360 100772 390416
rect 100708 390356 100772 390360
rect 102180 390416 102244 390420
rect 102180 390360 102194 390416
rect 102194 390360 102244 390416
rect 102180 390356 102244 390360
rect 106412 390356 106476 390420
rect 107700 390356 107764 390420
rect 115980 390416 116044 390420
rect 115980 390360 115994 390416
rect 115994 390360 116044 390416
rect 115980 390356 116044 390360
rect 118004 390356 118068 390420
rect 76420 390220 76484 390284
rect 89668 389132 89732 389196
rect 111748 388996 111812 389060
rect 99972 388860 100036 388924
rect 115060 388860 115124 388924
rect 83964 388784 84028 388788
rect 83964 388728 83978 388784
rect 83978 388728 84028 388784
rect 83964 388724 84028 388728
rect 95188 387772 95252 387836
rect 100524 387832 100588 387836
rect 100524 387776 100538 387832
rect 100538 387776 100588 387832
rect 100524 387772 100588 387776
rect 192340 386412 192404 386476
rect 95188 385596 95252 385660
rect 198596 385052 198660 385116
rect 120212 384236 120276 384300
rect 122604 382876 122668 382940
rect 356100 382604 356164 382668
rect 356468 382604 356532 382668
rect 356100 381924 356164 381988
rect 194548 381516 194612 381580
rect 67772 378660 67836 378724
rect 359412 378116 359476 378180
rect 179276 377300 179340 377364
rect 359412 376892 359476 376956
rect 199884 376484 199948 376548
rect 352236 376484 352300 376548
rect 354628 375728 354692 375732
rect 354628 375672 354678 375728
rect 354678 375672 354692 375728
rect 354628 375668 354692 375672
rect 194548 375260 194612 375324
rect 288756 375260 288820 375324
rect 356468 374036 356532 374100
rect 357572 373220 357636 373284
rect 180564 371860 180628 371924
rect 358860 371316 358924 371380
rect 198780 370772 198844 370836
rect 82676 370636 82740 370700
rect 213684 370636 213748 370700
rect 67772 370500 67836 370564
rect 250300 370500 250364 370564
rect 111564 369820 111628 369884
rect 121684 368460 121748 368524
rect 360332 368324 360396 368388
rect 200804 367780 200868 367844
rect 195100 366284 195164 366348
rect 118556 365664 118620 365668
rect 118556 365608 118606 365664
rect 118606 365608 118620 365664
rect 118556 365604 118620 365608
rect 81020 364924 81084 364988
rect 356284 364924 356348 364988
rect 114324 364244 114388 364308
rect 111748 363700 111812 363764
rect 190316 363700 190380 363764
rect 190316 363156 190380 363220
rect 240364 362476 240428 362540
rect 72740 362340 72804 362404
rect 154620 362340 154684 362404
rect 121684 362204 121748 362268
rect 67956 360844 68020 360908
rect 89668 360164 89732 360228
rect 206876 359484 206940 359548
rect 66116 359348 66180 359412
rect 69796 357444 69860 357508
rect 69060 354588 69124 354652
rect 69060 353908 69124 353972
rect 268332 353908 268396 353972
rect 180012 353500 180076 353564
rect 93716 353364 93780 353428
rect 209636 351324 209700 351388
rect 72924 350508 72988 350572
rect 286180 349828 286244 349892
rect 65932 347924 65996 347988
rect 99972 346972 100036 347036
rect 119476 345612 119540 345676
rect 66668 344388 66732 344452
rect 210740 344388 210804 344452
rect 291700 344388 291764 344452
rect 69612 344252 69676 344316
rect 286180 344312 286244 344316
rect 286180 344256 286230 344312
rect 286230 344256 286244 344312
rect 286180 344252 286244 344256
rect 157748 343028 157812 343092
rect 230428 342212 230492 342276
rect 354444 341532 354508 341596
rect 94452 340036 94516 340100
rect 109540 338404 109604 338468
rect 173204 338404 173268 338468
rect 170260 337316 170324 337380
rect 195100 337316 195164 337380
rect 188844 335956 188908 336020
rect 159404 335684 159468 335748
rect 241652 333372 241716 333436
rect 178540 331876 178604 331940
rect 162164 331332 162228 331396
rect 157932 330516 157996 330580
rect 252508 330516 252572 330580
rect 156828 329972 156892 330036
rect 69428 329564 69492 329628
rect 72924 329564 72988 329628
rect 75684 329428 75748 329492
rect 69428 328340 69492 328404
rect 156828 328204 156892 328268
rect 191604 326300 191668 326364
rect 69428 325484 69492 325548
rect 157748 325348 157812 325412
rect 157748 324396 157812 324460
rect 220860 323716 220924 323780
rect 247724 323716 247788 323780
rect 55076 320180 55140 320244
rect 281580 320180 281644 320244
rect 198412 318820 198476 318884
rect 191052 316780 191116 316844
rect 65932 315828 65996 315892
rect 242940 315012 243004 315076
rect 224172 314060 224236 314124
rect 161244 312564 161308 312628
rect 204484 311068 204548 311132
rect 352052 310388 352116 310452
rect 224724 309844 224788 309908
rect 179460 309028 179524 309092
rect 251220 308620 251284 308684
rect 157932 308484 157996 308548
rect 179460 308348 179524 308412
rect 180564 308348 180628 308412
rect 198596 307668 198660 307732
rect 159404 307124 159468 307188
rect 233740 306988 233804 307052
rect 219204 305628 219268 305692
rect 237420 303588 237484 303652
rect 304212 302228 304276 302292
rect 217548 301548 217612 301612
rect 244412 298284 244476 298348
rect 208164 297468 208228 297532
rect 199516 297332 199580 297396
rect 67956 296108 68020 296172
rect 214604 295972 214668 296036
rect 192340 295428 192404 295492
rect 255268 294068 255332 294132
rect 287100 293932 287164 293996
rect 169156 292572 169220 292636
rect 246804 291756 246868 291820
rect 198596 291076 198660 291140
rect 200620 291076 200684 291140
rect 246252 290048 246316 290052
rect 246252 289992 246302 290048
rect 246302 289992 246316 290048
rect 246252 289988 246316 289992
rect 191052 289852 191116 289916
rect 224172 289852 224236 289916
rect 187004 289776 187068 289780
rect 187004 289720 187054 289776
rect 187054 289720 187068 289776
rect 187004 289716 187068 289720
rect 160876 289172 160940 289236
rect 168972 289172 169036 289236
rect 238524 289172 238588 289236
rect 186820 289036 186884 289100
rect 226932 288492 226996 288556
rect 232084 287404 232148 287468
rect 283788 286316 283852 286380
rect 243676 285908 243740 285972
rect 212396 285772 212460 285836
rect 204484 285636 204548 285700
rect 218652 285636 218716 285700
rect 224172 285636 224236 285700
rect 228220 285636 228284 285700
rect 236500 285636 236564 285700
rect 192340 285092 192404 285156
rect 247724 285152 247788 285156
rect 247724 285096 247738 285152
rect 247738 285096 247788 285152
rect 247724 285092 247788 285096
rect 66668 284548 66732 284612
rect 244596 284412 244660 284476
rect 198780 284276 198844 284340
rect 192708 284004 192772 284068
rect 280292 284004 280356 284068
rect 205404 283928 205468 283932
rect 205404 283872 205418 283928
rect 205418 283872 205468 283928
rect 205404 283868 205468 283872
rect 214420 283928 214484 283932
rect 214420 283872 214470 283928
rect 214470 283872 214484 283928
rect 214420 283868 214484 283872
rect 216076 283928 216140 283932
rect 216076 283872 216126 283928
rect 216126 283872 216140 283928
rect 216076 283868 216140 283872
rect 222332 283868 222396 283932
rect 226012 283868 226076 283932
rect 229692 283868 229756 283932
rect 231900 283868 231964 283932
rect 236500 283868 236564 283932
rect 200068 283520 200132 283524
rect 200068 283464 200118 283520
rect 200118 283464 200132 283520
rect 200068 283460 200132 283464
rect 244596 283596 244660 283660
rect 198596 282916 198660 282980
rect 191788 282780 191852 282844
rect 192708 282780 192772 282844
rect 158484 281964 158548 282028
rect 195836 281556 195900 281620
rect 198780 281556 198844 281620
rect 199516 281556 199580 281620
rect 199332 281284 199396 281348
rect 200620 281284 200684 281348
rect 243492 281284 243556 281348
rect 69428 280740 69492 280804
rect 246252 280196 246316 280260
rect 156460 278020 156524 278084
rect 196940 277340 197004 277404
rect 200068 277340 200132 277404
rect 252508 275708 252572 275772
rect 65932 274136 65996 274140
rect 65932 274080 65946 274136
rect 65946 274080 65996 274136
rect 65932 274076 65996 274080
rect 248460 273124 248524 273188
rect 251220 273048 251284 273052
rect 251220 272992 251270 273048
rect 251270 272992 251284 273048
rect 251220 272988 251284 272992
rect 169524 271900 169588 271964
rect 181300 272444 181364 272508
rect 66116 271764 66180 271828
rect 191052 271084 191116 271148
rect 198412 270948 198476 271012
rect 250300 270404 250364 270468
rect 159956 270132 160020 270196
rect 163452 270132 163516 270196
rect 67772 269588 67836 269652
rect 260052 269180 260116 269244
rect 196756 268500 196820 268564
rect 196572 268364 196636 268428
rect 246804 267956 246868 268020
rect 67220 267412 67284 267476
rect 246620 267412 246684 267476
rect 246620 267004 246684 267068
rect 67772 266324 67836 266388
rect 197308 264148 197372 264212
rect 246804 263468 246868 263532
rect 197308 263060 197372 263124
rect 193812 262788 193876 262852
rect 244228 262516 244292 262580
rect 156828 261700 156892 261764
rect 249748 260884 249812 260948
rect 159220 260340 159284 260404
rect 244412 259524 244476 259588
rect 195100 259388 195164 259452
rect 191604 258708 191668 258772
rect 69428 255988 69492 256052
rect 191052 255580 191116 255644
rect 196940 255580 197004 255644
rect 243492 254084 243556 254148
rect 66668 252180 66732 252244
rect 199516 252180 199580 252244
rect 244044 251908 244108 251972
rect 243492 250004 243556 250068
rect 172468 249188 172532 249252
rect 199332 249052 199396 249116
rect 59124 247012 59188 247076
rect 245700 246468 245764 246532
rect 157932 246196 157996 246260
rect 191788 245652 191852 245716
rect 245700 245652 245764 245716
rect 199332 244836 199396 244900
rect 156828 244564 156892 244628
rect 191052 244564 191116 244628
rect 191788 244564 191852 244628
rect 200620 244020 200684 244084
rect 67220 243536 67284 243540
rect 67220 243480 67270 243536
rect 67270 243480 67284 243536
rect 67220 243476 67284 243480
rect 69428 243340 69492 243404
rect 192340 242116 192404 242180
rect 81020 242040 81084 242044
rect 81020 241984 81034 242040
rect 81034 241984 81084 242040
rect 81020 241980 81084 241984
rect 154620 242040 154684 242044
rect 154620 241984 154670 242040
rect 154670 241984 154684 242040
rect 154620 241980 154684 241984
rect 191788 241572 191852 241636
rect 83964 241300 84028 241364
rect 156460 241164 156524 241228
rect 156828 241028 156892 241092
rect 69612 240756 69676 240820
rect 302740 240756 302804 240820
rect 158484 240076 158548 240140
rect 208164 240076 208228 240140
rect 209636 240076 209700 240140
rect 210740 240136 210804 240140
rect 210740 240080 210754 240136
rect 210754 240080 210804 240136
rect 210740 240076 210804 240080
rect 213684 240076 213748 240140
rect 214604 240076 214668 240140
rect 217548 240136 217612 240140
rect 217548 240080 217562 240136
rect 217562 240080 217612 240136
rect 217548 240076 217612 240080
rect 219204 240076 219268 240140
rect 220860 240136 220924 240140
rect 220860 240080 220910 240136
rect 220910 240080 220924 240136
rect 220860 240076 220924 240080
rect 224724 240076 224788 240140
rect 226012 240076 226076 240140
rect 230428 240076 230492 240140
rect 232084 240076 232148 240140
rect 237420 240136 237484 240140
rect 237420 240080 237470 240136
rect 237470 240080 237484 240136
rect 237420 240076 237484 240080
rect 241652 240076 241716 240140
rect 243308 239940 243372 240004
rect 209636 238716 209700 238780
rect 206876 238580 206940 238644
rect 212396 238580 212460 238644
rect 244044 238036 244108 238100
rect 154068 237356 154132 237420
rect 199516 237356 199580 237420
rect 76420 237220 76484 237284
rect 216444 237356 216508 237420
rect 223620 237356 223684 237420
rect 242020 237356 242084 237420
rect 218652 237220 218716 237284
rect 193812 237084 193876 237148
rect 192340 236812 192404 236876
rect 82676 235860 82740 235924
rect 233740 235452 233804 235516
rect 205588 234636 205652 234700
rect 196756 234500 196820 234564
rect 188844 234364 188908 234428
rect 231900 234152 231964 234156
rect 231900 234096 231914 234152
rect 231914 234096 231964 234152
rect 231900 234092 231964 234096
rect 233004 234092 233068 234156
rect 191604 233820 191668 233884
rect 230428 233140 230492 233204
rect 193812 232596 193876 232660
rect 166212 231644 166276 231708
rect 205588 231508 205652 231572
rect 160876 230284 160940 230348
rect 175780 230148 175844 230212
rect 231900 229740 231964 229804
rect 412404 229740 412468 229804
rect 193812 228652 193876 228716
rect 179276 228380 179340 228444
rect 191052 228380 191116 228444
rect 244228 228380 244292 228444
rect 66668 228244 66732 228308
rect 414244 227020 414308 227084
rect 160692 226068 160756 226132
rect 184796 225932 184860 225996
rect 184796 225524 184860 225588
rect 298140 225524 298204 225588
rect 216076 224980 216140 225044
rect 169156 223348 169220 223412
rect 199332 222940 199396 223004
rect 195836 221852 195900 221916
rect 190316 220084 190380 220148
rect 234660 218588 234724 218652
rect 253060 217228 253124 217292
rect 69612 216276 69676 216340
rect 233188 216004 233252 216068
rect 222332 215248 222396 215252
rect 222332 215192 222382 215248
rect 222382 215192 222396 215248
rect 222332 215188 222396 215192
rect 161980 214916 162044 214980
rect 233004 214780 233068 214844
rect 232084 214372 232148 214436
rect 178540 212468 178604 212532
rect 223620 211108 223684 211172
rect 433380 210292 433444 210356
rect 173020 209340 173084 209404
rect 240364 207572 240428 207636
rect 214420 205728 214484 205732
rect 214420 205672 214470 205728
rect 214470 205672 214484 205728
rect 214420 205668 214484 205672
rect 216444 205396 216508 205460
rect 177804 202872 177868 202876
rect 177804 202816 177818 202872
rect 177818 202816 177868 202872
rect 177804 202812 177868 202816
rect 295932 202268 295996 202332
rect 157932 199956 157996 200020
rect 230612 199412 230676 199476
rect 244228 198732 244292 198796
rect 240732 198052 240796 198116
rect 245700 195876 245764 195940
rect 279004 195332 279068 195396
rect 284340 194516 284404 194580
rect 291148 192612 291212 192676
rect 244228 192476 244292 192540
rect 245700 191116 245764 191180
rect 287652 190980 287716 191044
rect 200620 189892 200684 189956
rect 75684 188260 75748 188324
rect 305500 187036 305564 187100
rect 299612 186900 299676 186964
rect 277164 186356 277228 186420
rect 285628 186356 285692 186420
rect 227668 185812 227732 185876
rect 237420 185676 237484 185740
rect 281764 185676 281828 185740
rect 188844 185540 188908 185604
rect 249932 185464 249996 185468
rect 249932 185408 249946 185464
rect 249946 185408 249996 185464
rect 249932 185404 249996 185408
rect 398604 184996 398668 185060
rect 162164 184316 162228 184380
rect 288572 183092 288636 183156
rect 159956 182956 160020 183020
rect 237604 181596 237668 181660
rect 298692 181460 298756 181524
rect 290596 180100 290660 180164
rect 180012 178740 180076 178804
rect 233372 178196 233436 178260
rect 112116 177924 112180 177988
rect 278820 178060 278884 178124
rect 280476 178060 280540 178124
rect 284524 177924 284588 177988
rect 98316 177516 98380 177580
rect 100708 177516 100772 177580
rect 105676 177516 105740 177580
rect 108068 177576 108132 177580
rect 108068 177520 108118 177576
rect 108118 177520 108132 177576
rect 108068 177516 108132 177520
rect 109540 177516 109604 177580
rect 114324 177576 114388 177580
rect 114324 177520 114374 177576
rect 114374 177520 114388 177576
rect 114324 177516 114388 177520
rect 121868 177516 121932 177580
rect 123156 177516 123220 177580
rect 124444 177516 124508 177580
rect 125732 177516 125796 177580
rect 130700 177516 130764 177580
rect 132356 177576 132420 177580
rect 132356 177520 132406 177576
rect 132406 177520 132420 177576
rect 132356 177516 132420 177520
rect 133092 177516 133156 177580
rect 148180 177516 148244 177580
rect 118372 177380 118436 177444
rect 104572 177244 104636 177308
rect 110644 177168 110708 177172
rect 110644 177112 110694 177168
rect 110694 177112 110708 177168
rect 110644 177108 110708 177112
rect 106964 176972 107028 177036
rect 164556 176972 164620 177036
rect 97028 176836 97092 176900
rect 101996 176836 102060 176900
rect 113220 176700 113284 176764
rect 115796 176760 115860 176764
rect 115796 176704 115846 176760
rect 115846 176704 115860 176760
rect 115796 176700 115860 176704
rect 119476 176760 119540 176764
rect 119476 176704 119526 176760
rect 119526 176704 119540 176760
rect 119476 176700 119540 176704
rect 120764 176760 120828 176764
rect 120764 176704 120814 176760
rect 120814 176704 120828 176760
rect 120764 176700 120828 176704
rect 127020 176760 127084 176764
rect 127020 176704 127070 176760
rect 127070 176704 127084 176760
rect 127020 176700 127084 176704
rect 129412 176760 129476 176764
rect 129412 176704 129462 176760
rect 129462 176704 129476 176760
rect 129412 176700 129476 176704
rect 158852 176700 158916 176764
rect 229140 176700 229204 176764
rect 226932 176564 226996 176628
rect 99420 176428 99484 176492
rect 103284 176428 103348 176492
rect 227668 176428 227732 176492
rect 228220 176292 228284 176356
rect 128124 175612 128188 175676
rect 116900 175476 116964 175540
rect 244228 175748 244292 175812
rect 277348 175748 277412 175812
rect 134380 175400 134444 175404
rect 134380 175344 134430 175400
rect 134430 175344 134444 175400
rect 134380 175340 134444 175344
rect 135668 175400 135732 175404
rect 135668 175344 135718 175400
rect 135718 175344 135732 175400
rect 135668 175340 135732 175344
rect 164556 174932 164620 174996
rect 280292 172484 280356 172548
rect 241652 168404 241716 168468
rect 280476 167860 280540 167924
rect 279372 167588 279436 167652
rect 236500 166772 236564 166836
rect 438900 166228 438964 166292
rect 233188 165684 233252 165748
rect 229140 163372 229204 163436
rect 281764 163236 281828 163300
rect 249012 161740 249076 161804
rect 248460 160652 248524 160716
rect 435036 159292 435100 159356
rect 281580 156436 281644 156500
rect 237604 156164 237668 156228
rect 238524 154396 238588 154460
rect 249932 153852 249996 153916
rect 244228 152492 244292 152556
rect 215892 150996 215956 151060
rect 230428 150588 230492 150652
rect 234660 149636 234724 149700
rect 264100 148956 264164 149020
rect 295932 149092 295996 149156
rect 237420 148276 237484 148340
rect 236500 146916 236564 146980
rect 230612 146296 230676 146300
rect 230612 146240 230626 146296
rect 230626 146240 230676 146296
rect 230612 146236 230676 146240
rect 232452 145556 232516 145620
rect 166212 144876 166276 144940
rect 231900 145284 231964 145348
rect 249748 144740 249812 144804
rect 231716 144060 231780 144124
rect 231716 142972 231780 143036
rect 230980 142836 231044 142900
rect 249012 142972 249076 143036
rect 242020 142836 242084 142900
rect 231164 142700 231228 142764
rect 244228 142488 244292 142492
rect 244228 142432 244278 142488
rect 244278 142432 244292 142488
rect 244228 142428 244292 142432
rect 424180 142156 424244 142220
rect 232084 142020 232148 142084
rect 237972 141340 238036 141404
rect 236500 141068 236564 141132
rect 440188 140796 440252 140860
rect 242020 140116 242084 140180
rect 441660 139980 441724 140044
rect 420868 139436 420932 139500
rect 425468 139496 425532 139500
rect 425468 139440 425518 139496
rect 425518 139440 425532 139496
rect 425468 139436 425532 139440
rect 426388 139436 426452 139500
rect 430620 139436 430684 139500
rect 436692 139436 436756 139500
rect 439084 139300 439148 139364
rect 233372 139164 233436 139228
rect 442028 138892 442092 138956
rect 245700 137804 245764 137868
rect 216812 137396 216876 137460
rect 229692 137260 229756 137324
rect 233740 135764 233804 135828
rect 398604 136172 398668 136236
rect 305500 135900 305564 135964
rect 284340 135084 284404 135148
rect 231164 134948 231228 135012
rect 249196 134404 249260 134468
rect 284524 134404 284588 134468
rect 285628 133588 285692 133652
rect 258580 132636 258644 132700
rect 229692 131412 229756 131476
rect 249012 130052 249076 130116
rect 267596 128420 267660 128484
rect 262812 127060 262876 127124
rect 360148 125428 360212 125492
rect 230980 125020 231044 125084
rect 353340 124068 353404 124132
rect 440188 121212 440252 121276
rect 439268 120804 439332 120868
rect 441660 119308 441724 119372
rect 230980 116180 231044 116244
rect 246252 116044 246316 116108
rect 439268 115908 439332 115972
rect 267780 113732 267844 113796
rect 266860 113324 266924 113388
rect 170260 112372 170324 112436
rect 439268 111284 439332 111348
rect 302740 111012 302804 111076
rect 283788 109924 283852 109988
rect 282132 109108 282196 109172
rect 397500 108292 397564 108356
rect 264100 107476 264164 107540
rect 232452 104212 232516 104276
rect 399892 103124 399956 103188
rect 170260 102444 170324 102508
rect 397500 102716 397564 102780
rect 258764 102308 258828 102372
rect 237972 102172 238036 102236
rect 290596 102172 290660 102236
rect 264100 101764 264164 101828
rect 287100 100948 287164 101012
rect 244228 100676 244292 100740
rect 260236 100132 260300 100196
rect 412404 99860 412468 99924
rect 414244 99860 414308 99924
rect 433380 99860 433444 99924
rect 435036 99860 435100 99924
rect 279372 99452 279436 99516
rect 400260 99180 400324 99244
rect 291700 97820 291764 97884
rect 434852 97880 434916 97884
rect 434852 97824 434866 97880
rect 434866 97824 434916 97880
rect 434852 97820 434916 97824
rect 229140 97004 229204 97068
rect 229140 96732 229204 96796
rect 255268 96460 255332 96524
rect 219204 95976 219268 95980
rect 219204 95920 219218 95976
rect 219218 95920 219268 95976
rect 219204 95916 219268 95920
rect 166396 95780 166460 95844
rect 224908 95508 224972 95572
rect 228956 95508 229020 95572
rect 205404 95100 205468 95164
rect 260052 94964 260116 95028
rect 100630 94752 100694 94756
rect 100630 94696 100666 94752
rect 100666 94696 100694 94752
rect 100630 94692 100694 94696
rect 120622 94752 120686 94756
rect 120622 94696 120630 94752
rect 120630 94696 120686 94752
rect 120622 94692 120686 94696
rect 151492 94692 151556 94756
rect 151766 94692 151830 94756
rect 267596 94420 267660 94484
rect 122052 94012 122116 94076
rect 114324 93876 114388 93940
rect 229692 93876 229756 93940
rect 95004 93740 95068 93804
rect 118188 93528 118252 93532
rect 118188 93472 118238 93528
rect 118238 93472 118252 93528
rect 118188 93468 118252 93472
rect 124076 93528 124140 93532
rect 124076 93472 124126 93528
rect 124126 93472 124140 93528
rect 124076 93468 124140 93472
rect 103284 93196 103348 93260
rect 110092 93256 110156 93260
rect 110092 93200 110142 93256
rect 110142 93200 110156 93256
rect 110092 93196 110156 93200
rect 115796 93060 115860 93124
rect 258764 93060 258828 93124
rect 286180 93060 286244 93124
rect 84332 92380 84396 92444
rect 108068 92440 108132 92444
rect 108068 92384 108118 92440
rect 108118 92384 108132 92440
rect 108068 92380 108132 92384
rect 110644 92380 110708 92444
rect 114876 92380 114940 92444
rect 116716 92440 116780 92444
rect 116716 92384 116766 92440
rect 116766 92384 116780 92440
rect 116716 92380 116780 92384
rect 125732 92440 125796 92444
rect 125732 92384 125782 92440
rect 125782 92384 125796 92440
rect 125732 92380 125796 92384
rect 133092 92440 133156 92444
rect 133092 92384 133142 92440
rect 133142 92384 133156 92440
rect 133092 92380 133156 92384
rect 120212 92244 120276 92308
rect 115428 92168 115492 92172
rect 115428 92112 115478 92168
rect 115478 92112 115492 92168
rect 115428 92108 115492 92112
rect 127572 92108 127636 92172
rect 104572 91972 104636 92036
rect 111196 91836 111260 91900
rect 100892 91700 100956 91764
rect 119660 91700 119724 91764
rect 130700 91760 130764 91764
rect 130700 91704 130750 91760
rect 130750 91704 130764 91760
rect 130700 91700 130764 91704
rect 151308 91700 151372 91764
rect 113220 91564 113284 91628
rect 99052 91428 99116 91492
rect 122788 91428 122852 91492
rect 85804 91292 85868 91356
rect 96660 91292 96724 91356
rect 101812 91292 101876 91356
rect 105492 91292 105556 91356
rect 106412 91292 106476 91356
rect 126468 91292 126532 91356
rect 151492 91352 151556 91356
rect 151492 91296 151542 91352
rect 151542 91296 151556 91352
rect 151492 91292 151556 91296
rect 74764 91156 74828 91220
rect 86724 91216 86788 91220
rect 86724 91160 86774 91216
rect 86774 91160 86788 91216
rect 86724 91156 86788 91160
rect 88012 91216 88076 91220
rect 88012 91160 88062 91216
rect 88062 91160 88076 91216
rect 88012 91156 88076 91160
rect 88932 91156 88996 91220
rect 90220 91156 90284 91220
rect 91324 91156 91388 91220
rect 92612 91156 92676 91220
rect 93900 91156 93964 91220
rect 96292 91216 96356 91220
rect 96292 91160 96342 91216
rect 96342 91160 96356 91216
rect 96292 91156 96356 91160
rect 97212 91156 97276 91220
rect 98132 91156 98196 91220
rect 99972 91156 100036 91220
rect 101996 91216 102060 91220
rect 101996 91160 102046 91216
rect 102046 91160 102060 91216
rect 101996 91156 102060 91160
rect 102732 91156 102796 91220
rect 104204 91156 104268 91220
rect 105676 91156 105740 91220
rect 106780 91156 106844 91220
rect 107700 91156 107764 91220
rect 109172 91216 109236 91220
rect 109172 91160 109222 91216
rect 109222 91160 109236 91216
rect 109172 91156 109236 91160
rect 109540 91156 109604 91220
rect 111932 91156 111996 91220
rect 112300 91156 112364 91220
rect 114324 91216 114388 91220
rect 114324 91160 114374 91216
rect 114374 91160 114388 91216
rect 114324 91156 114388 91160
rect 117084 91216 117148 91220
rect 117084 91160 117134 91216
rect 117134 91160 117148 91216
rect 117084 91156 117148 91160
rect 118004 91216 118068 91220
rect 118004 91160 118054 91216
rect 118054 91160 118068 91216
rect 118004 91156 118068 91160
rect 119292 91156 119356 91220
rect 121684 91156 121748 91220
rect 123156 91156 123220 91220
rect 125364 91216 125428 91220
rect 125364 91160 125414 91216
rect 125414 91160 125428 91216
rect 125364 91156 125428 91160
rect 126652 91156 126716 91220
rect 129412 91156 129476 91220
rect 132356 91216 132420 91220
rect 132356 91160 132406 91216
rect 132406 91160 132420 91216
rect 132356 91156 132420 91160
rect 134380 91156 134444 91220
rect 136036 91156 136100 91220
rect 151676 91216 151740 91220
rect 151676 91160 151726 91216
rect 151726 91160 151740 91216
rect 151676 91156 151740 91160
rect 152044 91156 152108 91220
rect 98500 91020 98564 91084
rect 124444 90884 124508 90948
rect 249196 90340 249260 90404
rect 442028 90340 442092 90404
rect 215892 89660 215956 89724
rect 304212 88980 304276 89044
rect 217180 88164 217244 88228
rect 282132 88164 282196 88228
rect 299612 86320 299676 86324
rect 299612 86264 299662 86320
rect 299662 86264 299676 86320
rect 299612 86260 299676 86264
rect 219204 84084 219268 84148
rect 264100 83404 264164 83468
rect 170260 81228 170324 81292
rect 166212 78508 166276 78572
rect 266860 77828 266924 77892
rect 426388 77828 426452 77892
rect 262812 76468 262876 76532
rect 166396 73068 166460 73132
rect 191052 69668 191116 69732
rect 430620 68172 430684 68236
rect 298140 66812 298204 66876
rect 291148 66132 291212 66196
rect 186820 64228 186884 64292
rect 267780 62732 267844 62796
rect 424180 60556 424244 60620
rect 436692 55796 436756 55860
rect 260236 53076 260300 53140
rect 233740 51716 233804 51780
rect 258580 44780 258644 44844
rect 249012 43420 249076 43484
rect 246252 39340 246316 39404
rect 224908 39204 224972 39268
rect 169524 37980 169588 38044
rect 65932 37844 65996 37908
rect 242020 36484 242084 36548
rect 439084 34444 439148 34508
rect 434852 30908 434916 30972
rect 281580 29548 281644 29612
rect 67772 24788 67836 24852
rect 287652 21388 287716 21452
rect 288756 21388 288820 21452
rect 172468 19892 172532 19956
rect 253060 19348 253124 19412
rect 55076 19212 55140 19276
rect 59124 15132 59188 15196
rect 425468 14452 425532 14516
rect 288756 12140 288820 12204
rect 299612 11732 299676 11796
rect 230980 11596 231044 11660
rect 288572 8196 288636 8260
rect 420868 7516 420932 7580
rect 188844 4932 188908 4996
rect 227668 4796 227732 4860
rect 298692 3980 298756 4044
rect 240732 3844 240796 3908
rect 268332 3436 268396 3500
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55075 320244 55141 320245
rect 55075 320180 55076 320244
rect 55140 320180 55141 320244
rect 55075 320179 55141 320180
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 55078 19277 55138 320179
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59123 247076 59189 247077
rect 59123 247012 59124 247076
rect 59188 247012 59189 247076
rect 59123 247011 59189 247012
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55075 19276 55141 19277
rect 55075 19212 55076 19276
rect 55140 19212 55141 19276
rect 55075 19211 55141 19212
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 -1306 56414 20898
rect 59126 15197 59186 247011
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59123 15196 59189 15197
rect 59123 15132 59124 15196
rect 59188 15132 59189 15196
rect 59123 15131 59189 15132
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 69611 702540 69677 702541
rect 69611 702476 69612 702540
rect 69676 702476 69677 702540
rect 69611 702475 69677 702476
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 591166 67574 608058
rect 69614 586530 69674 702475
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 591166 74414 614898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 591166 78134 618618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 591166 81854 622338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 591166 85574 626058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 88195 588572 88261 588573
rect 88195 588508 88196 588572
rect 88260 588508 88261 588572
rect 88195 588507 88261 588508
rect 69430 586470 69674 586530
rect 69430 582317 69490 586470
rect 88198 585717 88258 588507
rect 88195 585716 88261 585717
rect 88195 585652 88196 585716
rect 88260 585652 88261 585716
rect 88195 585651 88261 585652
rect 69427 582316 69493 582317
rect 69427 582252 69428 582316
rect 69492 582252 69493 582316
rect 69427 582251 69493 582252
rect 72679 579454 72999 579486
rect 72679 579218 72721 579454
rect 72957 579218 72999 579454
rect 72679 579134 72999 579218
rect 67771 578916 67837 578917
rect 67771 578852 67772 578916
rect 67836 578852 67837 578916
rect 72679 578898 72721 579134
rect 72957 578898 72999 579134
rect 72679 578866 72999 578898
rect 78609 579454 78929 579486
rect 78609 579218 78651 579454
rect 78887 579218 78929 579454
rect 78609 579134 78929 579218
rect 78609 578898 78651 579134
rect 78887 578898 78929 579134
rect 78609 578866 78929 578898
rect 84540 579454 84860 579486
rect 84540 579218 84582 579454
rect 84818 579218 84860 579454
rect 84540 579134 84860 579218
rect 84540 578898 84582 579134
rect 84818 578898 84860 579134
rect 84540 578866 84860 578898
rect 67771 578851 67837 578852
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 66667 556884 66733 556885
rect 66667 556820 66668 556884
rect 66732 556820 66733 556884
rect 66667 556819 66733 556820
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 66670 419661 66730 556819
rect 66954 536614 67574 537166
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 67774 535397 67834 578851
rect 75644 561454 75964 561486
rect 75644 561218 75686 561454
rect 75922 561218 75964 561454
rect 75644 561134 75964 561218
rect 75644 560898 75686 561134
rect 75922 560898 75964 561134
rect 75644 560866 75964 560898
rect 81575 561454 81895 561486
rect 81575 561218 81617 561454
rect 81853 561218 81895 561454
rect 81575 561134 81895 561218
rect 81575 560898 81617 561134
rect 81853 560898 81895 561134
rect 81575 560866 81895 560898
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91507 546548 91573 546549
rect 91507 546484 91508 546548
rect 91572 546484 91573 546548
rect 91507 546483 91573 546484
rect 72679 543454 72999 543486
rect 72679 543218 72721 543454
rect 72957 543218 72999 543454
rect 72679 543134 72999 543218
rect 68691 543012 68757 543013
rect 68691 542948 68692 543012
rect 68756 543010 68757 543012
rect 68756 542950 69122 543010
rect 68756 542948 68757 542950
rect 68691 542947 68757 542948
rect 67771 535396 67837 535397
rect 67771 535332 67772 535396
rect 67836 535332 67837 535396
rect 67771 535331 67837 535332
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 446407 67574 464058
rect 69062 452573 69122 542950
rect 72679 542898 72721 543134
rect 72957 542898 72999 543134
rect 72679 542866 72999 542898
rect 78609 543454 78929 543486
rect 78609 543218 78651 543454
rect 78887 543218 78929 543454
rect 78609 543134 78929 543218
rect 78609 542898 78651 543134
rect 78887 542898 78929 543134
rect 78609 542866 78929 542898
rect 84540 543454 84860 543486
rect 84540 543218 84582 543454
rect 84818 543218 84860 543454
rect 84540 543134 84860 543218
rect 84540 542898 84582 543134
rect 84818 542898 84860 543134
rect 84540 542866 84860 542898
rect 88195 541516 88261 541517
rect 88195 541452 88196 541516
rect 88260 541452 88261 541516
rect 88195 541451 88261 541452
rect 69611 535532 69677 535533
rect 69611 535468 69612 535532
rect 69676 535468 69677 535532
rect 69611 535467 69677 535468
rect 69059 452572 69125 452573
rect 69059 452508 69060 452572
rect 69124 452508 69125 452572
rect 69059 452507 69125 452508
rect 69062 451893 69122 452507
rect 69059 451892 69125 451893
rect 69059 451828 69060 451892
rect 69124 451828 69125 451892
rect 69059 451827 69125 451828
rect 66667 419660 66733 419661
rect 66667 419596 66668 419660
rect 66732 419596 66733 419660
rect 66667 419595 66733 419596
rect 67771 419660 67837 419661
rect 67771 419596 67772 419660
rect 67836 419596 67837 419660
rect 67771 419595 67837 419596
rect 65931 393276 65997 393277
rect 65931 393212 65932 393276
rect 65996 393212 65997 393276
rect 65931 393211 65997 393212
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 65934 347989 65994 393211
rect 66115 359412 66181 359413
rect 66115 359348 66116 359412
rect 66180 359348 66181 359412
rect 66115 359347 66181 359348
rect 65931 347988 65997 347989
rect 65931 347924 65932 347988
rect 65996 347924 65997 347988
rect 65931 347923 65997 347924
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 65934 315893 65994 347923
rect 65931 315892 65997 315893
rect 65931 315828 65932 315892
rect 65996 315828 65997 315892
rect 65931 315827 65997 315828
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 65931 274140 65997 274141
rect 65931 274076 65932 274140
rect 65996 274076 65997 274140
rect 65931 274075 65997 274076
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 65934 37909 65994 274075
rect 66118 271829 66178 359347
rect 66954 356614 67574 388356
rect 67774 378725 67834 419595
rect 69059 410004 69125 410005
rect 69059 409940 69060 410004
rect 69124 409940 69125 410004
rect 69059 409939 69125 409940
rect 67771 378724 67837 378725
rect 67771 378660 67772 378724
rect 67836 378660 67837 378724
rect 67771 378659 67837 378660
rect 67771 370564 67837 370565
rect 67771 370500 67772 370564
rect 67836 370500 67837 370564
rect 67771 370499 67837 370500
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66667 344452 66733 344453
rect 66667 344388 66668 344452
rect 66732 344388 66733 344452
rect 66667 344387 66733 344388
rect 66670 284613 66730 344387
rect 66954 331592 67574 356058
rect 66667 284612 66733 284613
rect 66667 284548 66668 284612
rect 66732 284548 66733 284612
rect 66667 284547 66733 284548
rect 66115 271828 66181 271829
rect 66115 271764 66116 271828
rect 66180 271764 66181 271828
rect 66115 271763 66181 271764
rect 67774 269653 67834 370499
rect 67955 360908 68021 360909
rect 67955 360844 67956 360908
rect 68020 360844 68021 360908
rect 67955 360843 68021 360844
rect 67958 296173 68018 360843
rect 69062 354653 69122 409939
rect 69614 390421 69674 535467
rect 73794 507454 74414 537166
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 72003 456108 72069 456109
rect 72003 456044 72004 456108
rect 72068 456044 72069 456108
rect 72003 456043 72069 456044
rect 71819 446452 71885 446453
rect 71819 446388 71820 446452
rect 71884 446388 71885 446452
rect 71819 446387 71885 446388
rect 71822 390557 71882 446387
rect 72006 445909 72066 456043
rect 73794 446407 74414 470898
rect 77514 511174 78134 537166
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 446407 78134 474618
rect 81234 514894 81854 537166
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 446407 81854 478338
rect 84954 518614 85574 537166
rect 88198 536757 88258 541451
rect 91510 541245 91570 546483
rect 91507 541244 91573 541245
rect 91507 541180 91508 541244
rect 91572 541180 91573 541244
rect 91507 541179 91573 541180
rect 88195 536756 88261 536757
rect 88195 536692 88196 536756
rect 88260 536692 88261 536756
rect 88195 536691 88261 536692
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446407 85574 482058
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 89667 469844 89733 469845
rect 89667 469780 89668 469844
rect 89732 469780 89733 469844
rect 89667 469779 89733 469780
rect 72003 445908 72069 445909
rect 72003 445844 72004 445908
rect 72068 445844 72069 445908
rect 72003 445843 72069 445844
rect 72739 445908 72805 445909
rect 72739 445844 72740 445908
rect 72804 445844 72805 445908
rect 72739 445843 72805 445844
rect 71819 390556 71885 390557
rect 71819 390492 71820 390556
rect 71884 390492 71885 390556
rect 71819 390491 71885 390492
rect 69611 390420 69677 390421
rect 69611 390356 69612 390420
rect 69676 390356 69677 390420
rect 69611 390355 69677 390356
rect 72742 362405 72802 445843
rect 72978 435454 73298 435486
rect 72978 435218 73020 435454
rect 73256 435218 73298 435454
rect 72978 435134 73298 435218
rect 72978 434898 73020 435134
rect 73256 434898 73298 435134
rect 72978 434866 73298 434898
rect 88338 417454 88658 417486
rect 88338 417218 88380 417454
rect 88616 417218 88658 417454
rect 88338 417134 88658 417218
rect 88338 416898 88380 417134
rect 88616 416898 88658 417134
rect 88338 416866 88658 416898
rect 72978 399454 73298 399486
rect 72978 399218 73020 399454
rect 73256 399218 73298 399454
rect 72978 399134 73298 399218
rect 72978 398898 73020 399134
rect 73256 398898 73298 399134
rect 72978 398866 73298 398898
rect 80467 391372 80533 391373
rect 80467 391308 80468 391372
rect 80532 391308 80533 391372
rect 80467 391307 80533 391308
rect 80470 390965 80530 391307
rect 80467 390964 80533 390965
rect 80467 390900 80468 390964
rect 80532 390900 80533 390964
rect 80467 390899 80533 390900
rect 89670 390421 89730 469779
rect 91139 458964 91205 458965
rect 91139 458900 91140 458964
rect 91204 458900 91205 458964
rect 91139 458899 91205 458900
rect 91142 390421 91202 458899
rect 91794 453454 92414 488898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 99971 538932 100037 538933
rect 99971 538868 99972 538932
rect 100036 538868 100037 538932
rect 99971 538867 100037 538868
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 96659 465764 96725 465765
rect 96659 465700 96660 465764
rect 96724 465700 96725 465764
rect 96659 465699 96725 465700
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 92611 456108 92677 456109
rect 92611 456044 92612 456108
rect 92676 456044 92677 456108
rect 92611 456043 92677 456044
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 446407 92414 452898
rect 92614 390421 92674 456043
rect 93899 449172 93965 449173
rect 93899 449108 93900 449172
rect 93964 449108 93965 449172
rect 93899 449107 93965 449108
rect 93715 445908 93781 445909
rect 93715 445844 93716 445908
rect 93780 445844 93781 445908
rect 93715 445843 93781 445844
rect 89667 390420 89733 390421
rect 89667 390356 89668 390420
rect 89732 390356 89733 390420
rect 89667 390355 89733 390356
rect 91139 390420 91205 390421
rect 91139 390356 91140 390420
rect 91204 390356 91205 390420
rect 91139 390355 91205 390356
rect 92611 390420 92677 390421
rect 92611 390356 92612 390420
rect 92676 390356 92677 390420
rect 92611 390355 92677 390356
rect 76419 390284 76485 390285
rect 76419 390220 76420 390284
rect 76484 390220 76485 390284
rect 76419 390219 76485 390220
rect 73794 363454 74414 388356
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 72739 362404 72805 362405
rect 72739 362340 72740 362404
rect 72804 362340 72805 362404
rect 72739 362339 72805 362340
rect 69795 357508 69861 357509
rect 69795 357444 69796 357508
rect 69860 357444 69861 357508
rect 69795 357443 69861 357444
rect 69059 354652 69125 354653
rect 69059 354588 69060 354652
rect 69124 354588 69125 354652
rect 69059 354587 69125 354588
rect 69062 353973 69122 354587
rect 69059 353972 69125 353973
rect 69059 353908 69060 353972
rect 69124 353908 69125 353972
rect 69059 353907 69125 353908
rect 69611 344316 69677 344317
rect 69611 344252 69612 344316
rect 69676 344252 69677 344316
rect 69611 344251 69677 344252
rect 69614 331230 69674 344251
rect 69246 331170 69674 331230
rect 69246 321570 69306 331170
rect 69427 329628 69493 329629
rect 69427 329564 69428 329628
rect 69492 329564 69493 329628
rect 69427 329563 69493 329564
rect 69430 328405 69490 329563
rect 69427 328404 69493 328405
rect 69427 328340 69428 328404
rect 69492 328340 69493 328404
rect 69427 328339 69493 328340
rect 69798 326770 69858 357443
rect 72923 350572 72989 350573
rect 72923 350508 72924 350572
rect 72988 350508 72989 350572
rect 72923 350507 72989 350508
rect 72926 329629 72986 350507
rect 73794 331592 74414 362898
rect 72923 329628 72989 329629
rect 72923 329564 72924 329628
rect 72988 329564 72989 329628
rect 72923 329563 72989 329564
rect 75683 329492 75749 329493
rect 75683 329428 75684 329492
rect 75748 329428 75749 329492
rect 75683 329427 75749 329428
rect 69430 326710 69858 326770
rect 69430 325549 69490 326710
rect 69427 325548 69493 325549
rect 69427 325484 69428 325548
rect 69492 325484 69493 325548
rect 69427 325483 69493 325484
rect 69246 321510 69674 321570
rect 67955 296172 68021 296173
rect 67955 296108 67956 296172
rect 68020 296108 68021 296172
rect 67955 296107 68021 296108
rect 69614 287070 69674 321510
rect 72978 291454 73298 291486
rect 72978 291218 73020 291454
rect 73256 291218 73298 291454
rect 72978 291134 73298 291218
rect 72978 290898 73020 291134
rect 73256 290898 73298 291134
rect 72978 290866 73298 290898
rect 69430 287010 69674 287070
rect 69430 280805 69490 287010
rect 69427 280804 69493 280805
rect 69427 280740 69428 280804
rect 69492 280740 69493 280804
rect 69427 280739 69493 280740
rect 67771 269652 67837 269653
rect 67771 269588 67772 269652
rect 67836 269588 67837 269652
rect 67771 269587 67837 269588
rect 67219 267476 67285 267477
rect 67219 267412 67220 267476
rect 67284 267412 67285 267476
rect 67219 267411 67285 267412
rect 66667 252244 66733 252245
rect 66667 252180 66668 252244
rect 66732 252180 66733 252244
rect 66667 252179 66733 252180
rect 66670 228309 66730 252179
rect 67222 243541 67282 267411
rect 67771 266388 67837 266389
rect 67771 266324 67772 266388
rect 67836 266324 67837 266388
rect 67771 266323 67837 266324
rect 67219 243540 67285 243541
rect 67219 243476 67220 243540
rect 67284 243476 67285 243540
rect 67219 243475 67285 243476
rect 66667 228308 66733 228309
rect 66667 228244 66668 228308
rect 66732 228244 66733 228308
rect 66667 228243 66733 228244
rect 66954 212614 67574 239592
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176600 67574 212058
rect 66954 68614 67574 93100
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 65931 37908 65997 37909
rect 65931 37844 65932 37908
rect 65996 37844 65997 37908
rect 65931 37843 65997 37844
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 67774 24853 67834 266323
rect 69427 256052 69493 256053
rect 69427 255988 69428 256052
rect 69492 255988 69493 256052
rect 69427 255987 69493 255988
rect 69430 248430 69490 255987
rect 72978 255454 73298 255486
rect 72978 255218 73020 255454
rect 73256 255218 73298 255454
rect 72978 255134 73298 255218
rect 72978 254898 73020 255134
rect 73256 254898 73298 255134
rect 72978 254866 73298 254898
rect 69430 248370 69674 248430
rect 69427 243404 69493 243405
rect 69427 243340 69428 243404
rect 69492 243340 69493 243404
rect 69427 243339 69493 243340
rect 69430 238770 69490 243339
rect 69614 240821 69674 248370
rect 69611 240820 69677 240821
rect 69611 240756 69612 240820
rect 69676 240756 69677 240820
rect 69611 240755 69677 240756
rect 69430 238710 69674 238770
rect 69614 216341 69674 238710
rect 73794 219454 74414 239592
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 69611 216340 69677 216341
rect 69611 216276 69612 216340
rect 69676 216276 69677 216340
rect 69611 216275 69677 216276
rect 73794 183454 74414 218898
rect 75686 188325 75746 329427
rect 76422 237285 76482 390219
rect 89670 389197 89730 390355
rect 89667 389196 89733 389197
rect 89667 389132 89668 389196
rect 89732 389132 89733 389196
rect 89667 389131 89733 389132
rect 83963 388788 84029 388789
rect 83963 388724 83964 388788
rect 84028 388724 84029 388788
rect 83963 388723 84029 388724
rect 77514 367174 78134 388356
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331592 78134 366618
rect 81234 370894 81854 388356
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 82675 370700 82741 370701
rect 82675 370636 82676 370700
rect 82740 370636 82741 370700
rect 82675 370635 82741 370636
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81019 364988 81085 364989
rect 81019 364924 81020 364988
rect 81084 364924 81085 364988
rect 81019 364923 81085 364924
rect 81022 242045 81082 364923
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 331592 81854 334338
rect 81019 242044 81085 242045
rect 81019 241980 81020 242044
rect 81084 241980 81085 242044
rect 81019 241979 81085 241980
rect 76419 237284 76485 237285
rect 76419 237220 76420 237284
rect 76484 237220 76485 237284
rect 76419 237219 76485 237220
rect 77514 223174 78134 239592
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 75683 188324 75749 188325
rect 75683 188260 75684 188324
rect 75748 188260 75749 188324
rect 75683 188259 75749 188260
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 176600 74414 182898
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 176600 78134 186618
rect 81234 226894 81854 239592
rect 82678 235925 82738 370635
rect 83966 241365 84026 388723
rect 84954 374614 85574 388356
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 89670 360229 89730 389131
rect 91794 381454 92414 388356
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 89667 360228 89733 360229
rect 89667 360164 89668 360228
rect 89732 360164 89733 360228
rect 89667 360163 89733 360164
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 331592 85574 338058
rect 91794 345454 92414 380898
rect 93718 353429 93778 445843
rect 93902 390421 93962 449107
rect 95187 447812 95253 447813
rect 95187 447748 95188 447812
rect 95252 447810 95253 447812
rect 95252 447750 95434 447810
rect 95252 447748 95253 447750
rect 95187 447747 95253 447748
rect 94451 444820 94517 444821
rect 94451 444756 94452 444820
rect 94516 444756 94517 444820
rect 94451 444755 94517 444756
rect 93899 390420 93965 390421
rect 93899 390356 93900 390420
rect 93964 390356 93965 390420
rect 93899 390355 93965 390356
rect 93715 353428 93781 353429
rect 93715 353364 93716 353428
rect 93780 353364 93781 353428
rect 93715 353363 93781 353364
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 331592 92414 344898
rect 94454 340101 94514 444755
rect 95374 390421 95434 447750
rect 95514 446407 96134 456618
rect 96662 390421 96722 465699
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 98131 457604 98197 457605
rect 98131 457540 98132 457604
rect 98196 457540 98197 457604
rect 98131 457539 98197 457540
rect 98134 390421 98194 457539
rect 99234 446407 99854 460338
rect 95371 390420 95437 390421
rect 95371 390356 95372 390420
rect 95436 390356 95437 390420
rect 95371 390355 95437 390356
rect 96659 390420 96725 390421
rect 96659 390356 96660 390420
rect 96724 390356 96725 390420
rect 96659 390355 96725 390356
rect 98131 390420 98197 390421
rect 98131 390356 98132 390420
rect 98196 390356 98197 390420
rect 98131 390355 98197 390356
rect 99974 388925 100034 538867
rect 102954 536614 103574 572058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 106411 538796 106477 538797
rect 106411 538732 106412 538796
rect 106476 538732 106477 538796
rect 106411 538731 106477 538732
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 100707 468484 100773 468485
rect 100707 468420 100708 468484
rect 100772 468420 100773 468484
rect 100707 468419 100773 468420
rect 100523 445772 100589 445773
rect 100523 445708 100524 445772
rect 100588 445708 100589 445772
rect 100523 445707 100589 445708
rect 99971 388924 100037 388925
rect 99971 388860 99972 388924
rect 100036 388860 100037 388924
rect 99971 388859 100037 388860
rect 95187 387836 95253 387837
rect 95187 387772 95188 387836
rect 95252 387772 95253 387836
rect 95187 387771 95253 387772
rect 95190 385661 95250 387771
rect 95187 385660 95253 385661
rect 95187 385596 95188 385660
rect 95252 385596 95253 385660
rect 95187 385595 95253 385596
rect 95514 385174 96134 388356
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 94451 340100 94517 340101
rect 94451 340036 94452 340100
rect 94516 340036 94517 340100
rect 94451 340035 94517 340036
rect 95514 331592 96134 348618
rect 99234 352894 99854 388356
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 331592 99854 352338
rect 99974 347037 100034 388859
rect 100526 387837 100586 445707
rect 100710 390421 100770 468419
rect 102954 464614 103574 500058
rect 104939 471204 105005 471205
rect 104939 471140 104940 471204
rect 105004 471140 105005 471204
rect 104939 471139 105005 471140
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102179 462908 102245 462909
rect 102179 462844 102180 462908
rect 102244 462844 102245 462908
rect 102179 462843 102245 462844
rect 102182 390421 102242 462843
rect 102954 446407 103574 464058
rect 103698 435454 104018 435486
rect 103698 435218 103740 435454
rect 103976 435218 104018 435454
rect 103698 435134 104018 435218
rect 103698 434898 103740 435134
rect 103976 434898 104018 435134
rect 103698 434866 104018 434898
rect 103698 399454 104018 399486
rect 103698 399218 103740 399454
rect 103976 399218 104018 399454
rect 103698 399134 104018 399218
rect 103698 398898 103740 399134
rect 103976 398898 104018 399134
rect 103698 398866 104018 398898
rect 104942 391101 105002 471139
rect 104939 391100 105005 391101
rect 104939 391036 104940 391100
rect 105004 391036 105005 391100
rect 104939 391035 105005 391036
rect 106414 390421 106474 538731
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 108987 467124 109053 467125
rect 108987 467060 108988 467124
rect 109052 467060 109053 467124
rect 108987 467059 109053 467060
rect 107699 465764 107765 465765
rect 107699 465700 107700 465764
rect 107764 465700 107765 465764
rect 107699 465699 107765 465700
rect 107702 390421 107762 465699
rect 108990 390557 109050 467059
rect 109794 446407 110414 470898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 115059 553484 115125 553485
rect 115059 553420 115060 553484
rect 115124 553420 115125 553484
rect 115059 553419 115125 553420
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 111747 457468 111813 457469
rect 111747 457404 111748 457468
rect 111812 457404 111813 457468
rect 111747 457403 111813 457404
rect 109539 444956 109605 444957
rect 109539 444892 109540 444956
rect 109604 444892 109605 444956
rect 109539 444891 109605 444892
rect 111563 444956 111629 444957
rect 111563 444892 111564 444956
rect 111628 444892 111629 444956
rect 111563 444891 111629 444892
rect 108987 390556 109053 390557
rect 108987 390492 108988 390556
rect 109052 390492 109053 390556
rect 108987 390491 109053 390492
rect 100707 390420 100773 390421
rect 100707 390356 100708 390420
rect 100772 390356 100773 390420
rect 100707 390355 100773 390356
rect 102179 390420 102245 390421
rect 102179 390356 102180 390420
rect 102244 390356 102245 390420
rect 102179 390355 102245 390356
rect 106411 390420 106477 390421
rect 106411 390356 106412 390420
rect 106476 390356 106477 390420
rect 106411 390355 106477 390356
rect 107699 390420 107765 390421
rect 107699 390356 107700 390420
rect 107764 390356 107765 390420
rect 107699 390355 107765 390356
rect 100523 387836 100589 387837
rect 100523 387772 100524 387836
rect 100588 387772 100589 387836
rect 100523 387771 100589 387772
rect 102954 356614 103574 388356
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 99971 347036 100037 347037
rect 99971 346972 99972 347036
rect 100036 346972 100037 347036
rect 99971 346971 100037 346972
rect 102954 331592 103574 356058
rect 109542 338469 109602 444891
rect 109794 363454 110414 388356
rect 111566 369885 111626 444891
rect 111750 389061 111810 457403
rect 113514 446407 114134 474618
rect 114323 445772 114389 445773
rect 114323 445708 114324 445772
rect 114388 445708 114389 445772
rect 114323 445707 114389 445708
rect 111747 389060 111813 389061
rect 111747 388996 111748 389060
rect 111812 388996 111813 389060
rect 111747 388995 111813 388996
rect 111563 369884 111629 369885
rect 111563 369820 111564 369884
rect 111628 369820 111629 369884
rect 111563 369819 111629 369820
rect 111750 363765 111810 388995
rect 113514 367174 114134 388356
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 111747 363764 111813 363765
rect 111747 363700 111748 363764
rect 111812 363700 111813 363764
rect 111747 363699 111813 363700
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109539 338468 109605 338469
rect 109539 338404 109540 338468
rect 109604 338404 109605 338468
rect 109539 338403 109605 338404
rect 109794 331592 110414 362898
rect 113514 331592 114134 366618
rect 114326 364309 114386 445707
rect 115062 388925 115122 553419
rect 117234 550894 117854 586338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 119475 579732 119541 579733
rect 119475 579668 119476 579732
rect 119540 579668 119541 579732
rect 119475 579667 119541 579668
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 115979 468484 116045 468485
rect 115979 468420 115980 468484
rect 116044 468420 116045 468484
rect 115979 468419 116045 468420
rect 115982 390421 116042 468419
rect 117234 446407 117854 478338
rect 118003 469844 118069 469845
rect 118003 469780 118004 469844
rect 118068 469780 118069 469844
rect 118003 469779 118069 469780
rect 118006 390421 118066 469779
rect 118555 445772 118621 445773
rect 118555 445708 118556 445772
rect 118620 445708 118621 445772
rect 118555 445707 118621 445708
rect 115979 390420 116045 390421
rect 115979 390356 115980 390420
rect 116044 390356 116045 390420
rect 115979 390355 116045 390356
rect 118003 390420 118069 390421
rect 118003 390356 118004 390420
rect 118068 390356 118069 390420
rect 118003 390355 118069 390356
rect 115059 388924 115125 388925
rect 115059 388860 115060 388924
rect 115124 388860 115125 388924
rect 115059 388859 115125 388860
rect 117234 370894 117854 388356
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 114323 364308 114389 364309
rect 114323 364244 114324 364308
rect 114388 364244 114389 364308
rect 114323 364243 114389 364244
rect 117234 334894 117854 370338
rect 118558 365669 118618 445707
rect 119478 436930 119538 579667
rect 120027 578372 120093 578373
rect 120027 578308 120028 578372
rect 120092 578308 120093 578372
rect 120027 578307 120093 578308
rect 120030 441630 120090 578307
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446407 121574 482058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 122603 449172 122669 449173
rect 122603 449108 122604 449172
rect 122668 449108 122669 449172
rect 122603 449107 122669 449108
rect 120030 441570 120458 441630
rect 119478 436870 120090 436930
rect 120030 431970 120090 436870
rect 120030 431910 120274 431970
rect 120214 430643 120274 431910
rect 120211 430642 120277 430643
rect 120211 430578 120212 430642
rect 120276 430578 120277 430642
rect 120211 430577 120277 430578
rect 119058 417454 119378 417486
rect 119058 417218 119100 417454
rect 119336 417218 119378 417454
rect 119058 417134 119378 417218
rect 119058 416898 119100 417134
rect 119336 416898 119378 417134
rect 119058 416866 119378 416898
rect 119475 392188 119541 392189
rect 119475 392124 119476 392188
rect 119540 392124 119541 392188
rect 119475 392123 119541 392124
rect 118555 365668 118621 365669
rect 118555 365604 118556 365668
rect 118620 365604 118621 365668
rect 118555 365603 118621 365604
rect 119478 345677 119538 392123
rect 120214 384301 120274 430577
rect 120398 428773 120458 441570
rect 120395 428772 120461 428773
rect 120395 428708 120396 428772
rect 120460 428708 120461 428772
rect 120395 428707 120461 428708
rect 122606 426325 122666 449107
rect 121683 426324 121749 426325
rect 121683 426260 121684 426324
rect 121748 426260 121749 426324
rect 121683 426259 121749 426260
rect 122603 426324 122669 426325
rect 122603 426260 122604 426324
rect 122668 426260 122669 426324
rect 122603 426259 122669 426260
rect 121499 419660 121565 419661
rect 121499 419596 121500 419660
rect 121564 419596 121565 419660
rect 121499 419595 121565 419596
rect 121502 390693 121562 419595
rect 121499 390692 121565 390693
rect 121499 390628 121500 390692
rect 121564 390628 121565 390692
rect 121499 390627 121565 390628
rect 120211 384300 120277 384301
rect 120211 384236 120212 384300
rect 120276 384236 120277 384300
rect 120211 384235 120277 384236
rect 120954 374614 121574 388356
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 119475 345676 119541 345677
rect 119475 345612 119476 345676
rect 119540 345612 119541 345676
rect 119475 345611 119541 345612
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 331592 117854 334338
rect 120954 338614 121574 374058
rect 121686 368525 121746 426259
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 122787 394772 122853 394773
rect 122787 394708 122788 394772
rect 122852 394708 122853 394772
rect 122787 394707 122853 394708
rect 122790 389190 122850 394707
rect 122606 389130 122850 389190
rect 122606 382941 122666 389130
rect 122603 382940 122669 382941
rect 122603 382876 122604 382940
rect 122668 382876 122669 382940
rect 122603 382875 122669 382876
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 121683 368524 121749 368525
rect 121683 368460 121684 368524
rect 121748 368460 121749 368524
rect 121683 368459 121749 368460
rect 121686 362269 121746 368459
rect 121683 362268 121749 362269
rect 121683 362204 121684 362268
rect 121748 362204 121749 362268
rect 121683 362203 121749 362204
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 331592 121574 338058
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 331592 128414 344898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 331592 132134 348618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 331592 135854 352338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 331592 139574 356058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 331592 146414 362898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331592 150134 366618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 160691 547908 160757 547909
rect 160691 547844 160692 547908
rect 160756 547844 160757 547908
rect 160691 547843 160757 547844
rect 159219 539748 159285 539749
rect 159219 539684 159220 539748
rect 159284 539684 159285 539748
rect 159219 539683 159285 539684
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156643 465220 156709 465221
rect 156643 465156 156644 465220
rect 156708 465156 156709 465220
rect 156643 465155 156709 465156
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 154067 442372 154133 442373
rect 154067 442308 154068 442372
rect 154132 442308 154133 442372
rect 154067 442307 154133 442308
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 331592 153854 334338
rect 88338 309454 88658 309486
rect 88338 309218 88380 309454
rect 88616 309218 88658 309454
rect 88338 309134 88658 309218
rect 88338 308898 88380 309134
rect 88616 308898 88658 309134
rect 88338 308866 88658 308898
rect 119058 309454 119378 309486
rect 119058 309218 119100 309454
rect 119336 309218 119378 309454
rect 119058 309134 119378 309218
rect 119058 308898 119100 309134
rect 119336 308898 119378 309134
rect 119058 308866 119378 308898
rect 149778 309454 150098 309486
rect 149778 309218 149820 309454
rect 150056 309218 150098 309454
rect 149778 309134 150098 309218
rect 149778 308898 149820 309134
rect 150056 308898 150098 309134
rect 149778 308866 150098 308898
rect 103698 291454 104018 291486
rect 103698 291218 103740 291454
rect 103976 291218 104018 291454
rect 103698 291134 104018 291218
rect 103698 290898 103740 291134
rect 103976 290898 104018 291134
rect 103698 290866 104018 290898
rect 134418 291454 134738 291486
rect 134418 291218 134460 291454
rect 134696 291218 134738 291454
rect 134418 291134 134738 291218
rect 134418 290898 134460 291134
rect 134696 290898 134738 291134
rect 134418 290866 134738 290898
rect 88338 273454 88658 273486
rect 88338 273218 88380 273454
rect 88616 273218 88658 273454
rect 88338 273134 88658 273218
rect 88338 272898 88380 273134
rect 88616 272898 88658 273134
rect 88338 272866 88658 272898
rect 119058 273454 119378 273486
rect 119058 273218 119100 273454
rect 119336 273218 119378 273454
rect 119058 273134 119378 273218
rect 119058 272898 119100 273134
rect 119336 272898 119378 273134
rect 119058 272866 119378 272898
rect 149778 273454 150098 273486
rect 149778 273218 149820 273454
rect 150056 273218 150098 273454
rect 149778 273134 150098 273218
rect 149778 272898 149820 273134
rect 150056 272898 150098 273134
rect 149778 272866 150098 272898
rect 103698 255454 104018 255486
rect 103698 255218 103740 255454
rect 103976 255218 104018 255454
rect 103698 255134 104018 255218
rect 103698 254898 103740 255134
rect 103976 254898 104018 255134
rect 103698 254866 104018 254898
rect 134418 255454 134738 255486
rect 134418 255218 134460 255454
rect 134696 255218 134738 255454
rect 134418 255134 134738 255218
rect 134418 254898 134460 255134
rect 134696 254898 134738 255134
rect 134418 254866 134738 254898
rect 83963 241364 84029 241365
rect 83963 241300 83964 241364
rect 84028 241300 84029 241364
rect 83963 241299 84029 241300
rect 82675 235924 82741 235925
rect 82675 235860 82676 235924
rect 82740 235860 82741 235924
rect 82675 235859 82741 235860
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 176600 81854 190338
rect 84954 230614 85574 239592
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 176600 85574 194058
rect 91794 237454 92414 239592
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 95514 205174 96134 239592
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 176600 96134 204618
rect 99234 208894 99854 239592
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 98315 177580 98381 177581
rect 98315 177516 98316 177580
rect 98380 177516 98381 177580
rect 98315 177515 98381 177516
rect 97027 176900 97093 176901
rect 97027 176836 97028 176900
rect 97092 176836 97093 176900
rect 97027 176835 97093 176836
rect 97030 175130 97090 176835
rect 96960 175070 97090 175130
rect 98318 175130 98378 177515
rect 99234 176600 99854 208338
rect 102954 212614 103574 239592
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 100707 177580 100773 177581
rect 100707 177516 100708 177580
rect 100772 177516 100773 177580
rect 100707 177515 100773 177516
rect 99419 176492 99485 176493
rect 99419 176428 99420 176492
rect 99484 176428 99485 176492
rect 99419 176427 99485 176428
rect 99422 175130 99482 176427
rect 98318 175070 98380 175130
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 177515
rect 101995 176900 102061 176901
rect 101995 176836 101996 176900
rect 102060 176836 102061 176900
rect 101995 176835 102061 176836
rect 101998 175130 102058 176835
rect 102954 176600 103574 212058
rect 109794 219454 110414 239592
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 105675 177580 105741 177581
rect 105675 177516 105676 177580
rect 105740 177516 105741 177580
rect 105675 177515 105741 177516
rect 108067 177580 108133 177581
rect 108067 177516 108068 177580
rect 108132 177516 108133 177580
rect 108067 177515 108133 177516
rect 109539 177580 109605 177581
rect 109539 177516 109540 177580
rect 109604 177516 109605 177580
rect 109539 177515 109605 177516
rect 104571 177308 104637 177309
rect 104571 177244 104572 177308
rect 104636 177244 104637 177308
rect 104571 177243 104637 177244
rect 103283 176492 103349 176493
rect 103283 176428 103284 176492
rect 103348 176428 103349 176492
rect 103283 176427 103349 176428
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176427
rect 104574 175130 104634 177243
rect 105678 175130 105738 177515
rect 106963 177036 107029 177037
rect 106963 176972 106964 177036
rect 107028 176972 107029 177036
rect 106963 176971 107029 176972
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 105738 175130
rect 106966 175130 107026 176971
rect 108070 175130 108130 177515
rect 109542 175130 109602 177515
rect 109794 176600 110414 182898
rect 113514 223174 114134 239592
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 112115 177988 112181 177989
rect 112115 177924 112116 177988
rect 112180 177924 112181 177988
rect 112115 177923 112181 177924
rect 110643 177172 110709 177173
rect 110643 177108 110644 177172
rect 110708 177108 110709 177172
rect 110643 177107 110709 177108
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109472 175070 109602 175130
rect 110646 175130 110706 177107
rect 112118 175130 112178 177923
rect 113219 176764 113285 176765
rect 113219 176700 113220 176764
rect 113284 176700 113285 176764
rect 113219 176699 113285 176700
rect 113222 175130 113282 176699
rect 113514 176600 114134 186618
rect 117234 226894 117854 239592
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 114323 177580 114389 177581
rect 114323 177516 114324 177580
rect 114388 177516 114389 177580
rect 114323 177515 114389 177516
rect 110646 175070 110756 175130
rect 109472 174494 109532 175070
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 113144 175070 113282 175130
rect 114326 175130 114386 177515
rect 115795 176764 115861 176765
rect 115795 176700 115796 176764
rect 115860 176700 115861 176764
rect 115795 176699 115861 176700
rect 115798 175130 115858 176699
rect 117234 176600 117854 190338
rect 120954 230614 121574 239592
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 118371 177444 118437 177445
rect 118371 177380 118372 177444
rect 118436 177380 118437 177444
rect 118371 177379 118437 177380
rect 116899 175540 116965 175541
rect 116899 175476 116900 175540
rect 116964 175476 116965 175540
rect 116899 175475 116965 175476
rect 114326 175070 114428 175130
rect 112056 174494 112116 175070
rect 113144 174494 113204 175070
rect 114368 174494 114428 175070
rect 115728 175070 115858 175130
rect 116902 175130 116962 175475
rect 118374 175130 118434 177379
rect 119475 176764 119541 176765
rect 119475 176700 119476 176764
rect 119540 176700 119541 176764
rect 119475 176699 119541 176700
rect 120763 176764 120829 176765
rect 120763 176700 120764 176764
rect 120828 176700 120829 176764
rect 120763 176699 120829 176700
rect 119478 175130 119538 176699
rect 120766 175130 120826 176699
rect 120954 176600 121574 194058
rect 127794 237454 128414 239592
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 121867 177580 121933 177581
rect 121867 177516 121868 177580
rect 121932 177516 121933 177580
rect 121867 177515 121933 177516
rect 123155 177580 123221 177581
rect 123155 177516 123156 177580
rect 123220 177516 123221 177580
rect 123155 177515 123221 177516
rect 124443 177580 124509 177581
rect 124443 177516 124444 177580
rect 124508 177516 124509 177580
rect 124443 177515 124509 177516
rect 125731 177580 125797 177581
rect 125731 177516 125732 177580
rect 125796 177516 125797 177580
rect 125731 177515 125797 177516
rect 121870 175130 121930 177515
rect 123158 175130 123218 177515
rect 124446 175130 124506 177515
rect 125734 175130 125794 177515
rect 127019 176764 127085 176765
rect 127019 176700 127020 176764
rect 127084 176700 127085 176764
rect 127019 176699 127085 176700
rect 127022 175130 127082 176699
rect 127794 176600 128414 200898
rect 131514 205174 132134 239592
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 130699 177580 130765 177581
rect 130699 177516 130700 177580
rect 130764 177516 130765 177580
rect 130699 177515 130765 177516
rect 129411 176764 129477 176765
rect 129411 176700 129412 176764
rect 129476 176700 129477 176764
rect 129411 176699 129477 176700
rect 128123 175676 128189 175677
rect 128123 175612 128124 175676
rect 128188 175612 128189 175676
rect 128123 175611 128189 175612
rect 128126 175130 128186 175611
rect 116902 175070 117012 175130
rect 115728 174494 115788 175070
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 119400 175070 119538 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 123072 175070 123218 175130
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 176699
rect 130702 175130 130762 177515
rect 131514 176600 132134 204618
rect 135234 208894 135854 239592
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 132355 177580 132421 177581
rect 132355 177516 132356 177580
rect 132420 177516 132421 177580
rect 132355 177515 132421 177516
rect 133091 177580 133157 177581
rect 133091 177516 133092 177580
rect 133156 177516 133157 177580
rect 133091 177515 133157 177516
rect 132358 175130 132418 177515
rect 129414 175070 129524 175130
rect 118312 174494 118372 175070
rect 119400 174494 119460 175070
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123072 174494 123132 175070
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 132048 175070 132418 175130
rect 133094 175130 133154 177515
rect 135234 176600 135854 208338
rect 138954 212614 139574 239592
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176600 139574 212058
rect 145794 219454 146414 239592
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 149514 223174 150134 239592
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 148179 177580 148245 177581
rect 148179 177516 148180 177580
rect 148244 177516 148245 177580
rect 148179 177515 148245 177516
rect 134379 175404 134445 175405
rect 134379 175340 134380 175404
rect 134444 175340 134445 175404
rect 134379 175339 134445 175340
rect 135667 175404 135733 175405
rect 135667 175340 135668 175404
rect 135732 175340 135733 175404
rect 135667 175339 135733 175340
rect 134382 175130 134442 175339
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 134360 175070 134442 175130
rect 135670 175130 135730 175339
rect 148182 175130 148242 177515
rect 149514 176600 150134 186618
rect 153234 226894 153854 239592
rect 154070 237421 154130 442307
rect 154619 362404 154685 362405
rect 154619 362340 154620 362404
rect 154684 362340 154685 362404
rect 154619 362339 154685 362340
rect 154622 242045 154682 362339
rect 156646 287070 156706 465155
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 157747 343092 157813 343093
rect 157747 343028 157748 343092
rect 157812 343028 157813 343092
rect 157747 343027 157813 343028
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 331592 157574 338058
rect 156827 330036 156893 330037
rect 156827 329972 156828 330036
rect 156892 329972 156893 330036
rect 156827 329971 156893 329972
rect 156830 328269 156890 329971
rect 156827 328268 156893 328269
rect 156827 328204 156828 328268
rect 156892 328204 156893 328268
rect 156827 328203 156893 328204
rect 157750 325413 157810 343027
rect 157931 330580 157997 330581
rect 157931 330516 157932 330580
rect 157996 330516 157997 330580
rect 157931 330515 157997 330516
rect 157747 325412 157813 325413
rect 157747 325348 157748 325412
rect 157812 325348 157813 325412
rect 157747 325347 157813 325348
rect 157750 324461 157810 325347
rect 157747 324460 157813 324461
rect 157747 324396 157748 324460
rect 157812 324396 157813 324460
rect 157747 324395 157813 324396
rect 157934 308549 157994 330515
rect 157931 308548 157997 308549
rect 157931 308484 157932 308548
rect 157996 308484 157997 308548
rect 157931 308483 157997 308484
rect 156646 287010 156890 287070
rect 156459 278084 156525 278085
rect 156459 278020 156460 278084
rect 156524 278020 156525 278084
rect 156459 278019 156525 278020
rect 154619 242044 154685 242045
rect 154619 241980 154620 242044
rect 154684 241980 154685 242044
rect 154619 241979 154685 241980
rect 156462 241229 156522 278019
rect 156830 261765 156890 287010
rect 158483 282028 158549 282029
rect 158483 281964 158484 282028
rect 158548 281964 158549 282028
rect 158483 281963 158549 281964
rect 156827 261764 156893 261765
rect 156827 261700 156828 261764
rect 156892 261700 156893 261764
rect 156827 261699 156893 261700
rect 157931 246260 157997 246261
rect 157931 246196 157932 246260
rect 157996 246196 157997 246260
rect 157931 246195 157997 246196
rect 156827 244628 156893 244629
rect 156827 244564 156828 244628
rect 156892 244564 156893 244628
rect 156827 244563 156893 244564
rect 156459 241228 156525 241229
rect 156459 241164 156460 241228
rect 156524 241164 156525 241228
rect 156459 241163 156525 241164
rect 156830 241093 156890 244563
rect 156827 241092 156893 241093
rect 156827 241028 156828 241092
rect 156892 241028 156893 241092
rect 156827 241027 156893 241028
rect 154067 237420 154133 237421
rect 154067 237356 154068 237420
rect 154132 237356 154133 237420
rect 154067 237355 154133 237356
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 176600 153854 190338
rect 156954 230614 157574 239592
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 157934 200021 157994 246195
rect 158486 240141 158546 281963
rect 159222 260405 159282 539683
rect 159403 335748 159469 335749
rect 159403 335684 159404 335748
rect 159468 335684 159469 335748
rect 159403 335683 159469 335684
rect 159406 307189 159466 335683
rect 159403 307188 159469 307189
rect 159403 307124 159404 307188
rect 159468 307124 159469 307188
rect 159403 307123 159469 307124
rect 159955 270196 160021 270197
rect 159955 270132 159956 270196
rect 160020 270132 160021 270196
rect 159955 270131 160021 270132
rect 159219 260404 159285 260405
rect 159219 260340 159220 260404
rect 159284 260340 159285 260404
rect 159219 260339 159285 260340
rect 158483 240140 158549 240141
rect 158483 240076 158484 240140
rect 158548 240076 158549 240140
rect 158483 240075 158549 240076
rect 157931 200020 157997 200021
rect 157931 199956 157932 200020
rect 157996 199956 157997 200020
rect 157931 199955 157997 199956
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 176600 157574 194058
rect 159958 183021 160018 270131
rect 160694 226133 160754 547843
rect 161243 542468 161309 542469
rect 161243 542404 161244 542468
rect 161308 542404 161309 542468
rect 161243 542403 161309 542404
rect 161246 312629 161306 542403
rect 163794 525454 164414 560898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 166211 557564 166277 557565
rect 166211 557500 166212 557564
rect 166276 557500 166277 557564
rect 166211 557499 166277 557500
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163451 518940 163517 518941
rect 163451 518876 163452 518940
rect 163516 518876 163517 518940
rect 163451 518875 163517 518876
rect 161979 514860 162045 514861
rect 161979 514796 161980 514860
rect 162044 514796 162045 514860
rect 161979 514795 162045 514796
rect 161243 312628 161309 312629
rect 161243 312564 161244 312628
rect 161308 312564 161309 312628
rect 161243 312563 161309 312564
rect 160875 289236 160941 289237
rect 160875 289172 160876 289236
rect 160940 289172 160941 289236
rect 160875 289171 160941 289172
rect 160878 230349 160938 289171
rect 160875 230348 160941 230349
rect 160875 230284 160876 230348
rect 160940 230284 160941 230348
rect 160875 230283 160941 230284
rect 160691 226132 160757 226133
rect 160691 226068 160692 226132
rect 160756 226068 160757 226132
rect 160691 226067 160757 226068
rect 161982 214981 162042 514795
rect 162163 331396 162229 331397
rect 162163 331332 162164 331396
rect 162228 331332 162229 331396
rect 162163 331331 162229 331332
rect 161979 214980 162045 214981
rect 161979 214916 161980 214980
rect 162044 214916 162045 214980
rect 161979 214915 162045 214916
rect 162166 184381 162226 331331
rect 163454 270197 163514 518875
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163451 270196 163517 270197
rect 163451 270132 163452 270196
rect 163516 270132 163517 270196
rect 163451 270131 163517 270132
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 166214 231709 166274 557499
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 168971 496908 169037 496909
rect 168971 496844 168972 496908
rect 169036 496844 169037 496908
rect 168971 496843 169037 496844
rect 171234 496894 171854 532338
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 168974 289237 169034 496843
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181299 543964 181365 543965
rect 181299 543900 181300 543964
rect 181364 543900 181365 543964
rect 181299 543899 181365 543900
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 175779 526420 175845 526421
rect 175779 526356 175780 526420
rect 175844 526356 175845 526420
rect 175779 526355 175845 526356
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 173019 401708 173085 401709
rect 173019 401644 173020 401708
rect 173084 401644 173085 401708
rect 173019 401643 173085 401644
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 170259 337380 170325 337381
rect 170259 337316 170260 337380
rect 170324 337316 170325 337380
rect 170259 337315 170325 337316
rect 169155 292636 169221 292637
rect 169155 292572 169156 292636
rect 169220 292572 169221 292636
rect 169155 292571 169221 292572
rect 168971 289236 169037 289237
rect 168971 289172 168972 289236
rect 169036 289172 169037 289236
rect 168971 289171 169037 289172
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 166211 231708 166277 231709
rect 166211 231644 166212 231708
rect 166276 231644 166277 231708
rect 166211 231643 166277 231644
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 162163 184380 162229 184381
rect 162163 184316 162164 184380
rect 162228 184316 162229 184380
rect 162163 184315 162229 184316
rect 159955 183020 160021 183021
rect 159955 182956 159956 183020
rect 160020 182956 160021 183020
rect 159955 182955 160021 182956
rect 158851 176764 158917 176765
rect 158851 176700 158852 176764
rect 158916 176700 158917 176764
rect 158851 176699 158917 176700
rect 158854 175130 158914 176699
rect 163794 176600 164414 200898
rect 167514 205174 168134 240618
rect 169158 223413 169218 292571
rect 169523 271964 169589 271965
rect 169523 271900 169524 271964
rect 169588 271900 169589 271964
rect 169523 271899 169589 271900
rect 169155 223412 169221 223413
rect 169155 223348 169156 223412
rect 169220 223348 169221 223412
rect 169155 223347 169221 223348
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 164555 177036 164621 177037
rect 164555 176972 164556 177036
rect 164620 176972 164621 177036
rect 164555 176971 164621 176972
rect 135670 175070 135780 175130
rect 148182 175070 148292 175130
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 164558 174997 164618 176971
rect 164555 174996 164621 174997
rect 164555 174932 164556 174996
rect 164620 174932 164621 174996
rect 164555 174931 164621 174932
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 69072 165454 69420 165486
rect 69072 165218 69128 165454
rect 69364 165218 69420 165454
rect 69072 165134 69420 165218
rect 69072 164898 69128 165134
rect 69364 164898 69420 165134
rect 69072 164866 69420 164898
rect 164136 165454 164484 165486
rect 164136 165218 164192 165454
rect 164428 165218 164484 165454
rect 164136 165134 164484 165218
rect 164136 164898 164192 165134
rect 164428 164898 164484 165134
rect 164136 164866 164484 164898
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 166211 144940 166277 144941
rect 166211 144876 166212 144940
rect 166276 144876 166277 144940
rect 166211 144875 166277 144876
rect 69072 129454 69420 129486
rect 69072 129218 69128 129454
rect 69364 129218 69420 129454
rect 69072 129134 69420 129218
rect 69072 128898 69128 129134
rect 69364 128898 69420 129134
rect 69072 128866 69420 128898
rect 164136 129454 164484 129486
rect 164136 129218 164192 129454
rect 164428 129218 164484 129454
rect 164136 129134 164484 129218
rect 164136 128898 164192 129134
rect 164428 128898 164484 129134
rect 164136 128866 164484 128898
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 85536 94890 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 85536 94830 85866 94890
rect 86624 94830 86786 94890
rect 87984 94830 88074 94890
rect 73794 75454 74414 93100
rect 74766 91221 74826 94830
rect 74763 91220 74829 91221
rect 74763 91156 74764 91220
rect 74828 91156 74829 91220
rect 74763 91155 74829 91156
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 67771 24852 67837 24853
rect 67771 24788 67772 24852
rect 67836 24788 67837 24852
rect 67771 24787 67837 24788
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 93100
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 93100
rect 84334 92445 84394 94830
rect 84331 92444 84397 92445
rect 84331 92380 84332 92444
rect 84396 92380 84397 92444
rect 84331 92379 84397 92380
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 93100
rect 85806 91357 85866 94830
rect 85803 91356 85869 91357
rect 85803 91292 85804 91356
rect 85868 91292 85869 91356
rect 85803 91291 85869 91292
rect 86726 91221 86786 94830
rect 88014 91221 88074 94830
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 88934 91221 88994 94830
rect 90222 91221 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 94920 94890 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 94920 94830 95066 94890
rect 96008 94830 96354 94890
rect 91326 91221 91386 94830
rect 86723 91220 86789 91221
rect 86723 91156 86724 91220
rect 86788 91156 86789 91220
rect 86723 91155 86789 91156
rect 88011 91220 88077 91221
rect 88011 91156 88012 91220
rect 88076 91156 88077 91220
rect 88011 91155 88077 91156
rect 88931 91220 88997 91221
rect 88931 91156 88932 91220
rect 88996 91156 88997 91220
rect 88931 91155 88997 91156
rect 90219 91220 90285 91221
rect 90219 91156 90220 91220
rect 90284 91156 90285 91220
rect 90219 91155 90285 91156
rect 91323 91220 91389 91221
rect 91323 91156 91324 91220
rect 91388 91156 91389 91220
rect 91323 91155 91389 91156
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 93100
rect 92614 91221 92674 94830
rect 93902 91221 93962 94830
rect 95006 93805 95066 94830
rect 95003 93804 95069 93805
rect 95003 93740 95004 93804
rect 95068 93740 95069 93804
rect 95003 93739 95069 93740
rect 92611 91220 92677 91221
rect 92611 91156 92612 91220
rect 92676 91156 92677 91220
rect 92611 91155 92677 91156
rect 93899 91220 93965 91221
rect 93899 91156 93900 91220
rect 93964 91156 93965 91220
rect 93899 91155 93965 91156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 93100
rect 96294 91221 96354 94830
rect 96662 94830 96748 94890
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 96662 91357 96722 94830
rect 96659 91356 96725 91357
rect 96659 91292 96660 91356
rect 96724 91292 96725 91356
rect 96659 91291 96725 91292
rect 97214 91221 97274 94830
rect 98134 91221 98194 94830
rect 96291 91220 96357 91221
rect 96291 91156 96292 91220
rect 96356 91156 96357 91220
rect 96291 91155 96357 91156
rect 97211 91220 97277 91221
rect 97211 91156 97212 91220
rect 97276 91156 97277 91220
rect 97211 91155 97277 91156
rect 98131 91220 98197 91221
rect 98131 91156 98132 91220
rect 98196 91156 98197 91220
rect 98131 91155 98197 91156
rect 98502 91085 98562 94830
rect 99054 94830 99196 94890
rect 99544 94890 99604 95200
rect 99544 94830 100034 94890
rect 99054 91493 99114 94830
rect 99051 91492 99117 91493
rect 99051 91428 99052 91492
rect 99116 91428 99117 91492
rect 99051 91427 99117 91428
rect 98499 91084 98565 91085
rect 98499 91020 98500 91084
rect 98564 91020 98565 91084
rect 98499 91019 98565 91020
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 93100
rect 99974 91221 100034 94830
rect 100632 94757 100692 95200
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 100954 94890
rect 100629 94756 100695 94757
rect 100629 94692 100630 94756
rect 100694 94692 100695 94756
rect 100629 94691 100695 94692
rect 100894 91765 100954 94830
rect 101814 94830 101916 94890
rect 101992 94890 102052 95200
rect 102944 94890 103004 95200
rect 101992 94830 102058 94890
rect 100891 91764 100957 91765
rect 100891 91700 100892 91764
rect 100956 91700 100957 91764
rect 100891 91699 100957 91700
rect 101814 91357 101874 94830
rect 101811 91356 101877 91357
rect 101811 91292 101812 91356
rect 101876 91292 101877 91356
rect 101811 91291 101877 91292
rect 101998 91221 102058 94830
rect 102734 94830 103004 94890
rect 103216 94890 103276 95200
rect 104304 94890 104364 95200
rect 103216 94830 103346 94890
rect 102734 91221 102794 94830
rect 103286 93261 103346 94830
rect 104206 94830 104364 94890
rect 104440 94890 104500 95200
rect 105392 94890 105452 95200
rect 105664 94890 105724 95200
rect 106480 94890 106540 95200
rect 104440 94830 104634 94890
rect 105392 94830 105554 94890
rect 105664 94830 105738 94890
rect 103283 93260 103349 93261
rect 103283 93196 103284 93260
rect 103348 93196 103349 93260
rect 103283 93195 103349 93196
rect 99971 91220 100037 91221
rect 99971 91156 99972 91220
rect 100036 91156 100037 91220
rect 99971 91155 100037 91156
rect 101995 91220 102061 91221
rect 101995 91156 101996 91220
rect 102060 91156 102061 91220
rect 101995 91155 102061 91156
rect 102731 91220 102797 91221
rect 102731 91156 102732 91220
rect 102796 91156 102797 91220
rect 102731 91155 102797 91156
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 93100
rect 104206 91221 104266 94830
rect 104574 92037 104634 94830
rect 104571 92036 104637 92037
rect 104571 91972 104572 92036
rect 104636 91972 104637 92036
rect 104571 91971 104637 91972
rect 105494 91357 105554 94830
rect 105491 91356 105557 91357
rect 105491 91292 105492 91356
rect 105556 91292 105557 91356
rect 105491 91291 105557 91292
rect 105678 91221 105738 94830
rect 106414 94830 106540 94890
rect 106616 94890 106676 95200
rect 107704 94890 107764 95200
rect 108112 94890 108172 95200
rect 106616 94830 106842 94890
rect 106414 91357 106474 94830
rect 106411 91356 106477 91357
rect 106411 91292 106412 91356
rect 106476 91292 106477 91356
rect 106411 91291 106477 91292
rect 106782 91221 106842 94830
rect 107702 94830 107764 94890
rect 108070 94830 108172 94890
rect 109064 94890 109124 95200
rect 109472 94890 109532 95200
rect 110152 94890 110212 95200
rect 110696 94890 110756 95200
rect 111240 94890 111300 95200
rect 109064 94830 109234 94890
rect 109472 94830 109602 94890
rect 107702 91221 107762 94830
rect 108070 92445 108130 94830
rect 108067 92444 108133 92445
rect 108067 92380 108068 92444
rect 108132 92380 108133 92444
rect 108067 92379 108133 92380
rect 109174 91221 109234 94830
rect 109542 91221 109602 94830
rect 110094 94830 110212 94890
rect 110646 94830 110756 94890
rect 111198 94830 111300 94890
rect 111920 94890 111980 95200
rect 112328 94890 112388 95200
rect 111920 94830 111994 94890
rect 110094 93261 110154 94830
rect 110091 93260 110157 93261
rect 110091 93196 110092 93260
rect 110156 93196 110157 93260
rect 110091 93195 110157 93196
rect 104203 91220 104269 91221
rect 104203 91156 104204 91220
rect 104268 91156 104269 91220
rect 104203 91155 104269 91156
rect 105675 91220 105741 91221
rect 105675 91156 105676 91220
rect 105740 91156 105741 91220
rect 105675 91155 105741 91156
rect 106779 91220 106845 91221
rect 106779 91156 106780 91220
rect 106844 91156 106845 91220
rect 106779 91155 106845 91156
rect 107699 91220 107765 91221
rect 107699 91156 107700 91220
rect 107764 91156 107765 91220
rect 107699 91155 107765 91156
rect 109171 91220 109237 91221
rect 109171 91156 109172 91220
rect 109236 91156 109237 91220
rect 109171 91155 109237 91156
rect 109539 91220 109605 91221
rect 109539 91156 109540 91220
rect 109604 91156 109605 91220
rect 109539 91155 109605 91156
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 93100
rect 110646 92445 110706 94830
rect 110643 92444 110709 92445
rect 110643 92380 110644 92444
rect 110708 92380 110709 92444
rect 110643 92379 110709 92380
rect 111198 91901 111258 94830
rect 111195 91900 111261 91901
rect 111195 91836 111196 91900
rect 111260 91836 111261 91900
rect 111195 91835 111261 91836
rect 111934 91221 111994 94830
rect 112302 94830 112388 94890
rect 113144 94890 113204 95200
rect 113688 94890 113748 95200
rect 114368 94890 114428 95200
rect 113144 94830 113282 94890
rect 113688 94830 114202 94890
rect 112302 91221 112362 94830
rect 113222 91629 113282 94830
rect 114142 93530 114202 94830
rect 114326 94830 114428 94890
rect 114776 94890 114836 95200
rect 115456 94890 115516 95200
rect 115864 94890 115924 95200
rect 114776 94830 114938 94890
rect 114326 93941 114386 94830
rect 114323 93940 114389 93941
rect 114323 93876 114324 93940
rect 114388 93876 114389 93940
rect 114323 93875 114389 93876
rect 114142 93470 114386 93530
rect 113219 91628 113285 91629
rect 113219 91564 113220 91628
rect 113284 91564 113285 91628
rect 113219 91563 113285 91564
rect 111931 91220 111997 91221
rect 111931 91156 111932 91220
rect 111996 91156 111997 91220
rect 111931 91155 111997 91156
rect 112299 91220 112365 91221
rect 112299 91156 112300 91220
rect 112364 91156 112365 91220
rect 112299 91155 112365 91156
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 79174 114134 93100
rect 114326 91221 114386 93470
rect 114878 92445 114938 94830
rect 115430 94830 115516 94890
rect 115798 94830 115924 94890
rect 116680 94890 116740 95200
rect 117088 94890 117148 95200
rect 116680 94830 116778 94890
rect 114875 92444 114941 92445
rect 114875 92380 114876 92444
rect 114940 92380 114941 92444
rect 114875 92379 114941 92380
rect 115430 92173 115490 94830
rect 115798 93125 115858 94830
rect 115795 93124 115861 93125
rect 115795 93060 115796 93124
rect 115860 93060 115861 93124
rect 115795 93059 115861 93060
rect 116718 92445 116778 94830
rect 117086 94830 117148 94890
rect 117904 94890 117964 95200
rect 118176 94890 118236 95200
rect 119400 94890 119460 95200
rect 117904 94830 118066 94890
rect 118176 94830 118250 94890
rect 116715 92444 116781 92445
rect 116715 92380 116716 92444
rect 116780 92380 116781 92444
rect 116715 92379 116781 92380
rect 115427 92172 115493 92173
rect 115427 92108 115428 92172
rect 115492 92108 115493 92172
rect 115427 92107 115493 92108
rect 117086 91221 117146 94830
rect 114323 91220 114389 91221
rect 114323 91156 114324 91220
rect 114388 91156 114389 91220
rect 114323 91155 114389 91156
rect 117083 91220 117149 91221
rect 117083 91156 117084 91220
rect 117148 91156 117149 91220
rect 117083 91155 117149 91156
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 82894 117854 93100
rect 118006 91221 118066 94830
rect 118190 93533 118250 94830
rect 119294 94830 119460 94890
rect 119536 94890 119596 95200
rect 120216 94890 120276 95200
rect 119536 94830 119722 94890
rect 118187 93532 118253 93533
rect 118187 93468 118188 93532
rect 118252 93468 118253 93532
rect 118187 93467 118253 93468
rect 119294 91221 119354 94830
rect 119662 91765 119722 94830
rect 120214 94830 120276 94890
rect 120214 92309 120274 94830
rect 120624 94757 120684 95200
rect 121712 94890 121772 95200
rect 121686 94830 121772 94890
rect 121984 94890 122044 95200
rect 122800 94890 122860 95200
rect 123208 94890 123268 95200
rect 121984 94830 122114 94890
rect 122800 94830 123034 94890
rect 120621 94756 120687 94757
rect 120621 94692 120622 94756
rect 120686 94692 120687 94756
rect 120621 94691 120687 94692
rect 120211 92308 120277 92309
rect 120211 92244 120212 92308
rect 120276 92244 120277 92308
rect 120211 92243 120277 92244
rect 119659 91764 119725 91765
rect 119659 91700 119660 91764
rect 119724 91700 119725 91764
rect 119659 91699 119725 91700
rect 118003 91220 118069 91221
rect 118003 91156 118004 91220
rect 118068 91156 118069 91220
rect 118003 91155 118069 91156
rect 119291 91220 119357 91221
rect 119291 91156 119292 91220
rect 119356 91156 119357 91220
rect 119291 91155 119357 91156
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 86614 121574 93100
rect 121686 91221 121746 94830
rect 122054 94077 122114 94830
rect 122051 94076 122117 94077
rect 122051 94012 122052 94076
rect 122116 94012 122117 94076
rect 122051 94011 122117 94012
rect 122974 93870 123034 94830
rect 122606 93810 123034 93870
rect 123158 94830 123268 94890
rect 124024 94890 124084 95200
rect 124432 94890 124492 95200
rect 125384 94890 125444 95200
rect 124024 94830 124138 94890
rect 124432 94830 124506 94890
rect 122606 91490 122666 93810
rect 122787 91492 122853 91493
rect 122787 91490 122788 91492
rect 122606 91430 122788 91490
rect 122787 91428 122788 91430
rect 122852 91428 122853 91492
rect 122787 91427 122853 91428
rect 123158 91221 123218 94830
rect 124078 93533 124138 94830
rect 124075 93532 124141 93533
rect 124075 93468 124076 93532
rect 124140 93468 124141 93532
rect 124075 93467 124141 93468
rect 121683 91220 121749 91221
rect 121683 91156 121684 91220
rect 121748 91156 121749 91220
rect 121683 91155 121749 91156
rect 123155 91220 123221 91221
rect 123155 91156 123156 91220
rect 123220 91156 123221 91220
rect 123155 91155 123221 91156
rect 124446 90949 124506 94830
rect 125366 94830 125444 94890
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125794 94890
rect 125366 91221 125426 94830
rect 125734 92445 125794 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 126608 94830 126714 94890
rect 125731 92444 125797 92445
rect 125731 92380 125732 92444
rect 125796 92380 125797 92444
rect 125731 92379 125797 92380
rect 126470 91357 126530 94830
rect 126467 91356 126533 91357
rect 126467 91292 126468 91356
rect 126532 91292 126533 91356
rect 126467 91291 126533 91292
rect 126654 91221 126714 94830
rect 127574 94830 128164 94890
rect 129328 94890 129388 95200
rect 130688 94890 130748 95200
rect 131912 94890 131972 95200
rect 133136 94890 133196 95200
rect 129328 94830 129474 94890
rect 130688 94830 130762 94890
rect 131912 94830 132418 94890
rect 127574 92173 127634 94830
rect 127571 92172 127637 92173
rect 127571 92108 127572 92172
rect 127636 92108 127637 92172
rect 127571 92107 127637 92108
rect 125363 91220 125429 91221
rect 125363 91156 125364 91220
rect 125428 91156 125429 91220
rect 125363 91155 125429 91156
rect 126651 91220 126717 91221
rect 126651 91156 126652 91220
rect 126716 91156 126717 91220
rect 126651 91155 126717 91156
rect 124443 90948 124509 90949
rect 124443 90884 124444 90948
rect 124508 90884 124509 90948
rect 124443 90883 124509 90884
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 93100
rect 129414 91221 129474 94830
rect 130702 91765 130762 94830
rect 130699 91764 130765 91765
rect 130699 91700 130700 91764
rect 130764 91700 130765 91764
rect 130699 91699 130765 91700
rect 129411 91220 129477 91221
rect 129411 91156 129412 91220
rect 129476 91156 129477 91220
rect 129411 91155 129477 91156
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 61174 132134 93100
rect 132358 91221 132418 94830
rect 133094 94830 133196 94890
rect 134360 94890 134420 95200
rect 135584 94890 135644 95200
rect 151496 94890 151556 95200
rect 134360 94830 134442 94890
rect 135584 94830 136098 94890
rect 133094 92445 133154 94830
rect 133091 92444 133157 92445
rect 133091 92380 133092 92444
rect 133156 92380 133157 92444
rect 133091 92379 133157 92380
rect 134382 91221 134442 94830
rect 132355 91220 132421 91221
rect 132355 91156 132356 91220
rect 132420 91156 132421 91220
rect 132355 91155 132421 91156
rect 134379 91220 134445 91221
rect 134379 91156 134380 91220
rect 134444 91156 134445 91220
rect 134379 91155 134445 91156
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 64894 135854 93100
rect 136038 91221 136098 94830
rect 151310 94830 151556 94890
rect 136035 91220 136101 91221
rect 136035 91156 136036 91220
rect 136100 91156 136101 91220
rect 136035 91155 136101 91156
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 93100
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 79174 150134 93100
rect 151310 91765 151370 94830
rect 151491 94756 151557 94757
rect 151491 94692 151492 94756
rect 151556 94692 151557 94756
rect 151491 94691 151557 94692
rect 151307 91764 151373 91765
rect 151307 91700 151308 91764
rect 151372 91700 151373 91764
rect 151307 91699 151373 91700
rect 151494 91357 151554 94691
rect 151632 94210 151692 95200
rect 151768 94757 151828 95200
rect 151904 94890 151964 95200
rect 151904 94830 152106 94890
rect 151765 94756 151831 94757
rect 151765 94692 151766 94756
rect 151830 94692 151831 94756
rect 151765 94691 151831 94692
rect 151632 94150 151738 94210
rect 151491 91356 151557 91357
rect 151491 91292 151492 91356
rect 151556 91292 151557 91356
rect 151491 91291 151557 91292
rect 151678 91221 151738 94150
rect 152046 91221 152106 94830
rect 151675 91220 151741 91221
rect 151675 91156 151676 91220
rect 151740 91156 151741 91220
rect 151675 91155 151741 91156
rect 152043 91220 152109 91221
rect 152043 91156 152044 91220
rect 152108 91156 152109 91220
rect 152043 91155 152109 91156
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 82894 153854 93100
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 86614 157574 93100
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 93100
rect 166214 78573 166274 144875
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 166395 95844 166461 95845
rect 166395 95780 166396 95844
rect 166460 95780 166461 95844
rect 166395 95779 166461 95780
rect 166211 78572 166277 78573
rect 166211 78508 166212 78572
rect 166276 78508 166277 78572
rect 166211 78507 166277 78508
rect 166398 73133 166458 95779
rect 166395 73132 166461 73133
rect 166395 73068 166396 73132
rect 166460 73068 166461 73132
rect 166395 73067 166461 73068
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 169526 38045 169586 271899
rect 170262 112437 170322 337315
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 172467 249252 172533 249253
rect 172467 249188 172468 249252
rect 172532 249188 172533 249252
rect 172467 249187 172533 249188
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 170259 112436 170325 112437
rect 170259 112372 170260 112436
rect 170324 112372 170325 112436
rect 170259 112371 170325 112372
rect 170259 102508 170325 102509
rect 170259 102444 170260 102508
rect 170324 102444 170325 102508
rect 170259 102443 170325 102444
rect 170262 81293 170322 102443
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 170259 81292 170325 81293
rect 170259 81228 170260 81292
rect 170324 81228 170325 81292
rect 170259 81227 170325 81228
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 169523 38044 169589 38045
rect 169523 37980 169524 38044
rect 169588 37980 169589 38044
rect 169523 37979 169589 37980
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 172470 19957 172530 249187
rect 173022 209405 173082 401643
rect 173203 396132 173269 396133
rect 173203 396068 173204 396132
rect 173268 396068 173269 396132
rect 173203 396067 173269 396068
rect 173206 338469 173266 396067
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 173203 338468 173269 338469
rect 173203 338404 173204 338468
rect 173268 338404 173269 338468
rect 173203 338403 173269 338404
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 175782 230213 175842 526355
rect 177803 430676 177869 430677
rect 177803 430612 177804 430676
rect 177868 430612 177869 430676
rect 177803 430611 177869 430612
rect 175779 230212 175845 230213
rect 175779 230148 175780 230212
rect 175844 230148 175845 230212
rect 175779 230147 175845 230148
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 173019 209404 173085 209405
rect 173019 209340 173020 209404
rect 173084 209340 173085 209404
rect 173019 209339 173085 209340
rect 174954 176614 175574 212058
rect 177806 202877 177866 430611
rect 179275 377364 179341 377365
rect 179275 377300 179276 377364
rect 179340 377300 179341 377364
rect 179275 377299 179341 377300
rect 178539 331940 178605 331941
rect 178539 331876 178540 331940
rect 178604 331876 178605 331940
rect 178539 331875 178605 331876
rect 178542 212533 178602 331875
rect 179278 228445 179338 377299
rect 180563 371924 180629 371925
rect 180563 371860 180564 371924
rect 180628 371860 180629 371924
rect 180563 371859 180629 371860
rect 180011 353564 180077 353565
rect 180011 353500 180012 353564
rect 180076 353500 180077 353564
rect 180011 353499 180077 353500
rect 179459 309092 179525 309093
rect 179459 309028 179460 309092
rect 179524 309028 179525 309092
rect 179459 309027 179525 309028
rect 179462 308413 179522 309027
rect 179459 308412 179525 308413
rect 179459 308348 179460 308412
rect 179524 308348 179525 308412
rect 179459 308347 179525 308348
rect 179275 228444 179341 228445
rect 179275 228380 179276 228444
rect 179340 228380 179341 228444
rect 179275 228379 179341 228380
rect 178539 212532 178605 212533
rect 178539 212468 178540 212532
rect 178604 212468 178605 212532
rect 178539 212467 178605 212468
rect 177803 202876 177869 202877
rect 177803 202812 177804 202876
rect 177868 202812 177869 202876
rect 177803 202811 177869 202812
rect 180014 178805 180074 353499
rect 180566 308413 180626 371859
rect 180563 308412 180629 308413
rect 180563 308348 180564 308412
rect 180628 308348 180629 308412
rect 180563 308347 180629 308348
rect 181302 272509 181362 543899
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 184795 449988 184861 449989
rect 184795 449924 184796 449988
rect 184860 449924 184861 449988
rect 184795 449923 184861 449924
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181299 272508 181365 272509
rect 181299 272444 181300 272508
rect 181364 272444 181365 272508
rect 181299 272443 181365 272444
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 184798 225997 184858 449923
rect 185514 439174 186134 474618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 191051 545324 191117 545325
rect 191051 545260 191052 545324
rect 191116 545260 191117 545324
rect 191051 545259 191117 545260
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 187003 447132 187069 447133
rect 187003 447068 187004 447132
rect 187068 447068 187069 447132
rect 187003 447067 187069 447068
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 187006 289781 187066 447067
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 188843 336020 188909 336021
rect 188843 335956 188844 336020
rect 188908 335956 188909 336020
rect 188843 335955 188909 335956
rect 187003 289780 187069 289781
rect 187003 289716 187004 289780
rect 187068 289716 187069 289780
rect 187003 289715 187069 289716
rect 186819 289100 186885 289101
rect 186819 289036 186820 289100
rect 186884 289036 186885 289100
rect 186819 289035 186885 289036
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 184795 225996 184861 225997
rect 184795 225932 184796 225996
rect 184860 225932 184861 225996
rect 184795 225931 184861 225932
rect 184798 225589 184858 225931
rect 184795 225588 184861 225589
rect 184795 225524 184796 225588
rect 184860 225524 184861 225588
rect 184795 225523 184861 225524
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 180011 178804 180077 178805
rect 180011 178740 180012 178804
rect 180076 178740 180077 178804
rect 180011 178739 180077 178740
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 172467 19956 172533 19957
rect 172467 19892 172468 19956
rect 172532 19892 172533 19956
rect 172467 19891 172533 19892
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 186822 64293 186882 289035
rect 188846 234429 188906 335955
rect 189234 334894 189854 370338
rect 190315 363764 190381 363765
rect 190315 363700 190316 363764
rect 190380 363700 190381 363764
rect 190315 363699 190381 363700
rect 190318 363221 190378 363699
rect 190315 363220 190381 363221
rect 190315 363156 190316 363220
rect 190380 363156 190381 363220
rect 190315 363155 190381 363156
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 188843 234428 188909 234429
rect 188843 234364 188844 234428
rect 188908 234364 188909 234428
rect 188843 234363 188909 234364
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 190318 220149 190378 363155
rect 191054 316845 191114 545259
rect 192954 518614 193574 554058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 197859 541244 197925 541245
rect 197859 541180 197860 541244
rect 197924 541180 197925 541244
rect 197859 541179 197925 541180
rect 195099 538524 195165 538525
rect 195099 538460 195100 538524
rect 195164 538460 195165 538524
rect 195099 538459 195165 538460
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192339 386476 192405 386477
rect 192339 386412 192340 386476
rect 192404 386412 192405 386476
rect 192339 386411 192405 386412
rect 191603 326364 191669 326365
rect 191603 326300 191604 326364
rect 191668 326300 191669 326364
rect 191603 326299 191669 326300
rect 191051 316844 191117 316845
rect 191051 316780 191052 316844
rect 191116 316780 191117 316844
rect 191051 316779 191117 316780
rect 191051 289916 191117 289917
rect 191051 289852 191052 289916
rect 191116 289852 191117 289916
rect 191051 289851 191117 289852
rect 191054 271149 191114 289851
rect 191051 271148 191117 271149
rect 191051 271084 191052 271148
rect 191116 271084 191117 271148
rect 191051 271083 191117 271084
rect 191606 258773 191666 326299
rect 192342 295493 192402 386411
rect 192954 374614 193574 410058
rect 194547 381580 194613 381581
rect 194547 381516 194548 381580
rect 194612 381516 194613 381580
rect 194547 381515 194613 381516
rect 194550 375325 194610 381515
rect 194547 375324 194613 375325
rect 194547 375260 194548 375324
rect 194612 375260 194613 375324
rect 194547 375259 194613 375260
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 195102 366349 195162 538459
rect 197862 526421 197922 541179
rect 199794 537993 200414 560898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 200803 545188 200869 545189
rect 200803 545124 200804 545188
rect 200868 545124 200869 545188
rect 200803 545123 200869 545124
rect 199331 535532 199397 535533
rect 199331 535468 199332 535532
rect 199396 535468 199397 535532
rect 199331 535467 199397 535468
rect 199334 527781 199394 535467
rect 199883 535260 199949 535261
rect 199883 535196 199884 535260
rect 199948 535196 199949 535260
rect 199883 535195 199949 535196
rect 199331 527780 199397 527781
rect 199331 527716 199332 527780
rect 199396 527716 199397 527780
rect 199331 527715 199397 527716
rect 197859 526420 197925 526421
rect 197859 526356 197860 526420
rect 197924 526356 197925 526420
rect 197859 526355 197925 526356
rect 198595 512548 198661 512549
rect 198595 512484 198596 512548
rect 198660 512484 198661 512548
rect 198595 512483 198661 512484
rect 196571 438972 196637 438973
rect 196571 438908 196572 438972
rect 196636 438908 196637 438972
rect 196571 438907 196637 438908
rect 195099 366348 195165 366349
rect 195099 366284 195100 366348
rect 195164 366284 195165 366348
rect 195099 366283 195165 366284
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 195099 337380 195165 337381
rect 195099 337316 195100 337380
rect 195164 337316 195165 337380
rect 195099 337315 195165 337316
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192339 295492 192405 295493
rect 192339 295428 192340 295492
rect 192404 295428 192405 295492
rect 192339 295427 192405 295428
rect 192342 285157 192402 295427
rect 192339 285156 192405 285157
rect 192339 285092 192340 285156
rect 192404 285092 192405 285156
rect 192339 285091 192405 285092
rect 192707 284068 192773 284069
rect 192707 284004 192708 284068
rect 192772 284004 192773 284068
rect 192707 284003 192773 284004
rect 192710 282845 192770 284003
rect 191787 282844 191853 282845
rect 191787 282780 191788 282844
rect 191852 282780 191853 282844
rect 191787 282779 191853 282780
rect 192707 282844 192773 282845
rect 192707 282780 192708 282844
rect 192772 282780 192773 282844
rect 192707 282779 192773 282780
rect 191603 258772 191669 258773
rect 191603 258708 191604 258772
rect 191668 258708 191669 258772
rect 191603 258707 191669 258708
rect 191051 255644 191117 255645
rect 191051 255580 191052 255644
rect 191116 255580 191117 255644
rect 191051 255579 191117 255580
rect 191054 244629 191114 255579
rect 191051 244628 191117 244629
rect 191051 244564 191052 244628
rect 191116 244564 191117 244628
rect 191051 244563 191117 244564
rect 191606 233885 191666 258707
rect 191790 245717 191850 282779
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 191787 245716 191853 245717
rect 191787 245652 191788 245716
rect 191852 245652 191853 245716
rect 191787 245651 191853 245652
rect 191787 244628 191853 244629
rect 191787 244564 191788 244628
rect 191852 244564 191853 244628
rect 191787 244563 191853 244564
rect 191790 241637 191850 244563
rect 192339 242180 192405 242181
rect 192339 242116 192340 242180
rect 192404 242116 192405 242180
rect 192339 242115 192405 242116
rect 191787 241636 191853 241637
rect 191787 241572 191788 241636
rect 191852 241572 191853 241636
rect 191787 241571 191853 241572
rect 192342 236877 192402 242115
rect 192339 236876 192405 236877
rect 192339 236812 192340 236876
rect 192404 236812 192405 236876
rect 192339 236811 192405 236812
rect 191603 233884 191669 233885
rect 191603 233820 191604 233884
rect 191668 233820 191669 233884
rect 191603 233819 191669 233820
rect 192954 230614 193574 266058
rect 193811 262852 193877 262853
rect 193811 262788 193812 262852
rect 193876 262788 193877 262852
rect 193811 262787 193877 262788
rect 193814 237149 193874 262787
rect 195102 259453 195162 337315
rect 195835 281620 195901 281621
rect 195835 281556 195836 281620
rect 195900 281556 195901 281620
rect 195835 281555 195901 281556
rect 195099 259452 195165 259453
rect 195099 259388 195100 259452
rect 195164 259388 195165 259452
rect 195099 259387 195165 259388
rect 193811 237148 193877 237149
rect 193811 237084 193812 237148
rect 193876 237084 193877 237148
rect 193811 237083 193877 237084
rect 193811 232660 193877 232661
rect 193811 232596 193812 232660
rect 193876 232596 193877 232660
rect 193811 232595 193877 232596
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 191051 228444 191117 228445
rect 191051 228380 191052 228444
rect 191116 228380 191117 228444
rect 191051 228379 191117 228380
rect 190315 220148 190381 220149
rect 190315 220084 190316 220148
rect 190380 220084 190381 220148
rect 190315 220083 190381 220084
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 188843 185604 188909 185605
rect 188843 185540 188844 185604
rect 188908 185540 188909 185604
rect 188843 185539 188909 185540
rect 186819 64292 186885 64293
rect 186819 64228 186820 64292
rect 186884 64228 186885 64292
rect 186819 64227 186885 64228
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 188846 4997 188906 185539
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 191054 69733 191114 228379
rect 192954 194614 193574 230058
rect 193814 228717 193874 232595
rect 193811 228716 193877 228717
rect 193811 228652 193812 228716
rect 193876 228652 193877 228716
rect 193811 228651 193877 228652
rect 195838 221917 195898 281555
rect 196574 268429 196634 438907
rect 198598 385117 198658 512483
rect 198779 458420 198845 458421
rect 198779 458356 198780 458420
rect 198844 458356 198845 458420
rect 198779 458355 198845 458356
rect 198595 385116 198661 385117
rect 198595 385052 198596 385116
rect 198660 385052 198661 385116
rect 198595 385051 198661 385052
rect 198411 318884 198477 318885
rect 198411 318820 198412 318884
rect 198476 318820 198477 318884
rect 198411 318819 198477 318820
rect 196939 277404 197005 277405
rect 196939 277340 196940 277404
rect 197004 277340 197005 277404
rect 196939 277339 197005 277340
rect 196755 268564 196821 268565
rect 196755 268500 196756 268564
rect 196820 268500 196821 268564
rect 196755 268499 196821 268500
rect 196571 268428 196637 268429
rect 196571 268364 196572 268428
rect 196636 268364 196637 268428
rect 196571 268363 196637 268364
rect 196758 234565 196818 268499
rect 196942 255645 197002 277339
rect 198414 271013 198474 318819
rect 198598 307733 198658 385051
rect 198782 370837 198842 458355
rect 199886 376549 199946 535195
rect 199883 376548 199949 376549
rect 199883 376484 199884 376548
rect 199948 376484 199949 376548
rect 199883 376483 199949 376484
rect 198779 370836 198845 370837
rect 198779 370772 198780 370836
rect 198844 370772 198845 370836
rect 198779 370771 198845 370772
rect 199794 345454 200414 375600
rect 200806 367845 200866 545123
rect 203514 537993 204134 564618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 537993 207854 568338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 537993 211574 572058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 537993 218414 542898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 537993 222134 546618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 537993 225854 550338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 537993 229574 554058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 537993 236414 560898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 537993 240134 564618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 537993 243854 568338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 537993 247574 572058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 537993 254414 542898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 537993 258134 546618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 537993 261854 550338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 537993 265574 554058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 537993 272414 560898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 537993 276134 564618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 537993 279854 568338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 537993 283574 572058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 537993 290414 542898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 537993 294134 546618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 537993 297854 550338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 537993 301574 554058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 537993 308414 560898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 537993 312134 564618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 537993 315854 568338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 537993 319574 572058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 537993 326414 542898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 537993 330134 546618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 537993 333854 550338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 537993 337574 554058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 537993 344414 560898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 537993 348134 564618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 537993 351854 568338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 353339 546684 353405 546685
rect 353339 546620 353340 546684
rect 353404 546620 353405 546684
rect 353339 546619 353405 546620
rect 352051 544100 352117 544101
rect 352051 544036 352052 544100
rect 352116 544036 352117 544100
rect 352051 544035 352117 544036
rect 219568 525454 219888 525486
rect 219568 525218 219610 525454
rect 219846 525218 219888 525454
rect 219568 525134 219888 525218
rect 219568 524898 219610 525134
rect 219846 524898 219888 525134
rect 219568 524866 219888 524898
rect 250288 525454 250608 525486
rect 250288 525218 250330 525454
rect 250566 525218 250608 525454
rect 250288 525134 250608 525218
rect 250288 524898 250330 525134
rect 250566 524898 250608 525134
rect 250288 524866 250608 524898
rect 281008 525454 281328 525486
rect 281008 525218 281050 525454
rect 281286 525218 281328 525454
rect 281008 525134 281328 525218
rect 281008 524898 281050 525134
rect 281286 524898 281328 525134
rect 281008 524866 281328 524898
rect 311728 525454 312048 525486
rect 311728 525218 311770 525454
rect 312006 525218 312048 525454
rect 311728 525134 312048 525218
rect 311728 524898 311770 525134
rect 312006 524898 312048 525134
rect 311728 524866 312048 524898
rect 342448 525454 342768 525486
rect 342448 525218 342490 525454
rect 342726 525218 342768 525454
rect 342448 525134 342768 525218
rect 342448 524898 342490 525134
rect 342726 524898 342768 525134
rect 342448 524866 342768 524898
rect 204208 507454 204528 507486
rect 204208 507218 204250 507454
rect 204486 507218 204528 507454
rect 204208 507134 204528 507218
rect 204208 506898 204250 507134
rect 204486 506898 204528 507134
rect 204208 506866 204528 506898
rect 234928 507454 235248 507486
rect 234928 507218 234970 507454
rect 235206 507218 235248 507454
rect 234928 507134 235248 507218
rect 234928 506898 234970 507134
rect 235206 506898 235248 507134
rect 234928 506866 235248 506898
rect 265648 507454 265968 507486
rect 265648 507218 265690 507454
rect 265926 507218 265968 507454
rect 265648 507134 265968 507218
rect 265648 506898 265690 507134
rect 265926 506898 265968 507134
rect 265648 506866 265968 506898
rect 296368 507454 296688 507486
rect 296368 507218 296410 507454
rect 296646 507218 296688 507454
rect 296368 507134 296688 507218
rect 296368 506898 296410 507134
rect 296646 506898 296688 507134
rect 296368 506866 296688 506898
rect 327088 507454 327408 507486
rect 327088 507218 327130 507454
rect 327366 507218 327408 507454
rect 327088 507134 327408 507218
rect 327088 506898 327130 507134
rect 327366 506898 327408 507134
rect 327088 506866 327408 506898
rect 219568 489454 219888 489486
rect 219568 489218 219610 489454
rect 219846 489218 219888 489454
rect 219568 489134 219888 489218
rect 219568 488898 219610 489134
rect 219846 488898 219888 489134
rect 219568 488866 219888 488898
rect 250288 489454 250608 489486
rect 250288 489218 250330 489454
rect 250566 489218 250608 489454
rect 250288 489134 250608 489218
rect 250288 488898 250330 489134
rect 250566 488898 250608 489134
rect 250288 488866 250608 488898
rect 281008 489454 281328 489486
rect 281008 489218 281050 489454
rect 281286 489218 281328 489454
rect 281008 489134 281328 489218
rect 281008 488898 281050 489134
rect 281286 488898 281328 489134
rect 281008 488866 281328 488898
rect 311728 489454 312048 489486
rect 311728 489218 311770 489454
rect 312006 489218 312048 489454
rect 311728 489134 312048 489218
rect 311728 488898 311770 489134
rect 312006 488898 312048 489134
rect 311728 488866 312048 488898
rect 342448 489454 342768 489486
rect 342448 489218 342490 489454
rect 342726 489218 342768 489454
rect 342448 489134 342768 489218
rect 342448 488898 342490 489134
rect 342726 488898 342768 489134
rect 342448 488866 342768 488898
rect 204208 471454 204528 471486
rect 204208 471218 204250 471454
rect 204486 471218 204528 471454
rect 204208 471134 204528 471218
rect 204208 470898 204250 471134
rect 204486 470898 204528 471134
rect 204208 470866 204528 470898
rect 234928 471454 235248 471486
rect 234928 471218 234970 471454
rect 235206 471218 235248 471454
rect 234928 471134 235248 471218
rect 234928 470898 234970 471134
rect 235206 470898 235248 471134
rect 234928 470866 235248 470898
rect 265648 471454 265968 471486
rect 265648 471218 265690 471454
rect 265926 471218 265968 471454
rect 265648 471134 265968 471218
rect 265648 470898 265690 471134
rect 265926 470898 265968 471134
rect 265648 470866 265968 470898
rect 296368 471454 296688 471486
rect 296368 471218 296410 471454
rect 296646 471218 296688 471454
rect 296368 471134 296688 471218
rect 296368 470898 296410 471134
rect 296646 470898 296688 471134
rect 296368 470866 296688 470898
rect 327088 471454 327408 471486
rect 327088 471218 327130 471454
rect 327366 471218 327408 471454
rect 327088 471134 327408 471218
rect 327088 470898 327130 471134
rect 327366 470898 327408 471134
rect 327088 470866 327408 470898
rect 219568 453454 219888 453486
rect 219568 453218 219610 453454
rect 219846 453218 219888 453454
rect 219568 453134 219888 453218
rect 219568 452898 219610 453134
rect 219846 452898 219888 453134
rect 219568 452866 219888 452898
rect 250288 453454 250608 453486
rect 250288 453218 250330 453454
rect 250566 453218 250608 453454
rect 250288 453134 250608 453218
rect 250288 452898 250330 453134
rect 250566 452898 250608 453134
rect 250288 452866 250608 452898
rect 281008 453454 281328 453486
rect 281008 453218 281050 453454
rect 281286 453218 281328 453454
rect 281008 453134 281328 453218
rect 281008 452898 281050 453134
rect 281286 452898 281328 453134
rect 281008 452866 281328 452898
rect 311728 453454 312048 453486
rect 311728 453218 311770 453454
rect 312006 453218 312048 453454
rect 311728 453134 312048 453218
rect 311728 452898 311770 453134
rect 312006 452898 312048 453134
rect 311728 452866 312048 452898
rect 342448 453454 342768 453486
rect 342448 453218 342490 453454
rect 342726 453218 342768 453454
rect 342448 453134 342768 453218
rect 342448 452898 342490 453134
rect 342726 452898 342768 453134
rect 342448 452866 342768 452898
rect 204208 435454 204528 435486
rect 204208 435218 204250 435454
rect 204486 435218 204528 435454
rect 204208 435134 204528 435218
rect 204208 434898 204250 435134
rect 204486 434898 204528 435134
rect 204208 434866 204528 434898
rect 234928 435454 235248 435486
rect 234928 435218 234970 435454
rect 235206 435218 235248 435454
rect 234928 435134 235248 435218
rect 234928 434898 234970 435134
rect 235206 434898 235248 435134
rect 234928 434866 235248 434898
rect 265648 435454 265968 435486
rect 265648 435218 265690 435454
rect 265926 435218 265968 435454
rect 265648 435134 265968 435218
rect 265648 434898 265690 435134
rect 265926 434898 265968 435134
rect 265648 434866 265968 434898
rect 296368 435454 296688 435486
rect 296368 435218 296410 435454
rect 296646 435218 296688 435454
rect 296368 435134 296688 435218
rect 296368 434898 296410 435134
rect 296646 434898 296688 435134
rect 296368 434866 296688 434898
rect 327088 435454 327408 435486
rect 327088 435218 327130 435454
rect 327366 435218 327408 435454
rect 327088 435134 327408 435218
rect 327088 434898 327130 435134
rect 327366 434898 327408 435134
rect 327088 434866 327408 434898
rect 219568 417454 219888 417486
rect 219568 417218 219610 417454
rect 219846 417218 219888 417454
rect 219568 417134 219888 417218
rect 219568 416898 219610 417134
rect 219846 416898 219888 417134
rect 219568 416866 219888 416898
rect 250288 417454 250608 417486
rect 250288 417218 250330 417454
rect 250566 417218 250608 417454
rect 250288 417134 250608 417218
rect 250288 416898 250330 417134
rect 250566 416898 250608 417134
rect 250288 416866 250608 416898
rect 281008 417454 281328 417486
rect 281008 417218 281050 417454
rect 281286 417218 281328 417454
rect 281008 417134 281328 417218
rect 281008 416898 281050 417134
rect 281286 416898 281328 417134
rect 281008 416866 281328 416898
rect 311728 417454 312048 417486
rect 311728 417218 311770 417454
rect 312006 417218 312048 417454
rect 311728 417134 312048 417218
rect 311728 416898 311770 417134
rect 312006 416898 312048 417134
rect 311728 416866 312048 416898
rect 342448 417454 342768 417486
rect 342448 417218 342490 417454
rect 342726 417218 342768 417454
rect 342448 417134 342768 417218
rect 342448 416898 342490 417134
rect 342726 416898 342768 417134
rect 342448 416866 342768 416898
rect 204208 399454 204528 399486
rect 204208 399218 204250 399454
rect 204486 399218 204528 399454
rect 204208 399134 204528 399218
rect 204208 398898 204250 399134
rect 204486 398898 204528 399134
rect 204208 398866 204528 398898
rect 234928 399454 235248 399486
rect 234928 399218 234970 399454
rect 235206 399218 235248 399454
rect 234928 399134 235248 399218
rect 234928 398898 234970 399134
rect 235206 398898 235248 399134
rect 234928 398866 235248 398898
rect 265648 399454 265968 399486
rect 265648 399218 265690 399454
rect 265926 399218 265968 399454
rect 265648 399134 265968 399218
rect 265648 398898 265690 399134
rect 265926 398898 265968 399134
rect 265648 398866 265968 398898
rect 296368 399454 296688 399486
rect 296368 399218 296410 399454
rect 296646 399218 296688 399454
rect 296368 399134 296688 399218
rect 296368 398898 296410 399134
rect 296646 398898 296688 399134
rect 296368 398866 296688 398898
rect 327088 399454 327408 399486
rect 327088 399218 327130 399454
rect 327366 399218 327408 399454
rect 327088 399134 327408 399218
rect 327088 398898 327130 399134
rect 327366 398898 327408 399134
rect 327088 398866 327408 398898
rect 219568 381454 219888 381486
rect 219568 381218 219610 381454
rect 219846 381218 219888 381454
rect 219568 381134 219888 381218
rect 219568 380898 219610 381134
rect 219846 380898 219888 381134
rect 219568 380866 219888 380898
rect 250288 381454 250608 381486
rect 250288 381218 250330 381454
rect 250566 381218 250608 381454
rect 250288 381134 250608 381218
rect 250288 380898 250330 381134
rect 250566 380898 250608 381134
rect 250288 380866 250608 380898
rect 281008 381454 281328 381486
rect 281008 381218 281050 381454
rect 281286 381218 281328 381454
rect 281008 381134 281328 381218
rect 281008 380898 281050 381134
rect 281286 380898 281328 381134
rect 281008 380866 281328 380898
rect 311728 381454 312048 381486
rect 311728 381218 311770 381454
rect 312006 381218 312048 381454
rect 311728 381134 312048 381218
rect 311728 380898 311770 381134
rect 312006 380898 312048 381134
rect 311728 380866 312048 380898
rect 342448 381454 342768 381486
rect 342448 381218 342490 381454
rect 342726 381218 342768 381454
rect 342448 381134 342768 381218
rect 342448 380898 342490 381134
rect 342726 380898 342768 381134
rect 342448 380866 342768 380898
rect 200803 367844 200869 367845
rect 200803 367780 200804 367844
rect 200868 367780 200869 367844
rect 200803 367779 200869 367780
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 198595 307732 198661 307733
rect 198595 307668 198596 307732
rect 198660 307668 198661 307732
rect 198595 307667 198661 307668
rect 199515 297396 199581 297397
rect 199515 297332 199516 297396
rect 199580 297332 199581 297396
rect 199515 297331 199581 297332
rect 198595 291140 198661 291141
rect 198595 291076 198596 291140
rect 198660 291076 198661 291140
rect 198595 291075 198661 291076
rect 198598 282981 198658 291075
rect 198779 284340 198845 284341
rect 198779 284276 198780 284340
rect 198844 284276 198845 284340
rect 198779 284275 198845 284276
rect 198595 282980 198661 282981
rect 198595 282916 198596 282980
rect 198660 282916 198661 282980
rect 198595 282915 198661 282916
rect 198782 281621 198842 284275
rect 199518 281621 199578 297331
rect 199794 286182 200414 308898
rect 203514 349174 204134 375600
rect 206875 359548 206941 359549
rect 206875 359484 206876 359548
rect 206940 359484 206941 359548
rect 206875 359483 206941 359484
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 200619 291140 200685 291141
rect 200619 291076 200620 291140
rect 200684 291076 200685 291140
rect 200619 291075 200685 291076
rect 200067 283524 200133 283525
rect 200067 283460 200068 283524
rect 200132 283460 200133 283524
rect 200067 283459 200133 283460
rect 200070 283250 200130 283459
rect 199886 283190 200130 283250
rect 198779 281620 198845 281621
rect 198779 281556 198780 281620
rect 198844 281556 198845 281620
rect 198779 281555 198845 281556
rect 199515 281620 199581 281621
rect 199515 281556 199516 281620
rect 199580 281556 199581 281620
rect 199515 281555 199581 281556
rect 199331 281348 199397 281349
rect 199331 281284 199332 281348
rect 199396 281284 199397 281348
rect 199331 281283 199397 281284
rect 198411 271012 198477 271013
rect 198411 270948 198412 271012
rect 198476 270948 198477 271012
rect 198411 270947 198477 270948
rect 197307 264212 197373 264213
rect 197307 264148 197308 264212
rect 197372 264148 197373 264212
rect 197307 264147 197373 264148
rect 197310 263125 197370 264147
rect 197307 263124 197373 263125
rect 197307 263060 197308 263124
rect 197372 263060 197373 263124
rect 197307 263059 197373 263060
rect 196939 255644 197005 255645
rect 196939 255580 196940 255644
rect 197004 255580 197005 255644
rect 196939 255579 197005 255580
rect 199334 249117 199394 281283
rect 199886 277410 199946 283190
rect 200622 281349 200682 291075
rect 203514 286182 204134 312618
rect 204483 311132 204549 311133
rect 204483 311068 204484 311132
rect 204548 311068 204549 311132
rect 204483 311067 204549 311068
rect 204486 285701 204546 311067
rect 204483 285700 204549 285701
rect 204483 285636 204484 285700
rect 204548 285636 204549 285700
rect 204483 285635 204549 285636
rect 205403 283932 205469 283933
rect 205403 283868 205404 283932
rect 205468 283868 205469 283932
rect 205403 283867 205469 283868
rect 200619 281348 200685 281349
rect 200619 281284 200620 281348
rect 200684 281284 200685 281348
rect 200619 281283 200685 281284
rect 199886 277405 200130 277410
rect 199886 277404 200133 277405
rect 199886 277350 200068 277404
rect 200067 277340 200068 277350
rect 200132 277340 200133 277404
rect 200067 277339 200133 277340
rect 204408 255454 204728 255486
rect 204408 255218 204450 255454
rect 204686 255218 204728 255454
rect 204408 255134 204728 255218
rect 204408 254898 204450 255134
rect 204686 254898 204728 255134
rect 204408 254866 204728 254898
rect 199515 252244 199581 252245
rect 199515 252180 199516 252244
rect 199580 252180 199581 252244
rect 199515 252179 199581 252180
rect 199331 249116 199397 249117
rect 199331 249052 199332 249116
rect 199396 249052 199397 249116
rect 199331 249051 199397 249052
rect 199331 244900 199397 244901
rect 199331 244836 199332 244900
rect 199396 244836 199397 244900
rect 199331 244835 199397 244836
rect 196755 234564 196821 234565
rect 196755 234500 196756 234564
rect 196820 234500 196821 234564
rect 196755 234499 196821 234500
rect 199334 223005 199394 244835
rect 199518 237421 199578 252179
rect 200619 244084 200685 244085
rect 200619 244020 200620 244084
rect 200684 244020 200685 244084
rect 200619 244019 200685 244020
rect 199794 237454 200414 238182
rect 199515 237420 199581 237421
rect 199515 237356 199516 237420
rect 199580 237356 199581 237420
rect 199515 237355 199581 237356
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199331 223004 199397 223005
rect 199331 222940 199332 223004
rect 199396 222940 199397 223004
rect 199331 222939 199397 222940
rect 195835 221916 195901 221917
rect 195835 221852 195836 221916
rect 195900 221852 195901 221916
rect 195835 221851 195901 221852
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 191051 69732 191117 69733
rect 191051 69668 191052 69732
rect 191116 69668 191117 69732
rect 191051 69667 191117 69668
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 188843 4996 188909 4997
rect 188843 4932 188844 4996
rect 188908 4932 188909 4996
rect 188843 4931 188909 4932
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 200622 189957 200682 244019
rect 203514 205174 204134 238182
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 200619 189956 200685 189957
rect 200619 189892 200620 189956
rect 200684 189892 200685 189956
rect 200619 189891 200685 189892
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 205406 95165 205466 283867
rect 206878 238645 206938 359483
rect 207234 352894 207854 375600
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 210954 356614 211574 375600
rect 213683 370700 213749 370701
rect 213683 370636 213684 370700
rect 213748 370636 213749 370700
rect 213683 370635 213749 370636
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 209635 351388 209701 351389
rect 209635 351324 209636 351388
rect 209700 351324 209701 351388
rect 209635 351323 209701 351324
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 286182 207854 316338
rect 208163 297532 208229 297533
rect 208163 297468 208164 297532
rect 208228 297468 208229 297532
rect 208163 297467 208229 297468
rect 208166 240141 208226 297467
rect 209638 240141 209698 351323
rect 210739 344452 210805 344453
rect 210739 344388 210740 344452
rect 210804 344388 210805 344452
rect 210739 344387 210805 344388
rect 210742 240141 210802 344387
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 286182 211574 320058
rect 212395 285836 212461 285837
rect 212395 285772 212396 285836
rect 212460 285772 212461 285836
rect 212395 285771 212461 285772
rect 208163 240140 208229 240141
rect 208163 240076 208164 240140
rect 208228 240076 208229 240140
rect 208163 240075 208229 240076
rect 209635 240140 209701 240141
rect 209635 240076 209636 240140
rect 209700 240076 209701 240140
rect 209635 240075 209701 240076
rect 210739 240140 210805 240141
rect 210739 240076 210740 240140
rect 210804 240076 210805 240140
rect 210739 240075 210805 240076
rect 209638 238781 209698 240075
rect 209635 238780 209701 238781
rect 209635 238716 209636 238780
rect 209700 238716 209701 238780
rect 209635 238715 209701 238716
rect 212398 238645 212458 285771
rect 213686 240141 213746 370635
rect 217794 363454 218414 375600
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217547 301612 217613 301613
rect 217547 301548 217548 301612
rect 217612 301548 217613 301612
rect 217547 301547 217613 301548
rect 214603 296036 214669 296037
rect 214603 295972 214604 296036
rect 214668 295972 214669 296036
rect 214603 295971 214669 295972
rect 214419 283932 214485 283933
rect 214419 283868 214420 283932
rect 214484 283868 214485 283932
rect 214419 283867 214485 283868
rect 213683 240140 213749 240141
rect 213683 240076 213684 240140
rect 213748 240076 213749 240140
rect 213683 240075 213749 240076
rect 206875 238644 206941 238645
rect 206875 238580 206876 238644
rect 206940 238580 206941 238644
rect 206875 238579 206941 238580
rect 212395 238644 212461 238645
rect 212395 238580 212396 238644
rect 212460 238580 212461 238644
rect 212395 238579 212461 238580
rect 205587 234700 205653 234701
rect 205587 234636 205588 234700
rect 205652 234636 205653 234700
rect 205587 234635 205653 234636
rect 205590 231573 205650 234635
rect 205587 231572 205653 231573
rect 205587 231508 205588 231572
rect 205652 231508 205653 231572
rect 205587 231507 205653 231508
rect 207234 208894 207854 238182
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 205403 95164 205469 95165
rect 205403 95100 205404 95164
rect 205468 95100 205469 95164
rect 205403 95099 205469 95100
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 212614 211574 238182
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 214422 205733 214482 283867
rect 214606 240141 214666 295971
rect 216075 283932 216141 283933
rect 216075 283868 216076 283932
rect 216140 283868 216141 283932
rect 216075 283867 216141 283868
rect 214603 240140 214669 240141
rect 214603 240076 214604 240140
rect 214668 240076 214669 240140
rect 214603 240075 214669 240076
rect 216078 225045 216138 283867
rect 217550 240141 217610 301547
rect 217794 291454 218414 326898
rect 221514 367174 222134 375600
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 220859 323780 220925 323781
rect 220859 323716 220860 323780
rect 220924 323716 220925 323780
rect 220859 323715 220925 323716
rect 219203 305692 219269 305693
rect 219203 305628 219204 305692
rect 219268 305628 219269 305692
rect 219203 305627 219269 305628
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 286182 218414 290898
rect 218651 285700 218717 285701
rect 218651 285636 218652 285700
rect 218716 285636 218717 285700
rect 218651 285635 218717 285636
rect 217547 240140 217613 240141
rect 217547 240076 217548 240140
rect 217612 240076 217613 240140
rect 217547 240075 217613 240076
rect 216443 237420 216509 237421
rect 216443 237356 216444 237420
rect 216508 237356 216509 237420
rect 216443 237355 216509 237356
rect 216075 225044 216141 225045
rect 216075 224980 216076 225044
rect 216140 224980 216141 225044
rect 216075 224979 216141 224980
rect 214419 205732 214485 205733
rect 214419 205668 214420 205732
rect 214484 205668 214485 205732
rect 214419 205667 214485 205668
rect 216446 205461 216506 237355
rect 217794 219454 218414 238182
rect 218654 237285 218714 285635
rect 219206 240141 219266 305627
rect 219768 273454 220088 273486
rect 219768 273218 219810 273454
rect 220046 273218 220088 273454
rect 219768 273134 220088 273218
rect 219768 272898 219810 273134
rect 220046 272898 220088 273134
rect 219768 272866 220088 272898
rect 220862 240141 220922 323715
rect 221514 295174 222134 330618
rect 225234 370894 225854 375600
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 224171 314124 224237 314125
rect 224171 314060 224172 314124
rect 224236 314060 224237 314124
rect 224171 314059 224237 314060
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 286182 222134 294618
rect 224174 289917 224234 314059
rect 224723 309908 224789 309909
rect 224723 309844 224724 309908
rect 224788 309844 224789 309908
rect 224723 309843 224789 309844
rect 224171 289916 224237 289917
rect 224171 289852 224172 289916
rect 224236 289852 224237 289916
rect 224171 289851 224237 289852
rect 224174 285701 224234 289851
rect 224171 285700 224237 285701
rect 224171 285636 224172 285700
rect 224236 285636 224237 285700
rect 224171 285635 224237 285636
rect 222331 283932 222397 283933
rect 222331 283868 222332 283932
rect 222396 283868 222397 283932
rect 222331 283867 222397 283868
rect 219203 240140 219269 240141
rect 219203 240076 219204 240140
rect 219268 240076 219269 240140
rect 219203 240075 219269 240076
rect 220859 240140 220925 240141
rect 220859 240076 220860 240140
rect 220924 240076 220925 240140
rect 220859 240075 220925 240076
rect 218651 237284 218717 237285
rect 218651 237220 218652 237284
rect 218716 237220 218717 237284
rect 218651 237219 218717 237220
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 216443 205460 216509 205461
rect 216443 205396 216444 205460
rect 216508 205396 216509 205460
rect 216443 205395 216509 205396
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 178000 218414 182898
rect 221514 223174 222134 238182
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 222334 215253 222394 283867
rect 224726 240141 224786 309843
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 286182 225854 298338
rect 228954 374614 229574 375600
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 235794 345454 236414 375600
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 230427 342276 230493 342277
rect 230427 342212 230428 342276
rect 230492 342212 230493 342276
rect 230427 342211 230493 342212
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 226931 288556 226997 288557
rect 226931 288492 226932 288556
rect 226996 288492 226997 288556
rect 226931 288491 226997 288492
rect 226011 283932 226077 283933
rect 226011 283868 226012 283932
rect 226076 283868 226077 283932
rect 226011 283867 226077 283868
rect 226014 240141 226074 283867
rect 224723 240140 224789 240141
rect 224723 240076 224724 240140
rect 224788 240076 224789 240140
rect 224723 240075 224789 240076
rect 226011 240140 226077 240141
rect 226011 240076 226012 240140
rect 226076 240076 226077 240140
rect 226011 240075 226077 240076
rect 223619 237420 223685 237421
rect 223619 237356 223620 237420
rect 223684 237356 223685 237420
rect 223619 237355 223685 237356
rect 222331 215252 222397 215253
rect 222331 215188 222332 215252
rect 222396 215188 222397 215252
rect 222331 215187 222397 215188
rect 223622 211173 223682 237355
rect 225234 226894 225854 238182
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 223619 211172 223685 211173
rect 223619 211108 223620 211172
rect 223684 211108 223685 211172
rect 223619 211107 223685 211108
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 178000 222134 186618
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 178000 225854 190338
rect 226934 176629 226994 288491
rect 228954 286182 229574 302058
rect 228219 285700 228285 285701
rect 228219 285636 228220 285700
rect 228284 285636 228285 285700
rect 228219 285635 228285 285636
rect 227667 185876 227733 185877
rect 227667 185812 227668 185876
rect 227732 185812 227733 185876
rect 227667 185811 227733 185812
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 226931 176628 226997 176629
rect 226931 176564 226932 176628
rect 226996 176564 226997 176628
rect 226931 176563 226997 176564
rect 227670 176493 227730 185811
rect 227667 176492 227733 176493
rect 227667 176428 227668 176492
rect 227732 176428 227733 176492
rect 227667 176427 227733 176428
rect 210954 176294 211574 176378
rect 228222 176357 228282 285635
rect 229691 283932 229757 283933
rect 229691 283868 229692 283932
rect 229756 283868 229757 283932
rect 229691 283867 229757 283868
rect 228954 230614 229574 238182
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 178000 229574 194058
rect 229139 176764 229205 176765
rect 229139 176700 229140 176764
rect 229204 176700 229205 176764
rect 229139 176699 229205 176700
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 228219 176356 228285 176357
rect 228219 176292 228220 176356
rect 228284 176292 228285 176356
rect 228219 176291 228285 176292
rect 210954 140614 211574 176058
rect 221207 165454 221527 165486
rect 221207 165218 221249 165454
rect 221485 165218 221527 165454
rect 221207 165134 221527 165218
rect 221207 164898 221249 165134
rect 221485 164898 221527 165134
rect 221207 164866 221527 164898
rect 224471 165454 224791 165486
rect 224471 165218 224513 165454
rect 224749 165218 224791 165454
rect 224471 165134 224791 165218
rect 224471 164898 224513 165134
rect 224749 164898 224791 165134
rect 224471 164866 224791 164898
rect 229142 163437 229202 176699
rect 229139 163436 229205 163437
rect 229139 163372 229140 163436
rect 229204 163372 229205 163436
rect 229139 163371 229205 163372
rect 215891 151060 215957 151061
rect 215891 150996 215892 151060
rect 215956 150996 215957 151060
rect 215891 150995 215957 150996
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 215894 89725 215954 150995
rect 219575 147454 219895 147486
rect 219575 147218 219617 147454
rect 219853 147218 219895 147454
rect 219575 147134 219895 147218
rect 219575 146898 219617 147134
rect 219853 146898 219895 147134
rect 219575 146866 219895 146898
rect 222839 147454 223159 147486
rect 222839 147218 222881 147454
rect 223117 147218 223159 147454
rect 222839 147134 223159 147218
rect 222839 146898 222881 147134
rect 223117 146898 223159 147134
rect 222839 146866 223159 146898
rect 226103 147454 226423 147486
rect 226103 147218 226145 147454
rect 226381 147218 226423 147454
rect 226103 147134 226423 147218
rect 226103 146898 226145 147134
rect 226381 146898 226423 147134
rect 226103 146866 226423 146898
rect 216811 137460 216877 137461
rect 216811 137396 216812 137460
rect 216876 137396 216877 137460
rect 216811 137395 216877 137396
rect 216814 132510 216874 137395
rect 229694 137325 229754 283867
rect 230430 240141 230490 342211
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 233739 307052 233805 307053
rect 233739 306988 233740 307052
rect 233804 306988 233805 307052
rect 233739 306987 233805 306988
rect 232083 287468 232149 287469
rect 232083 287404 232084 287468
rect 232148 287404 232149 287468
rect 232083 287403 232149 287404
rect 231899 283932 231965 283933
rect 231899 283868 231900 283932
rect 231964 283868 231965 283932
rect 231899 283867 231965 283868
rect 230427 240140 230493 240141
rect 230427 240076 230428 240140
rect 230492 240076 230493 240140
rect 230427 240075 230493 240076
rect 231902 234157 231962 283867
rect 232086 240141 232146 287403
rect 232083 240140 232149 240141
rect 232083 240076 232084 240140
rect 232148 240076 232149 240140
rect 232083 240075 232149 240076
rect 233742 235517 233802 306987
rect 235794 286182 236414 308898
rect 239514 349174 240134 375600
rect 240363 362540 240429 362541
rect 240363 362476 240364 362540
rect 240428 362476 240429 362540
rect 240363 362475 240429 362476
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 237419 303652 237485 303653
rect 237419 303588 237420 303652
rect 237484 303588 237485 303652
rect 237419 303587 237485 303588
rect 236499 285700 236565 285701
rect 236499 285636 236500 285700
rect 236564 285636 236565 285700
rect 236499 285635 236565 285636
rect 236502 283933 236562 285635
rect 236499 283932 236565 283933
rect 236499 283868 236500 283932
rect 236564 283868 236565 283932
rect 236499 283867 236565 283868
rect 235128 255454 235448 255486
rect 235128 255218 235170 255454
rect 235406 255218 235448 255454
rect 235128 255134 235448 255218
rect 235128 254898 235170 255134
rect 235406 254898 235448 255134
rect 235128 254866 235448 254898
rect 235794 237454 236414 238182
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 233739 235516 233805 235517
rect 233739 235452 233740 235516
rect 233804 235452 233805 235516
rect 233739 235451 233805 235452
rect 231899 234156 231965 234157
rect 231899 234092 231900 234156
rect 231964 234092 231965 234156
rect 231899 234091 231965 234092
rect 233003 234156 233069 234157
rect 233003 234092 233004 234156
rect 233068 234092 233069 234156
rect 233003 234091 233069 234092
rect 230427 233204 230493 233205
rect 230427 233140 230428 233204
rect 230492 233140 230493 233204
rect 230427 233139 230493 233140
rect 230430 150653 230490 233139
rect 231899 229804 231965 229805
rect 231899 229740 231900 229804
rect 231964 229740 231965 229804
rect 231899 229739 231965 229740
rect 230611 199476 230677 199477
rect 230611 199412 230612 199476
rect 230676 199412 230677 199476
rect 230611 199411 230677 199412
rect 230427 150652 230493 150653
rect 230427 150588 230428 150652
rect 230492 150588 230493 150652
rect 230427 150587 230493 150588
rect 230614 146301 230674 199411
rect 230611 146300 230677 146301
rect 230611 146236 230612 146300
rect 230676 146236 230677 146300
rect 230611 146235 230677 146236
rect 231902 145349 231962 229739
rect 233006 214845 233066 234091
rect 234659 218652 234725 218653
rect 234659 218588 234660 218652
rect 234724 218588 234725 218652
rect 234659 218587 234725 218588
rect 233187 216068 233253 216069
rect 233187 216004 233188 216068
rect 233252 216004 233253 216068
rect 233187 216003 233253 216004
rect 233003 214844 233069 214845
rect 233003 214780 233004 214844
rect 233068 214780 233069 214844
rect 233003 214779 233069 214780
rect 232083 214436 232149 214437
rect 232083 214372 232084 214436
rect 232148 214372 232149 214436
rect 232083 214371 232149 214372
rect 231899 145348 231965 145349
rect 231899 145284 231900 145348
rect 231964 145284 231965 145348
rect 231899 145283 231965 145284
rect 231715 144124 231781 144125
rect 231715 144060 231716 144124
rect 231780 144060 231781 144124
rect 231715 144059 231781 144060
rect 231718 143037 231778 144059
rect 231715 143036 231781 143037
rect 231715 142972 231716 143036
rect 231780 142972 231781 143036
rect 231715 142971 231781 142972
rect 230979 142900 231045 142901
rect 230979 142836 230980 142900
rect 231044 142836 231045 142900
rect 230979 142835 231045 142836
rect 229691 137324 229757 137325
rect 229691 137260 229692 137324
rect 229756 137260 229757 137324
rect 229691 137259 229757 137260
rect 216814 132450 217242 132510
rect 215891 89724 215957 89725
rect 215891 89660 215892 89724
rect 215956 89660 215957 89724
rect 215891 89659 215957 89660
rect 217182 88229 217242 132450
rect 229691 131476 229757 131477
rect 229691 131412 229692 131476
rect 229756 131412 229757 131476
rect 229691 131411 229757 131412
rect 221207 129454 221527 129486
rect 221207 129218 221249 129454
rect 221485 129218 221527 129454
rect 221207 129134 221527 129218
rect 221207 128898 221249 129134
rect 221485 128898 221527 129134
rect 221207 128866 221527 128898
rect 224471 129454 224791 129486
rect 224471 129218 224513 129454
rect 224749 129218 224791 129454
rect 224471 129134 224791 129218
rect 224471 128898 224513 129134
rect 224749 128898 224791 129134
rect 224471 128866 224791 128898
rect 219575 111454 219895 111486
rect 219575 111218 219617 111454
rect 219853 111218 219895 111454
rect 219575 111134 219895 111218
rect 219575 110898 219617 111134
rect 219853 110898 219895 111134
rect 219575 110866 219895 110898
rect 222839 111454 223159 111486
rect 222839 111218 222881 111454
rect 223117 111218 223159 111454
rect 222839 111134 223159 111218
rect 222839 110898 222881 111134
rect 223117 110898 223159 111134
rect 222839 110866 223159 110898
rect 226103 111454 226423 111486
rect 226103 111218 226145 111454
rect 226381 111218 226423 111454
rect 226103 111134 226423 111218
rect 226103 110898 226145 111134
rect 226381 110898 226423 111134
rect 226103 110866 226423 110898
rect 229139 97068 229205 97069
rect 229139 97004 229140 97068
rect 229204 97004 229205 97068
rect 229139 97003 229205 97004
rect 229142 96930 229202 97003
rect 227670 96870 229202 96930
rect 219203 95980 219269 95981
rect 219203 95916 219204 95980
rect 219268 95916 219269 95980
rect 219203 95915 219269 95916
rect 217179 88228 217245 88229
rect 217179 88164 217180 88228
rect 217244 88164 217245 88228
rect 217179 88163 217245 88164
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 94000
rect 219206 84149 219266 95915
rect 224907 95572 224973 95573
rect 224907 95508 224908 95572
rect 224972 95508 224973 95572
rect 224907 95507 224973 95508
rect 219203 84148 219269 84149
rect 219203 84084 219204 84148
rect 219268 84084 219269 84148
rect 219203 84083 219269 84084
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 94000
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 224910 39269 224970 95507
rect 225234 82894 225854 94000
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 224907 39268 224973 39269
rect 224907 39204 224908 39268
rect 224972 39204 224973 39268
rect 224907 39203 224973 39204
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 227670 4861 227730 96870
rect 229139 96796 229205 96797
rect 229139 96732 229140 96796
rect 229204 96732 229205 96796
rect 229139 96731 229205 96732
rect 229142 96630 229202 96731
rect 228958 96570 229202 96630
rect 228958 95573 229018 96570
rect 228955 95572 229021 95573
rect 228955 95508 228956 95572
rect 229020 95508 229021 95572
rect 228955 95507 229021 95508
rect 228954 86614 229574 94000
rect 229694 93941 229754 131411
rect 230982 125085 231042 142835
rect 231163 142764 231229 142765
rect 231163 142700 231164 142764
rect 231228 142700 231229 142764
rect 231163 142699 231229 142700
rect 231166 135013 231226 142699
rect 232086 142085 232146 214371
rect 233190 165749 233250 216003
rect 233371 178260 233437 178261
rect 233371 178196 233372 178260
rect 233436 178196 233437 178260
rect 233371 178195 233437 178196
rect 233187 165748 233253 165749
rect 233187 165684 233188 165748
rect 233252 165684 233253 165748
rect 233187 165683 233253 165684
rect 232451 145620 232517 145621
rect 232451 145556 232452 145620
rect 232516 145556 232517 145620
rect 232451 145555 232517 145556
rect 232083 142084 232149 142085
rect 232083 142020 232084 142084
rect 232148 142020 232149 142084
rect 232083 142019 232149 142020
rect 231163 135012 231229 135013
rect 231163 134948 231164 135012
rect 231228 134948 231229 135012
rect 231163 134947 231229 134948
rect 230979 125084 231045 125085
rect 230979 125020 230980 125084
rect 231044 125020 231045 125084
rect 230979 125019 231045 125020
rect 230979 116244 231045 116245
rect 230979 116180 230980 116244
rect 231044 116180 231045 116244
rect 230979 116179 231045 116180
rect 229691 93940 229757 93941
rect 229691 93876 229692 93940
rect 229756 93876 229757 93940
rect 229691 93875 229757 93876
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 227667 4860 227733 4861
rect 227667 4796 227668 4860
rect 227732 4796 227733 4860
rect 227667 4795 227733 4796
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 230982 11661 231042 116179
rect 232454 104277 232514 145555
rect 233374 139229 233434 178195
rect 234662 149701 234722 218587
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 236502 166837 236562 283867
rect 237422 240141 237482 303587
rect 238523 289236 238589 289237
rect 238523 289172 238524 289236
rect 238588 289172 238589 289236
rect 238523 289171 238589 289172
rect 237419 240140 237485 240141
rect 237419 240076 237420 240140
rect 237484 240076 237485 240140
rect 237419 240075 237485 240076
rect 237419 185740 237485 185741
rect 237419 185676 237420 185740
rect 237484 185676 237485 185740
rect 237419 185675 237485 185676
rect 236499 166836 236565 166837
rect 236499 166772 236500 166836
rect 236564 166772 236565 166836
rect 236499 166771 236565 166772
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 234659 149700 234725 149701
rect 234659 149636 234660 149700
rect 234724 149636 234725 149700
rect 234659 149635 234725 149636
rect 233371 139228 233437 139229
rect 233371 139164 233372 139228
rect 233436 139164 233437 139228
rect 233371 139163 233437 139164
rect 233739 135828 233805 135829
rect 233739 135764 233740 135828
rect 233804 135764 233805 135828
rect 233739 135763 233805 135764
rect 232451 104276 232517 104277
rect 232451 104212 232452 104276
rect 232516 104212 232517 104276
rect 232451 104211 232517 104212
rect 233742 51781 233802 135763
rect 235794 129454 236414 164898
rect 237422 148341 237482 185675
rect 237603 181660 237669 181661
rect 237603 181596 237604 181660
rect 237668 181596 237669 181660
rect 237603 181595 237669 181596
rect 237606 156229 237666 181595
rect 237603 156228 237669 156229
rect 237603 156164 237604 156228
rect 237668 156164 237669 156228
rect 237603 156163 237669 156164
rect 238526 154461 238586 289171
rect 239514 286182 240134 312618
rect 239514 205174 240134 238182
rect 240366 207637 240426 362475
rect 243234 352894 243854 375600
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 241651 333436 241717 333437
rect 241651 333372 241652 333436
rect 241716 333372 241717 333436
rect 241651 333371 241717 333372
rect 241654 240141 241714 333371
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 242939 315076 243005 315077
rect 242939 315012 242940 315076
rect 243004 315012 243005 315076
rect 242939 315011 243005 315012
rect 242942 282570 243002 315011
rect 243234 286182 243854 316338
rect 246954 356614 247574 375600
rect 250299 370564 250365 370565
rect 250299 370500 250300 370564
rect 250364 370500 250365 370564
rect 250299 370499 250365 370500
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 247723 323780 247789 323781
rect 247723 323716 247724 323780
rect 247788 323716 247789 323780
rect 247723 323715 247789 323716
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 244411 298348 244477 298349
rect 244411 298284 244412 298348
rect 244476 298284 244477 298348
rect 244411 298283 244477 298284
rect 243675 285972 243741 285973
rect 243675 285908 243676 285972
rect 243740 285908 243741 285972
rect 243675 285907 243741 285908
rect 242942 282510 243554 282570
rect 243494 281349 243554 282510
rect 243491 281348 243557 281349
rect 243491 281284 243492 281348
rect 243556 281284 243557 281348
rect 243491 281283 243557 281284
rect 243678 277410 243738 285907
rect 243126 277350 243738 277410
rect 243126 267750 243186 277350
rect 243126 267690 243554 267750
rect 243494 254149 243554 267690
rect 244227 262580 244293 262581
rect 244227 262516 244228 262580
rect 244292 262516 244293 262580
rect 244227 262515 244293 262516
rect 243491 254148 243557 254149
rect 243491 254084 243492 254148
rect 243556 254084 243557 254148
rect 243491 254083 243557 254084
rect 244043 251972 244109 251973
rect 244043 251908 244044 251972
rect 244108 251908 244109 251972
rect 244043 251907 244109 251908
rect 243491 250068 243557 250069
rect 243491 250004 243492 250068
rect 243556 250004 243557 250068
rect 243491 250003 243557 250004
rect 243494 248430 243554 250003
rect 243310 248370 243554 248430
rect 241651 240140 241717 240141
rect 241651 240076 241652 240140
rect 241716 240076 241717 240140
rect 241651 240075 241717 240076
rect 240363 207636 240429 207637
rect 240363 207572 240364 207636
rect 240428 207572 240429 207636
rect 240363 207571 240429 207572
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 169174 240134 204618
rect 240731 198116 240797 198117
rect 240731 198052 240732 198116
rect 240796 198052 240797 198116
rect 240731 198051 240797 198052
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 238523 154460 238589 154461
rect 238523 154396 238524 154460
rect 238588 154396 238589 154460
rect 238523 154395 238589 154396
rect 237419 148340 237485 148341
rect 237419 148276 237420 148340
rect 237484 148276 237485 148340
rect 237419 148275 237485 148276
rect 236499 146980 236565 146981
rect 236499 146916 236500 146980
rect 236564 146916 236565 146980
rect 236499 146915 236565 146916
rect 236502 141133 236562 146915
rect 237971 141404 238037 141405
rect 237971 141340 237972 141404
rect 238036 141340 238037 141404
rect 237971 141339 238037 141340
rect 236499 141132 236565 141133
rect 236499 141068 236500 141132
rect 236564 141068 236565 141132
rect 236499 141067 236565 141068
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 237974 102237 238034 141339
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 237971 102236 238037 102237
rect 237971 102172 237972 102236
rect 238036 102172 238037 102236
rect 237971 102171 238037 102172
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 233739 51780 233805 51781
rect 233739 51716 233740 51780
rect 233804 51716 233805 51780
rect 233739 51715 233805 51716
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 230979 11660 231045 11661
rect 230979 11596 230980 11660
rect 231044 11596 231045 11660
rect 230979 11595 231045 11596
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 240734 3909 240794 198051
rect 241654 168469 241714 240075
rect 243310 240005 243370 248370
rect 243307 240004 243373 240005
rect 243307 239940 243308 240004
rect 243372 239940 243373 240004
rect 243307 239939 243373 239940
rect 242019 237420 242085 237421
rect 242019 237356 242020 237420
rect 242084 237356 242085 237420
rect 242019 237355 242085 237356
rect 241651 168468 241717 168469
rect 241651 168404 241652 168468
rect 241716 168404 241717 168468
rect 241651 168403 241717 168404
rect 242022 142901 242082 237355
rect 243234 208894 243854 238182
rect 244046 238101 244106 251907
rect 244043 238100 244109 238101
rect 244043 238036 244044 238100
rect 244108 238036 244109 238100
rect 244043 238035 244109 238036
rect 244230 228445 244290 262515
rect 244414 259589 244474 298283
rect 246803 291820 246869 291821
rect 246803 291756 246804 291820
rect 246868 291756 246869 291820
rect 246803 291755 246869 291756
rect 246251 290052 246317 290053
rect 246251 289988 246252 290052
rect 246316 289988 246317 290052
rect 246251 289987 246317 289988
rect 244595 284476 244661 284477
rect 244595 284412 244596 284476
rect 244660 284412 244661 284476
rect 244595 284411 244661 284412
rect 244598 283661 244658 284411
rect 244595 283660 244661 283661
rect 244595 283596 244596 283660
rect 244660 283596 244661 283660
rect 244595 283595 244661 283596
rect 246254 280261 246314 289987
rect 246251 280260 246317 280261
rect 246251 280196 246252 280260
rect 246316 280196 246317 280260
rect 246251 280195 246317 280196
rect 246806 277410 246866 291755
rect 246622 277350 246866 277410
rect 246954 284614 247574 320058
rect 247726 285157 247786 323715
rect 247723 285156 247789 285157
rect 247723 285092 247724 285156
rect 247788 285092 247789 285156
rect 247723 285091 247789 285092
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 246622 267477 246682 277350
rect 246803 268020 246869 268021
rect 246803 267956 246804 268020
rect 246868 267956 246869 268020
rect 246803 267955 246869 267956
rect 246619 267476 246685 267477
rect 246619 267412 246620 267476
rect 246684 267412 246685 267476
rect 246619 267411 246685 267412
rect 246622 267069 246682 267411
rect 246619 267068 246685 267069
rect 246619 267004 246620 267068
rect 246684 267004 246685 267068
rect 246619 267003 246685 267004
rect 246806 263533 246866 267955
rect 246803 263532 246869 263533
rect 246803 263468 246804 263532
rect 246868 263468 246869 263532
rect 246803 263467 246869 263468
rect 244411 259588 244477 259589
rect 244411 259524 244412 259588
rect 244476 259524 244477 259588
rect 244411 259523 244477 259524
rect 246954 248614 247574 284058
rect 248459 273188 248525 273189
rect 248459 273124 248460 273188
rect 248524 273124 248525 273188
rect 248459 273123 248525 273124
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 245699 246532 245765 246533
rect 245699 246468 245700 246532
rect 245764 246468 245765 246532
rect 245699 246467 245765 246468
rect 245702 245717 245762 246467
rect 245699 245716 245765 245717
rect 245699 245652 245700 245716
rect 245764 245652 245765 245716
rect 245699 245651 245765 245652
rect 244227 228444 244293 228445
rect 244227 228380 244228 228444
rect 244292 228380 244293 228444
rect 244227 228379 244293 228380
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 172894 243854 208338
rect 244227 198796 244293 198797
rect 244227 198732 244228 198796
rect 244292 198732 244293 198796
rect 244227 198731 244293 198732
rect 244230 192541 244290 198731
rect 245702 195941 245762 245651
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 245699 195940 245765 195941
rect 245699 195876 245700 195940
rect 245764 195876 245765 195940
rect 245699 195875 245765 195876
rect 244227 192540 244293 192541
rect 244227 192476 244228 192540
rect 244292 192476 244293 192540
rect 244227 192475 244293 192476
rect 245699 191180 245765 191181
rect 245699 191116 245700 191180
rect 245764 191116 245765 191180
rect 245699 191115 245765 191116
rect 244227 175812 244293 175813
rect 244227 175748 244228 175812
rect 244292 175748 244293 175812
rect 244227 175747 244293 175748
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 242019 142900 242085 142901
rect 242019 142836 242020 142900
rect 242084 142836 242085 142900
rect 242019 142835 242085 142836
rect 242019 140180 242085 140181
rect 242019 140116 242020 140180
rect 242084 140116 242085 140180
rect 242019 140115 242085 140116
rect 242022 36549 242082 140115
rect 243234 136894 243854 172338
rect 244230 152557 244290 175747
rect 244227 152556 244293 152557
rect 244227 152492 244228 152556
rect 244292 152492 244293 152556
rect 244227 152491 244293 152492
rect 244227 142492 244293 142493
rect 244227 142428 244228 142492
rect 244292 142428 244293 142492
rect 244227 142427 244293 142428
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 244230 100741 244290 142427
rect 245702 137869 245762 191115
rect 246954 176614 247574 212058
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 248462 160717 248522 273123
rect 250302 270469 250362 370499
rect 253794 363454 254414 375600
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 252507 330580 252573 330581
rect 252507 330516 252508 330580
rect 252572 330516 252573 330580
rect 252507 330515 252573 330516
rect 251219 308684 251285 308685
rect 251219 308620 251220 308684
rect 251284 308620 251285 308684
rect 251219 308619 251285 308620
rect 251222 273053 251282 308619
rect 252510 275773 252570 330515
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 257514 367174 258134 375600
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 255267 294132 255333 294133
rect 255267 294068 255268 294132
rect 255332 294068 255333 294132
rect 255267 294067 255333 294068
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 252507 275772 252573 275773
rect 252507 275708 252508 275772
rect 252572 275708 252573 275772
rect 252507 275707 252573 275708
rect 251219 273052 251285 273053
rect 251219 272988 251220 273052
rect 251284 272988 251285 273052
rect 251219 272987 251285 272988
rect 250299 270468 250365 270469
rect 250299 270404 250300 270468
rect 250364 270404 250365 270468
rect 250299 270403 250365 270404
rect 249747 260948 249813 260949
rect 249747 260884 249748 260948
rect 249812 260884 249813 260948
rect 249747 260883 249813 260884
rect 249011 161804 249077 161805
rect 249011 161740 249012 161804
rect 249076 161740 249077 161804
rect 249011 161739 249077 161740
rect 248459 160716 248525 160717
rect 248459 160652 248460 160716
rect 248524 160652 248525 160716
rect 248459 160651 248525 160652
rect 249014 143037 249074 161739
rect 249750 144805 249810 260883
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253059 217292 253125 217293
rect 253059 217228 253060 217292
rect 253124 217228 253125 217292
rect 253059 217227 253125 217228
rect 249931 185468 249997 185469
rect 249931 185404 249932 185468
rect 249996 185404 249997 185468
rect 249931 185403 249997 185404
rect 249934 153917 249994 185403
rect 249931 153916 249997 153917
rect 249931 153852 249932 153916
rect 249996 153852 249997 153916
rect 249931 153851 249997 153852
rect 249747 144804 249813 144805
rect 249747 144740 249748 144804
rect 249812 144740 249813 144804
rect 249747 144739 249813 144740
rect 249011 143036 249077 143037
rect 249011 142972 249012 143036
rect 249076 142972 249077 143036
rect 249011 142971 249077 142972
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 245699 137868 245765 137869
rect 245699 137804 245700 137868
rect 245764 137804 245765 137868
rect 245699 137803 245765 137804
rect 246251 116108 246317 116109
rect 246251 116044 246252 116108
rect 246316 116044 246317 116108
rect 246251 116043 246317 116044
rect 244227 100740 244293 100741
rect 244227 100676 244228 100740
rect 244292 100676 244293 100740
rect 244227 100675 244293 100676
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 242019 36548 242085 36549
rect 242019 36484 242020 36548
rect 242084 36484 242085 36548
rect 242019 36483 242085 36484
rect 243234 28894 243854 64338
rect 246254 39405 246314 116043
rect 246954 104614 247574 140058
rect 249195 134468 249261 134469
rect 249195 134404 249196 134468
rect 249260 134404 249261 134468
rect 249195 134403 249261 134404
rect 249011 130116 249077 130117
rect 249011 130052 249012 130116
rect 249076 130052 249077 130116
rect 249011 130051 249077 130052
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246251 39404 246317 39405
rect 246251 39340 246252 39404
rect 246316 39340 246317 39404
rect 246251 39339 246317 39340
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 240731 3908 240797 3909
rect 240731 3844 240732 3908
rect 240796 3844 240797 3908
rect 240731 3843 240797 3844
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 68058
rect 249014 43485 249074 130051
rect 249198 90405 249258 134403
rect 249195 90404 249261 90405
rect 249195 90340 249196 90404
rect 249260 90340 249261 90404
rect 249195 90339 249261 90340
rect 249011 43484 249077 43485
rect 249011 43420 249012 43484
rect 249076 43420 249077 43484
rect 249011 43419 249077 43420
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253062 19413 253122 217227
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 255270 96525 255330 294067
rect 257514 259174 258134 294618
rect 261234 370894 261854 375600
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 260051 269244 260117 269245
rect 260051 269180 260052 269244
rect 260116 269180 260117 269244
rect 260051 269179 260117 269180
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 258579 132700 258645 132701
rect 258579 132636 258580 132700
rect 258644 132636 258645 132700
rect 258579 132635 258645 132636
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 255267 96524 255333 96525
rect 255267 96460 255268 96524
rect 255332 96460 255333 96524
rect 255267 96459 255333 96460
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253059 19412 253125 19413
rect 253059 19348 253060 19412
rect 253124 19348 253125 19412
rect 253059 19347 253125 19348
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 258582 44845 258642 132635
rect 258763 102372 258829 102373
rect 258763 102308 258764 102372
rect 258828 102308 258829 102372
rect 258763 102307 258829 102308
rect 258766 93125 258826 102307
rect 260054 95029 260114 269179
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 264954 374614 265574 375600
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 268331 353972 268397 353973
rect 268331 353908 268332 353972
rect 268396 353908 268397 353972
rect 268331 353907 268397 353908
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264099 149020 264165 149021
rect 264099 148956 264100 149020
rect 264164 148956 264165 149020
rect 264099 148955 264165 148956
rect 262811 127124 262877 127125
rect 262811 127060 262812 127124
rect 262876 127060 262877 127124
rect 262811 127059 262877 127060
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 260235 100196 260301 100197
rect 260235 100132 260236 100196
rect 260300 100132 260301 100196
rect 260235 100131 260301 100132
rect 260051 95028 260117 95029
rect 260051 94964 260052 95028
rect 260116 94964 260117 95028
rect 260051 94963 260117 94964
rect 258763 93124 258829 93125
rect 258763 93060 258764 93124
rect 258828 93060 258829 93124
rect 258763 93059 258829 93060
rect 260238 53141 260298 100131
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 260235 53140 260301 53141
rect 260235 53076 260236 53140
rect 260300 53076 260301 53140
rect 260235 53075 260301 53076
rect 261234 46894 261854 82338
rect 262814 76533 262874 127059
rect 264102 107541 264162 148955
rect 264954 122614 265574 158058
rect 267595 128484 267661 128485
rect 267595 128420 267596 128484
rect 267660 128420 267661 128484
rect 267595 128419 267661 128420
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264099 107540 264165 107541
rect 264099 107476 264100 107540
rect 264164 107476 264165 107540
rect 264099 107475 264165 107476
rect 264099 101828 264165 101829
rect 264099 101764 264100 101828
rect 264164 101764 264165 101828
rect 264099 101763 264165 101764
rect 264102 83469 264162 101763
rect 264954 86614 265574 122058
rect 266859 113388 266925 113389
rect 266859 113324 266860 113388
rect 266924 113324 266925 113388
rect 266859 113323 266925 113324
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264099 83468 264165 83469
rect 264099 83404 264100 83468
rect 264164 83404 264165 83468
rect 264099 83403 264165 83404
rect 262811 76532 262877 76533
rect 262811 76468 262812 76532
rect 262876 76468 262877 76532
rect 262811 76467 262877 76468
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 258579 44844 258645 44845
rect 258579 44780 258580 44844
rect 258644 44780 258645 44844
rect 258579 44779 258645 44780
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 86058
rect 266862 77893 266922 113323
rect 267598 94485 267658 128419
rect 267779 113796 267845 113797
rect 267779 113732 267780 113796
rect 267844 113732 267845 113796
rect 267779 113731 267845 113732
rect 267595 94484 267661 94485
rect 267595 94420 267596 94484
rect 267660 94420 267661 94484
rect 267595 94419 267661 94420
rect 266859 77892 266925 77893
rect 266859 77828 266860 77892
rect 266924 77828 266925 77892
rect 266859 77827 266925 77828
rect 267782 62797 267842 113731
rect 267779 62796 267845 62797
rect 267779 62732 267780 62796
rect 267844 62732 267845 62796
rect 267779 62731 267845 62732
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 268334 3501 268394 353907
rect 271794 345454 272414 375600
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 178000 272414 200898
rect 275514 349174 276134 375600
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 178000 276134 204618
rect 279234 352894 279854 375600
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 282954 356614 283574 375600
rect 288755 375324 288821 375325
rect 288755 375260 288756 375324
rect 288820 375260 288821 375324
rect 288755 375259 288821 375260
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 286179 349892 286245 349893
rect 286179 349828 286180 349892
rect 286244 349828 286245 349892
rect 286179 349827 286245 349828
rect 286182 344317 286242 349827
rect 286179 344316 286245 344317
rect 286179 344252 286180 344316
rect 286244 344252 286245 344316
rect 286179 344251 286245 344252
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 281579 320244 281645 320245
rect 281579 320180 281580 320244
rect 281644 320180 281645 320244
rect 281579 320179 281645 320180
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 280291 284068 280357 284069
rect 280291 284004 280292 284068
rect 280356 284004 280357 284068
rect 280291 284003 280357 284004
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279003 195396 279069 195397
rect 279003 195332 279004 195396
rect 279068 195332 279069 195396
rect 279003 195331 279069 195332
rect 277163 186420 277229 186421
rect 277163 186356 277164 186420
rect 277228 186356 277229 186420
rect 277163 186355 277229 186356
rect 277166 176670 277226 186355
rect 278819 178124 278885 178125
rect 278819 178060 278820 178124
rect 278884 178060 278885 178124
rect 278819 178059 278885 178060
rect 277166 176610 277410 176670
rect 277350 175813 277410 176610
rect 277347 175812 277413 175813
rect 277347 175748 277348 175812
rect 277412 175748 277413 175812
rect 277347 175747 277413 175748
rect 272207 165454 272527 165486
rect 272207 165218 272249 165454
rect 272485 165218 272527 165454
rect 272207 165134 272527 165218
rect 272207 164898 272249 165134
rect 272485 164898 272527 165134
rect 272207 164866 272527 164898
rect 275471 165454 275791 165486
rect 275471 165218 275513 165454
rect 275749 165218 275791 165454
rect 275471 165134 275791 165218
rect 275471 164898 275513 165134
rect 275749 164898 275791 165134
rect 275471 164866 275791 164898
rect 270575 147454 270895 147486
rect 270575 147218 270617 147454
rect 270853 147218 270895 147454
rect 270575 147134 270895 147218
rect 270575 146898 270617 147134
rect 270853 146898 270895 147134
rect 270575 146866 270895 146898
rect 273839 147454 274159 147486
rect 273839 147218 273881 147454
rect 274117 147218 274159 147454
rect 273839 147134 274159 147218
rect 273839 146898 273881 147134
rect 274117 146898 274159 147134
rect 273839 146866 274159 146898
rect 277103 147454 277423 147486
rect 277103 147218 277145 147454
rect 277381 147218 277423 147454
rect 277103 147134 277423 147218
rect 277103 146898 277145 147134
rect 277381 146898 277423 147134
rect 277103 146866 277423 146898
rect 272207 129454 272527 129486
rect 272207 129218 272249 129454
rect 272485 129218 272527 129454
rect 272207 129134 272527 129218
rect 272207 128898 272249 129134
rect 272485 128898 272527 129134
rect 272207 128866 272527 128898
rect 275471 129454 275791 129486
rect 275471 129218 275513 129454
rect 275749 129218 275791 129454
rect 275471 129134 275791 129218
rect 275471 128898 275513 129134
rect 275749 128898 275791 129134
rect 275471 128866 275791 128898
rect 278822 113190 278882 178059
rect 279006 176670 279066 195331
rect 279234 178000 279854 208338
rect 279006 176610 279434 176670
rect 279374 167653 279434 176610
rect 280294 172549 280354 284003
rect 280475 178124 280541 178125
rect 280475 178060 280476 178124
rect 280540 178060 280541 178124
rect 280475 178059 280541 178060
rect 280291 172548 280357 172549
rect 280291 172484 280292 172548
rect 280356 172484 280357 172548
rect 280291 172483 280357 172484
rect 280478 167925 280538 178059
rect 280475 167924 280541 167925
rect 280475 167860 280476 167924
rect 280540 167860 280541 167924
rect 280475 167859 280541 167860
rect 279371 167652 279437 167653
rect 279371 167588 279372 167652
rect 279436 167588 279437 167652
rect 279371 167587 279437 167588
rect 281582 156501 281642 320179
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 283787 286380 283853 286381
rect 283787 286316 283788 286380
rect 283852 286316 283853 286380
rect 283787 286315 283853 286316
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 281763 185740 281829 185741
rect 281763 185676 281764 185740
rect 281828 185676 281829 185740
rect 281763 185675 281829 185676
rect 281766 163301 281826 185675
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 281763 163300 281829 163301
rect 281763 163236 281764 163300
rect 281828 163236 281829 163300
rect 281763 163235 281829 163236
rect 281579 156500 281645 156501
rect 281579 156436 281580 156500
rect 281644 156436 281645 156500
rect 281579 156435 281645 156436
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 278822 113130 279434 113190
rect 270575 111454 270895 111486
rect 270575 111218 270617 111454
rect 270853 111218 270895 111454
rect 270575 111134 270895 111218
rect 270575 110898 270617 111134
rect 270853 110898 270895 111134
rect 270575 110866 270895 110898
rect 273839 111454 274159 111486
rect 273839 111218 273881 111454
rect 274117 111218 274159 111454
rect 273839 111134 274159 111218
rect 273839 110898 273881 111134
rect 274117 110898 274159 111134
rect 273839 110866 274159 110898
rect 277103 111454 277423 111486
rect 277103 111218 277145 111454
rect 277381 111218 277423 111454
rect 277103 111134 277423 111218
rect 277103 110898 277145 111134
rect 277381 110898 277423 111134
rect 277103 110866 277423 110898
rect 279374 99517 279434 113130
rect 282131 109172 282197 109173
rect 282131 109108 282132 109172
rect 282196 109108 282197 109172
rect 282131 109107 282197 109108
rect 279371 99516 279437 99517
rect 279371 99452 279372 99516
rect 279436 99452 279437 99516
rect 279371 99451 279437 99452
rect 271794 93454 272414 94000
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 268331 3500 268397 3501
rect 268331 3436 268332 3500
rect 268396 3436 268397 3500
rect 268331 3435 268397 3436
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 61174 276134 94000
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 64894 279854 94000
rect 282134 88229 282194 109107
rect 282954 104614 283574 140058
rect 283790 109989 283850 286315
rect 284339 194580 284405 194581
rect 284339 194516 284340 194580
rect 284404 194516 284405 194580
rect 284339 194515 284405 194516
rect 284342 135149 284402 194515
rect 285627 186420 285693 186421
rect 285627 186356 285628 186420
rect 285692 186356 285693 186420
rect 285627 186355 285693 186356
rect 284523 177988 284589 177989
rect 284523 177924 284524 177988
rect 284588 177924 284589 177988
rect 284523 177923 284589 177924
rect 284339 135148 284405 135149
rect 284339 135084 284340 135148
rect 284404 135084 284405 135148
rect 284339 135083 284405 135084
rect 284526 134469 284586 177923
rect 284523 134468 284589 134469
rect 284523 134404 284524 134468
rect 284588 134404 284589 134468
rect 284523 134403 284589 134404
rect 285630 133653 285690 186355
rect 285627 133652 285693 133653
rect 285627 133588 285628 133652
rect 285692 133588 285693 133652
rect 285627 133587 285693 133588
rect 283787 109988 283853 109989
rect 283787 109924 283788 109988
rect 283852 109924 283853 109988
rect 283787 109923 283853 109924
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282131 88228 282197 88229
rect 282131 88164 282132 88228
rect 282196 88164 282197 88228
rect 282131 88163 282197 88164
rect 282134 84210 282194 88163
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 281582 84150 282194 84210
rect 281582 29613 281642 84150
rect 282954 68614 283574 104058
rect 286182 93125 286242 344251
rect 287099 293996 287165 293997
rect 287099 293932 287100 293996
rect 287164 293932 287165 293996
rect 287099 293931 287165 293932
rect 287102 101013 287162 293931
rect 287651 191044 287717 191045
rect 287651 190980 287652 191044
rect 287716 190980 287717 191044
rect 287651 190979 287717 190980
rect 287654 190470 287714 190979
rect 288758 190470 288818 375259
rect 287654 190410 288818 190470
rect 289794 363454 290414 375600
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 293514 367174 294134 375600
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 291699 344452 291765 344453
rect 291699 344388 291700 344452
rect 291764 344388 291765 344452
rect 291699 344387 291765 344388
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 287099 101012 287165 101013
rect 287099 100948 287100 101012
rect 287164 100948 287165 101012
rect 287099 100947 287165 100948
rect 286179 93124 286245 93125
rect 286179 93060 286180 93124
rect 286244 93060 286245 93124
rect 286179 93059 286245 93060
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 281579 29612 281645 29613
rect 281579 29548 281580 29612
rect 281644 29548 281645 29612
rect 281579 29547 281645 29548
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 287654 21453 287714 190410
rect 289794 183454 290414 218898
rect 291147 192676 291213 192677
rect 291147 192612 291148 192676
rect 291212 192612 291213 192676
rect 291147 192611 291213 192612
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 288571 183156 288637 183157
rect 288571 183092 288572 183156
rect 288636 183092 288637 183156
rect 288571 183091 288637 183092
rect 289794 183134 290414 183218
rect 287651 21452 287717 21453
rect 287651 21388 287652 21452
rect 287716 21388 287717 21452
rect 287651 21387 287717 21388
rect 288574 8261 288634 183091
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 290595 180164 290661 180165
rect 290595 180100 290596 180164
rect 290660 180100 290661 180164
rect 290595 180099 290661 180100
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 290598 102237 290658 180099
rect 290595 102236 290661 102237
rect 290595 102172 290596 102236
rect 290660 102172 290661 102236
rect 290595 102171 290661 102172
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 291150 66197 291210 192611
rect 291702 97885 291762 344387
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 297234 370894 297854 375600
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 295931 202332 295997 202333
rect 295931 202268 295932 202332
rect 295996 202268 295997 202332
rect 295931 202267 295997 202268
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 295934 149157 295994 202267
rect 297234 190894 297854 226338
rect 300954 374614 301574 375600
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 307794 345454 308414 375600
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 304211 302292 304277 302293
rect 304211 302228 304212 302292
rect 304276 302228 304277 302292
rect 304211 302227 304277 302228
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 302739 240820 302805 240821
rect 302739 240756 302740 240820
rect 302804 240756 302805 240820
rect 302739 240755 302805 240756
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 298139 225588 298205 225589
rect 298139 225524 298140 225588
rect 298204 225524 298205 225588
rect 298139 225523 298205 225524
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 295931 149156 295997 149157
rect 295931 149092 295932 149156
rect 295996 149092 295997 149156
rect 295931 149091 295997 149092
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 291699 97884 291765 97885
rect 291699 97820 291700 97884
rect 291764 97820 291765 97884
rect 291699 97819 291765 97820
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 291147 66196 291213 66197
rect 291147 66132 291148 66196
rect 291212 66132 291213 66196
rect 291147 66131 291213 66132
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 288755 21452 288821 21453
rect 288755 21388 288756 21452
rect 288820 21388 288821 21452
rect 288755 21387 288821 21388
rect 288758 12205 288818 21387
rect 288755 12204 288821 12205
rect 288755 12140 288756 12204
rect 288820 12140 288821 12204
rect 288755 12139 288821 12140
rect 288571 8260 288637 8261
rect 288571 8196 288572 8260
rect 288636 8196 288637 8260
rect 288571 8195 288637 8196
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 298142 66877 298202 225523
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 299611 186964 299677 186965
rect 299611 186900 299612 186964
rect 299676 186900 299677 186964
rect 299611 186899 299677 186900
rect 298691 181524 298757 181525
rect 298691 181460 298692 181524
rect 298756 181460 298757 181524
rect 298691 181459 298757 181460
rect 298139 66876 298205 66877
rect 298139 66812 298140 66876
rect 298204 66812 298205 66876
rect 298139 66811 298205 66812
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 298694 4045 298754 181459
rect 299614 86325 299674 186899
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 302742 111077 302802 240755
rect 302739 111076 302805 111077
rect 302739 111012 302740 111076
rect 302804 111012 302805 111076
rect 302739 111011 302805 111012
rect 304214 89045 304274 302227
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 305499 187100 305565 187101
rect 305499 187036 305500 187100
rect 305564 187036 305565 187100
rect 305499 187035 305565 187036
rect 305502 135965 305562 187035
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 305499 135964 305565 135965
rect 305499 135900 305500 135964
rect 305564 135900 305565 135964
rect 305499 135899 305565 135900
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 304211 89044 304277 89045
rect 304211 88980 304212 89044
rect 304276 88980 304277 89044
rect 304211 88979 304277 88980
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 299611 86324 299677 86325
rect 299611 86260 299612 86324
rect 299676 86260 299677 86324
rect 299611 86259 299677 86260
rect 300954 86294 301574 86378
rect 299614 11797 299674 86259
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 299611 11796 299677 11797
rect 299611 11732 299612 11796
rect 299676 11732 299677 11796
rect 299611 11731 299677 11732
rect 298691 4044 298757 4045
rect 298691 3980 298692 4044
rect 298756 3980 298757 4044
rect 298691 3979 298757 3980
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 349174 312134 375600
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 352894 315854 375600
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 356614 319574 375600
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 363454 326414 375600
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 367174 330134 375600
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 370894 333854 375600
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 374614 337574 375600
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 345454 344414 375600
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 349174 348134 375600
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 352894 351854 375600
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 352054 310453 352114 544035
rect 352235 541244 352301 541245
rect 352235 541180 352236 541244
rect 352300 541180 352301 541244
rect 352235 541179 352301 541180
rect 352238 376549 352298 541179
rect 352235 376548 352301 376549
rect 352235 376484 352236 376548
rect 352300 376484 352301 376548
rect 352235 376483 352301 376484
rect 352051 310452 352117 310453
rect 352051 310388 352052 310452
rect 352116 310388 352117 310452
rect 352051 310387 352117 310388
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 353342 124133 353402 546619
rect 354954 537993 355574 572058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 356099 542468 356165 542469
rect 356099 542404 356100 542468
rect 356164 542404 356165 542468
rect 356099 542403 356165 542404
rect 356102 485790 356162 542403
rect 360147 514996 360213 514997
rect 360147 514932 360148 514996
rect 360212 514932 360213 514996
rect 360147 514931 360213 514932
rect 356283 499900 356349 499901
rect 356283 499836 356284 499900
rect 356348 499836 356349 499900
rect 356283 499835 356349 499836
rect 356286 499590 356346 499835
rect 356286 499530 356714 499590
rect 356102 485730 356530 485790
rect 356283 480180 356349 480181
rect 356283 480116 356284 480180
rect 356348 480116 356349 480180
rect 356283 480115 356349 480116
rect 356286 479770 356346 480115
rect 354814 479710 356346 479770
rect 354814 473370 354874 479710
rect 356470 476130 356530 485730
rect 354446 473310 354874 473370
rect 356102 476070 356530 476130
rect 354446 389190 354506 473310
rect 354446 389130 354690 389190
rect 354630 379530 354690 389130
rect 356102 382669 356162 476070
rect 356654 470610 356714 499530
rect 360150 485790 360210 514931
rect 359966 485730 360210 485790
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 359966 476130 360026 485730
rect 359966 476070 360210 476130
rect 356286 470550 356714 470610
rect 356286 386430 356346 470550
rect 357571 438972 357637 438973
rect 357571 438908 357572 438972
rect 357636 438908 357637 438972
rect 357571 438907 357637 438908
rect 356286 386370 356530 386430
rect 356470 383210 356530 386370
rect 356286 383150 356530 383210
rect 356099 382668 356165 382669
rect 356099 382604 356100 382668
rect 356164 382604 356165 382668
rect 356099 382603 356165 382604
rect 356099 381988 356165 381989
rect 356099 381924 356100 381988
rect 356164 381924 356165 381988
rect 356099 381923 356165 381924
rect 356102 381850 356162 381923
rect 354446 379470 354690 379530
rect 354814 381790 356162 381850
rect 354446 375730 354506 379470
rect 354627 375732 354693 375733
rect 354627 375730 354628 375732
rect 354446 375670 354628 375730
rect 354627 375668 354628 375670
rect 354692 375668 354693 375732
rect 354627 375667 354693 375668
rect 354814 347790 354874 381790
rect 354446 347730 354874 347790
rect 354954 356614 355574 375600
rect 356286 364989 356346 383150
rect 356467 382668 356533 382669
rect 356467 382604 356468 382668
rect 356532 382604 356533 382668
rect 356467 382603 356533 382604
rect 356470 374101 356530 382603
rect 356467 374100 356533 374101
rect 356467 374036 356468 374100
rect 356532 374036 356533 374100
rect 356467 374035 356533 374036
rect 357574 373285 357634 438907
rect 358859 409460 358925 409461
rect 358859 409396 358860 409460
rect 358924 409396 358925 409460
rect 358859 409395 358925 409396
rect 357571 373284 357637 373285
rect 357571 373220 357572 373284
rect 357636 373220 357637 373284
rect 357571 373219 357637 373220
rect 358862 371381 358922 409395
rect 360150 389190 360210 476070
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 360331 396948 360397 396949
rect 360331 396884 360332 396948
rect 360396 396884 360397 396948
rect 360331 396883 360397 396884
rect 359966 389130 360210 389190
rect 359966 379530 360026 389130
rect 359966 379470 360210 379530
rect 359411 378180 359477 378181
rect 359411 378116 359412 378180
rect 359476 378116 359477 378180
rect 359411 378115 359477 378116
rect 359414 376957 359474 378115
rect 359411 376956 359477 376957
rect 359411 376892 359412 376956
rect 359476 376892 359477 376956
rect 359411 376891 359477 376892
rect 358859 371380 358925 371381
rect 358859 371316 358860 371380
rect 358924 371316 358925 371380
rect 358859 371315 358925 371316
rect 356283 364988 356349 364989
rect 356283 364924 356284 364988
rect 356348 364924 356349 364988
rect 356283 364923 356349 364924
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354446 341597 354506 347730
rect 354443 341596 354509 341597
rect 354443 341532 354444 341596
rect 354508 341532 354509 341596
rect 354443 341531 354509 341532
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 353339 124132 353405 124133
rect 353339 124068 353340 124132
rect 353404 124068 353405 124132
rect 353339 124067 353405 124068
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 104614 355574 140058
rect 360150 125493 360210 379470
rect 360334 368389 360394 396883
rect 360331 368388 360397 368389
rect 360331 368324 360332 368388
rect 360396 368324 360397 368388
rect 360331 368323 360397 368324
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 360147 125492 360213 125493
rect 360147 125428 360148 125492
rect 360212 125428 360213 125492
rect 360147 125427 360213 125428
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 398603 185060 398669 185061
rect 398603 184996 398604 185060
rect 398668 184996 398669 185060
rect 398603 184995 398669 184996
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 142000 398414 146898
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 398606 136237 398666 184995
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 142000 402134 150618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 142000 405854 154338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 412403 229804 412469 229805
rect 412403 229740 412404 229804
rect 412468 229740 412469 229804
rect 412403 229739 412469 229740
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 142000 409574 158058
rect 412406 137730 412466 229739
rect 414243 227084 414309 227085
rect 414243 227020 414244 227084
rect 414308 227020 414309 227084
rect 414243 227019 414309 227020
rect 412406 137670 412834 137730
rect 398603 136236 398669 136237
rect 398603 136172 398604 136236
rect 398668 136172 398669 136236
rect 398603 136171 398669 136172
rect 402544 129454 402864 129486
rect 402544 129218 402586 129454
rect 402822 129218 402864 129454
rect 402544 129134 402864 129218
rect 402544 128898 402586 129134
rect 402822 128898 402864 129134
rect 402544 128866 402864 128898
rect 405744 129454 406064 129486
rect 405744 129218 405786 129454
rect 406022 129218 406064 129454
rect 405744 129134 406064 129218
rect 405744 128898 405786 129134
rect 406022 128898 406064 129134
rect 405744 128866 406064 128898
rect 408944 129454 409264 129486
rect 408944 129218 408986 129454
rect 409222 129218 409264 129454
rect 408944 129134 409264 129218
rect 408944 128898 408986 129134
rect 409222 128898 409264 129134
rect 408944 128866 409264 128898
rect 412144 129454 412464 129486
rect 412144 129218 412186 129454
rect 412422 129218 412464 129454
rect 412144 129134 412464 129218
rect 412144 128898 412186 129134
rect 412422 128898 412464 129134
rect 412144 128866 412464 128898
rect 404144 111454 404464 111486
rect 404144 111218 404186 111454
rect 404422 111218 404464 111454
rect 404144 111134 404464 111218
rect 404144 110898 404186 111134
rect 404422 110898 404464 111134
rect 404144 110866 404464 110898
rect 407344 111454 407664 111486
rect 407344 111218 407386 111454
rect 407622 111218 407664 111454
rect 407344 111134 407664 111218
rect 407344 110898 407386 111134
rect 407622 110898 407664 111134
rect 407344 110866 407664 110898
rect 410544 111454 410864 111486
rect 410544 111218 410586 111454
rect 410822 111218 410864 111454
rect 410544 111134 410864 111218
rect 410544 110898 410586 111134
rect 410822 110898 410864 111134
rect 410544 110866 410864 110898
rect 397499 108356 397565 108357
rect 397499 108292 397500 108356
rect 397564 108292 397565 108356
rect 397499 108291 397565 108292
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 397502 102781 397562 108291
rect 399891 103188 399957 103189
rect 399891 103124 399892 103188
rect 399956 103124 399957 103188
rect 399891 103123 399957 103124
rect 399894 103050 399954 103123
rect 399894 102990 400322 103050
rect 397499 102780 397565 102781
rect 397499 102716 397500 102780
rect 397564 102716 397565 102780
rect 397499 102715 397565 102716
rect 400262 99245 400322 102990
rect 412774 101690 412834 137670
rect 413744 111454 414064 111486
rect 413744 111218 413786 111454
rect 414022 111218 414064 111454
rect 413744 111134 414064 111218
rect 413744 110898 413786 111134
rect 414022 110898 414064 111134
rect 413744 110866 414064 110898
rect 412406 101630 412834 101690
rect 412406 99925 412466 101630
rect 414246 99925 414306 227019
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 142000 416414 164898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 142000 420134 168618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 142000 423854 172338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433379 210356 433445 210357
rect 433379 210292 433380 210356
rect 433444 210292 433445 210356
rect 433379 210291 433445 210292
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 424179 142220 424245 142221
rect 424179 142156 424180 142220
rect 424244 142156 424245 142220
rect 424179 142155 424245 142156
rect 420867 139500 420933 139501
rect 420867 139436 420868 139500
rect 420932 139436 420933 139500
rect 420867 139435 420933 139436
rect 415344 129454 415664 129486
rect 415344 129218 415386 129454
rect 415622 129218 415664 129454
rect 415344 129134 415664 129218
rect 415344 128898 415386 129134
rect 415622 128898 415664 129134
rect 415344 128866 415664 128898
rect 418544 129454 418864 129486
rect 418544 129218 418586 129454
rect 418822 129218 418864 129454
rect 418544 129134 418864 129218
rect 418544 128898 418586 129134
rect 418822 128898 418864 129134
rect 418544 128866 418864 128898
rect 416944 111454 417264 111486
rect 416944 111218 416986 111454
rect 417222 111218 417264 111454
rect 416944 111134 417264 111218
rect 416944 110898 416986 111134
rect 417222 110898 417264 111134
rect 416944 110866 417264 110898
rect 420144 111454 420464 111486
rect 420144 111218 420186 111454
rect 420422 111218 420464 111454
rect 420144 111134 420464 111218
rect 420144 110898 420186 111134
rect 420422 110898 420464 111134
rect 420144 110866 420464 110898
rect 412403 99924 412469 99925
rect 412403 99860 412404 99924
rect 412468 99860 412469 99924
rect 412403 99859 412469 99860
rect 414243 99924 414309 99925
rect 414243 99860 414244 99924
rect 414308 99860 414309 99924
rect 414243 99859 414309 99860
rect 400259 99244 400325 99245
rect 400259 99180 400260 99244
rect 400324 99180 400325 99244
rect 400259 99179 400325 99180
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 75454 398414 98000
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 79174 402134 98000
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 82894 405854 98000
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 86614 409574 98000
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 93454 416414 98000
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 97174 420134 98000
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 420870 7581 420930 139435
rect 421744 129454 422064 129486
rect 421744 129218 421786 129454
rect 422022 129218 422064 129454
rect 421744 129134 422064 129218
rect 421744 128898 421786 129134
rect 422022 128898 422064 129134
rect 421744 128866 422064 128898
rect 423344 111454 423664 111486
rect 423344 111218 423386 111454
rect 423622 111218 423664 111454
rect 423344 111134 423664 111218
rect 423344 110898 423386 111134
rect 423622 110898 423664 111134
rect 423344 110866 423664 110898
rect 423234 64894 423854 98000
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 424182 60621 424242 142155
rect 426954 142000 427574 176058
rect 425467 139500 425533 139501
rect 425467 139436 425468 139500
rect 425532 139436 425533 139500
rect 425467 139435 425533 139436
rect 426387 139500 426453 139501
rect 426387 139436 426388 139500
rect 426452 139436 426453 139500
rect 426387 139435 426453 139436
rect 430619 139500 430685 139501
rect 430619 139436 430620 139500
rect 430684 139436 430685 139500
rect 430619 139435 430685 139436
rect 424944 129454 425264 129486
rect 424944 129218 424986 129454
rect 425222 129218 425264 129454
rect 424944 129134 425264 129218
rect 424944 128898 424986 129134
rect 425222 128898 425264 129134
rect 424944 128866 425264 128898
rect 424179 60620 424245 60621
rect 424179 60556 424180 60620
rect 424244 60556 424245 60620
rect 424179 60555 424245 60556
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 420867 7580 420933 7581
rect 420867 7516 420868 7580
rect 420932 7516 420933 7580
rect 420867 7515 420933 7516
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 -5146 423854 28338
rect 425470 14517 425530 139435
rect 426390 77893 426450 139435
rect 428144 129454 428464 129486
rect 428144 129218 428186 129454
rect 428422 129218 428464 129454
rect 428144 129134 428464 129218
rect 428144 128898 428186 129134
rect 428422 128898 428464 129134
rect 428144 128866 428464 128898
rect 426544 111454 426864 111486
rect 426544 111218 426586 111454
rect 426822 111218 426864 111454
rect 426544 111134 426864 111218
rect 426544 110898 426586 111134
rect 426822 110898 426864 111134
rect 426544 110866 426864 110898
rect 429744 111454 430064 111486
rect 429744 111218 429786 111454
rect 430022 111218 430064 111454
rect 429744 111134 430064 111218
rect 429744 110898 429786 111134
rect 430022 110898 430064 111134
rect 429744 110866 430064 110898
rect 426387 77892 426453 77893
rect 426387 77828 426388 77892
rect 426452 77828 426453 77892
rect 426387 77827 426453 77828
rect 426954 68614 427574 98000
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 430622 68237 430682 139435
rect 431344 129454 431664 129486
rect 431344 129218 431386 129454
rect 431622 129218 431664 129454
rect 431344 129134 431664 129218
rect 431344 128898 431386 129134
rect 431622 128898 431664 129134
rect 431344 128866 431664 128898
rect 432944 111454 433264 111486
rect 432944 111218 432986 111454
rect 433222 111218 433264 111454
rect 432944 111134 433264 111218
rect 432944 110898 432986 111134
rect 433222 110898 433264 111134
rect 432944 110866 433264 110898
rect 433382 99925 433442 210291
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 435035 159356 435101 159357
rect 435035 159292 435036 159356
rect 435100 159292 435101 159356
rect 435035 159291 435101 159292
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 142000 434414 146898
rect 434544 129454 434864 129486
rect 434544 129218 434586 129454
rect 434822 129218 434864 129454
rect 434544 129134 434864 129218
rect 434544 128898 434586 129134
rect 434822 128898 434864 129134
rect 434544 128866 434864 128898
rect 435038 99925 435098 159291
rect 437514 151174 438134 186618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 438899 166292 438965 166293
rect 438899 166228 438900 166292
rect 438964 166228 438965 166292
rect 438899 166227 438965 166228
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 142000 438134 150618
rect 436691 139500 436757 139501
rect 436691 139436 436692 139500
rect 436756 139436 436757 139500
rect 436691 139435 436757 139436
rect 436144 111454 436464 111486
rect 436144 111218 436186 111454
rect 436422 111218 436464 111454
rect 436144 111134 436464 111218
rect 436144 110898 436186 111134
rect 436422 110898 436464 111134
rect 436144 110866 436464 110898
rect 433379 99924 433445 99925
rect 433379 99860 433380 99924
rect 433444 99860 433445 99924
rect 433379 99859 433445 99860
rect 435035 99924 435101 99925
rect 435035 99860 435036 99924
rect 435100 99860 435101 99924
rect 435035 99859 435101 99860
rect 433794 75454 434414 98000
rect 434851 97884 434917 97885
rect 434851 97820 434852 97884
rect 434916 97820 434917 97884
rect 434851 97819 434917 97820
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 430619 68236 430685 68237
rect 430619 68172 430620 68236
rect 430684 68172 430685 68236
rect 430619 68171 430685 68172
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 425467 14516 425533 14517
rect 425467 14452 425468 14516
rect 425532 14452 425533 14516
rect 425467 14451 425533 14452
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 434854 30973 434914 97819
rect 436694 55861 436754 139435
rect 437744 129454 438064 129486
rect 437744 129218 437786 129454
rect 438022 129218 438064 129454
rect 437744 129134 438064 129218
rect 437744 128898 437786 129134
rect 438022 128898 438064 129134
rect 437744 128866 438064 128898
rect 438902 125490 438962 166227
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 142000 441854 154338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 440187 140860 440253 140861
rect 440187 140796 440188 140860
rect 440252 140796 440253 140860
rect 440187 140795 440253 140796
rect 439083 139364 439149 139365
rect 439083 139300 439084 139364
rect 439148 139300 439149 139364
rect 439083 139299 439149 139300
rect 439086 125610 439146 139299
rect 439086 125550 439514 125610
rect 438902 125430 439330 125490
rect 439270 120869 439330 125430
rect 439267 120868 439333 120869
rect 439267 120804 439268 120868
rect 439332 120804 439333 120868
rect 439267 120803 439333 120804
rect 439454 118690 439514 125550
rect 440190 121277 440250 140795
rect 441659 140044 441725 140045
rect 441659 139980 441660 140044
rect 441724 139980 441725 140044
rect 441659 139979 441725 139980
rect 440187 121276 440253 121277
rect 440187 121212 440188 121276
rect 440252 121212 440253 121276
rect 440187 121211 440253 121212
rect 441662 119373 441722 139979
rect 442027 138956 442093 138957
rect 442027 138892 442028 138956
rect 442092 138892 442093 138956
rect 442027 138891 442093 138892
rect 441659 119372 441725 119373
rect 441659 119308 441660 119372
rect 441724 119308 441725 119372
rect 441659 119307 441725 119308
rect 438902 118630 439514 118690
rect 438902 115950 438962 118630
rect 439267 115972 439333 115973
rect 438902 115890 439146 115950
rect 439267 115908 439268 115972
rect 439332 115908 439333 115972
rect 439267 115907 439333 115908
rect 437514 79174 438134 98000
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 436691 55860 436757 55861
rect 436691 55796 436692 55860
rect 436756 55796 436757 55860
rect 436691 55795 436757 55796
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 434851 30972 434917 30973
rect 434851 30908 434852 30972
rect 434916 30908 434917 30972
rect 434851 30907 434917 30908
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 7174 438134 42618
rect 439086 34509 439146 115890
rect 439270 111349 439330 115907
rect 439267 111348 439333 111349
rect 439267 111284 439268 111348
rect 439332 111284 439333 111348
rect 439267 111283 439333 111284
rect 441234 82894 441854 98000
rect 442030 90405 442090 138891
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 442027 90404 442093 90405
rect 442027 90340 442028 90404
rect 442092 90340 442093 90404
rect 442027 90339 442093 90340
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 439083 34508 439149 34509
rect 439083 34444 439084 34508
rect 439148 34444 439149 34508
rect 439083 34443 439149 34444
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 72721 579218 72957 579454
rect 72721 578898 72957 579134
rect 78651 579218 78887 579454
rect 78651 578898 78887 579134
rect 84582 579218 84818 579454
rect 84582 578898 84818 579134
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 75686 561218 75922 561454
rect 75686 560898 75922 561134
rect 81617 561218 81853 561454
rect 81617 560898 81853 561134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 72721 543218 72957 543454
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 72721 542898 72957 543134
rect 78651 543218 78887 543454
rect 78651 542898 78887 543134
rect 84582 543218 84818 543454
rect 84582 542898 84818 543134
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 73020 435218 73256 435454
rect 73020 434898 73256 435134
rect 88380 417218 88616 417454
rect 88380 416898 88616 417134
rect 73020 399218 73256 399454
rect 73020 398898 73256 399134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73020 291218 73256 291454
rect 73020 290898 73256 291134
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73020 255218 73256 255454
rect 73020 254898 73256 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 103740 435218 103976 435454
rect 103740 434898 103976 435134
rect 103740 399218 103976 399454
rect 103740 398898 103976 399134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 119100 417218 119336 417454
rect 119100 416898 119336 417134
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 88380 309218 88616 309454
rect 88380 308898 88616 309134
rect 119100 309218 119336 309454
rect 119100 308898 119336 309134
rect 149820 309218 150056 309454
rect 149820 308898 150056 309134
rect 103740 291218 103976 291454
rect 103740 290898 103976 291134
rect 134460 291218 134696 291454
rect 134460 290898 134696 291134
rect 88380 273218 88616 273454
rect 88380 272898 88616 273134
rect 119100 273218 119336 273454
rect 119100 272898 119336 273134
rect 149820 273218 150056 273454
rect 149820 272898 150056 273134
rect 103740 255218 103976 255454
rect 103740 254898 103976 255134
rect 134460 255218 134696 255454
rect 134460 254898 134696 255134
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 69128 165218 69364 165454
rect 69128 164898 69364 165134
rect 164192 165218 164428 165454
rect 164192 164898 164428 165134
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 69128 129218 69364 129454
rect 69128 128898 69364 129134
rect 164192 129218 164428 129454
rect 164192 128898 164428 129134
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 219610 525218 219846 525454
rect 219610 524898 219846 525134
rect 250330 525218 250566 525454
rect 250330 524898 250566 525134
rect 281050 525218 281286 525454
rect 281050 524898 281286 525134
rect 311770 525218 312006 525454
rect 311770 524898 312006 525134
rect 342490 525218 342726 525454
rect 342490 524898 342726 525134
rect 204250 507218 204486 507454
rect 204250 506898 204486 507134
rect 234970 507218 235206 507454
rect 234970 506898 235206 507134
rect 265690 507218 265926 507454
rect 265690 506898 265926 507134
rect 296410 507218 296646 507454
rect 296410 506898 296646 507134
rect 327130 507218 327366 507454
rect 327130 506898 327366 507134
rect 219610 489218 219846 489454
rect 219610 488898 219846 489134
rect 250330 489218 250566 489454
rect 250330 488898 250566 489134
rect 281050 489218 281286 489454
rect 281050 488898 281286 489134
rect 311770 489218 312006 489454
rect 311770 488898 312006 489134
rect 342490 489218 342726 489454
rect 342490 488898 342726 489134
rect 204250 471218 204486 471454
rect 204250 470898 204486 471134
rect 234970 471218 235206 471454
rect 234970 470898 235206 471134
rect 265690 471218 265926 471454
rect 265690 470898 265926 471134
rect 296410 471218 296646 471454
rect 296410 470898 296646 471134
rect 327130 471218 327366 471454
rect 327130 470898 327366 471134
rect 219610 453218 219846 453454
rect 219610 452898 219846 453134
rect 250330 453218 250566 453454
rect 250330 452898 250566 453134
rect 281050 453218 281286 453454
rect 281050 452898 281286 453134
rect 311770 453218 312006 453454
rect 311770 452898 312006 453134
rect 342490 453218 342726 453454
rect 342490 452898 342726 453134
rect 204250 435218 204486 435454
rect 204250 434898 204486 435134
rect 234970 435218 235206 435454
rect 234970 434898 235206 435134
rect 265690 435218 265926 435454
rect 265690 434898 265926 435134
rect 296410 435218 296646 435454
rect 296410 434898 296646 435134
rect 327130 435218 327366 435454
rect 327130 434898 327366 435134
rect 219610 417218 219846 417454
rect 219610 416898 219846 417134
rect 250330 417218 250566 417454
rect 250330 416898 250566 417134
rect 281050 417218 281286 417454
rect 281050 416898 281286 417134
rect 311770 417218 312006 417454
rect 311770 416898 312006 417134
rect 342490 417218 342726 417454
rect 342490 416898 342726 417134
rect 204250 399218 204486 399454
rect 204250 398898 204486 399134
rect 234970 399218 235206 399454
rect 234970 398898 235206 399134
rect 265690 399218 265926 399454
rect 265690 398898 265926 399134
rect 296410 399218 296646 399454
rect 296410 398898 296646 399134
rect 327130 399218 327366 399454
rect 327130 398898 327366 399134
rect 219610 381218 219846 381454
rect 219610 380898 219846 381134
rect 250330 381218 250566 381454
rect 250330 380898 250566 381134
rect 281050 381218 281286 381454
rect 281050 380898 281286 381134
rect 311770 381218 312006 381454
rect 311770 380898 312006 381134
rect 342490 381218 342726 381454
rect 342490 380898 342726 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 204450 255218 204686 255454
rect 204450 254898 204686 255134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 219810 273218 220046 273454
rect 219810 272898 220046 273134
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 221249 165218 221485 165454
rect 221249 164898 221485 165134
rect 224513 165218 224749 165454
rect 224513 164898 224749 165134
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 219617 147218 219853 147454
rect 219617 146898 219853 147134
rect 222881 147218 223117 147454
rect 222881 146898 223117 147134
rect 226145 147218 226381 147454
rect 226145 146898 226381 147134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 235170 255218 235406 255454
rect 235170 254898 235406 255134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 221249 129218 221485 129454
rect 221249 128898 221485 129134
rect 224513 129218 224749 129454
rect 224513 128898 224749 129134
rect 219617 111218 219853 111454
rect 219617 110898 219853 111134
rect 222881 111218 223117 111454
rect 222881 110898 223117 111134
rect 226145 111218 226381 111454
rect 226145 110898 226381 111134
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 272249 165218 272485 165454
rect 272249 164898 272485 165134
rect 275513 165218 275749 165454
rect 275513 164898 275749 165134
rect 270617 147218 270853 147454
rect 270617 146898 270853 147134
rect 273881 147218 274117 147454
rect 273881 146898 274117 147134
rect 277145 147218 277381 147454
rect 277145 146898 277381 147134
rect 272249 129218 272485 129454
rect 272249 128898 272485 129134
rect 275513 129218 275749 129454
rect 275513 128898 275749 129134
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 270617 111218 270853 111454
rect 270617 110898 270853 111134
rect 273881 111218 274117 111454
rect 273881 110898 274117 111134
rect 277145 111218 277381 111454
rect 277145 110898 277381 111134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 402586 129218 402822 129454
rect 402586 128898 402822 129134
rect 405786 129218 406022 129454
rect 405786 128898 406022 129134
rect 408986 129218 409222 129454
rect 408986 128898 409222 129134
rect 412186 129218 412422 129454
rect 412186 128898 412422 129134
rect 404186 111218 404422 111454
rect 404186 110898 404422 111134
rect 407386 111218 407622 111454
rect 407386 110898 407622 111134
rect 410586 111218 410822 111454
rect 410586 110898 410822 111134
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 413786 111218 414022 111454
rect 413786 110898 414022 111134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 415386 129218 415622 129454
rect 415386 128898 415622 129134
rect 418586 129218 418822 129454
rect 418586 128898 418822 129134
rect 416986 111218 417222 111454
rect 416986 110898 417222 111134
rect 420186 111218 420422 111454
rect 420186 110898 420422 111134
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 421786 129218 422022 129454
rect 421786 128898 422022 129134
rect 423386 111218 423622 111454
rect 423386 110898 423622 111134
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 424986 129218 425222 129454
rect 424986 128898 425222 129134
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 428186 129218 428422 129454
rect 428186 128898 428422 129134
rect 426586 111218 426822 111454
rect 426586 110898 426822 111134
rect 429786 111218 430022 111454
rect 429786 110898 430022 111134
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 431386 129218 431622 129454
rect 431386 128898 431622 129134
rect 432986 111218 433222 111454
rect 432986 110898 433222 111134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 434586 129218 434822 129454
rect 434586 128898 434822 129134
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 436186 111218 436422 111454
rect 436186 110898 436422 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 437786 129218 438022 129454
rect 437786 128898 438022 129134
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 72721 579454
rect 72957 579218 78651 579454
rect 78887 579218 84582 579454
rect 84818 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 72721 579134
rect 72957 578898 78651 579134
rect 78887 578898 84582 579134
rect 84818 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 75686 561454
rect 75922 561218 81617 561454
rect 81853 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 75686 561134
rect 75922 560898 81617 561134
rect 81853 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 72721 543454
rect 72957 543218 78651 543454
rect 78887 543218 84582 543454
rect 84818 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 72721 543134
rect 72957 542898 78651 543134
rect 78887 542898 84582 543134
rect 84818 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 219610 525454
rect 219846 525218 250330 525454
rect 250566 525218 281050 525454
rect 281286 525218 311770 525454
rect 312006 525218 342490 525454
rect 342726 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 219610 525134
rect 219846 524898 250330 525134
rect 250566 524898 281050 525134
rect 281286 524898 311770 525134
rect 312006 524898 342490 525134
rect 342726 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 204250 507454
rect 204486 507218 234970 507454
rect 235206 507218 265690 507454
rect 265926 507218 296410 507454
rect 296646 507218 327130 507454
rect 327366 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 204250 507134
rect 204486 506898 234970 507134
rect 235206 506898 265690 507134
rect 265926 506898 296410 507134
rect 296646 506898 327130 507134
rect 327366 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 219610 489454
rect 219846 489218 250330 489454
rect 250566 489218 281050 489454
rect 281286 489218 311770 489454
rect 312006 489218 342490 489454
rect 342726 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 219610 489134
rect 219846 488898 250330 489134
rect 250566 488898 281050 489134
rect 281286 488898 311770 489134
rect 312006 488898 342490 489134
rect 342726 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 204250 471454
rect 204486 471218 234970 471454
rect 235206 471218 265690 471454
rect 265926 471218 296410 471454
rect 296646 471218 327130 471454
rect 327366 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 204250 471134
rect 204486 470898 234970 471134
rect 235206 470898 265690 471134
rect 265926 470898 296410 471134
rect 296646 470898 327130 471134
rect 327366 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 219610 453454
rect 219846 453218 250330 453454
rect 250566 453218 281050 453454
rect 281286 453218 311770 453454
rect 312006 453218 342490 453454
rect 342726 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 219610 453134
rect 219846 452898 250330 453134
rect 250566 452898 281050 453134
rect 281286 452898 311770 453134
rect 312006 452898 342490 453134
rect 342726 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73020 435454
rect 73256 435218 103740 435454
rect 103976 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 204250 435454
rect 204486 435218 234970 435454
rect 235206 435218 265690 435454
rect 265926 435218 296410 435454
rect 296646 435218 327130 435454
rect 327366 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73020 435134
rect 73256 434898 103740 435134
rect 103976 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 204250 435134
rect 204486 434898 234970 435134
rect 235206 434898 265690 435134
rect 265926 434898 296410 435134
rect 296646 434898 327130 435134
rect 327366 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 88380 417454
rect 88616 417218 119100 417454
rect 119336 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 219610 417454
rect 219846 417218 250330 417454
rect 250566 417218 281050 417454
rect 281286 417218 311770 417454
rect 312006 417218 342490 417454
rect 342726 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 88380 417134
rect 88616 416898 119100 417134
rect 119336 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 219610 417134
rect 219846 416898 250330 417134
rect 250566 416898 281050 417134
rect 281286 416898 311770 417134
rect 312006 416898 342490 417134
rect 342726 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73020 399454
rect 73256 399218 103740 399454
rect 103976 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 204250 399454
rect 204486 399218 234970 399454
rect 235206 399218 265690 399454
rect 265926 399218 296410 399454
rect 296646 399218 327130 399454
rect 327366 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73020 399134
rect 73256 398898 103740 399134
rect 103976 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 204250 399134
rect 204486 398898 234970 399134
rect 235206 398898 265690 399134
rect 265926 398898 296410 399134
rect 296646 398898 327130 399134
rect 327366 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 219610 381454
rect 219846 381218 250330 381454
rect 250566 381218 281050 381454
rect 281286 381218 311770 381454
rect 312006 381218 342490 381454
rect 342726 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 219610 381134
rect 219846 380898 250330 381134
rect 250566 380898 281050 381134
rect 281286 380898 311770 381134
rect 312006 380898 342490 381134
rect 342726 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 88380 309454
rect 88616 309218 119100 309454
rect 119336 309218 149820 309454
rect 150056 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 88380 309134
rect 88616 308898 119100 309134
rect 119336 308898 149820 309134
rect 150056 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73020 291454
rect 73256 291218 103740 291454
rect 103976 291218 134460 291454
rect 134696 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73020 291134
rect 73256 290898 103740 291134
rect 103976 290898 134460 291134
rect 134696 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 88380 273454
rect 88616 273218 119100 273454
rect 119336 273218 149820 273454
rect 150056 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 219810 273454
rect 220046 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 88380 273134
rect 88616 272898 119100 273134
rect 119336 272898 149820 273134
rect 150056 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 219810 273134
rect 220046 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73020 255454
rect 73256 255218 103740 255454
rect 103976 255218 134460 255454
rect 134696 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 204450 255454
rect 204686 255218 235170 255454
rect 235406 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73020 255134
rect 73256 254898 103740 255134
rect 103976 254898 134460 255134
rect 134696 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 204450 255134
rect 204686 254898 235170 255134
rect 235406 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 69128 165454
rect 69364 165218 164192 165454
rect 164428 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 221249 165454
rect 221485 165218 224513 165454
rect 224749 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 272249 165454
rect 272485 165218 275513 165454
rect 275749 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 69128 165134
rect 69364 164898 164192 165134
rect 164428 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 221249 165134
rect 221485 164898 224513 165134
rect 224749 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 272249 165134
rect 272485 164898 275513 165134
rect 275749 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 219617 147454
rect 219853 147218 222881 147454
rect 223117 147218 226145 147454
rect 226381 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 270617 147454
rect 270853 147218 273881 147454
rect 274117 147218 277145 147454
rect 277381 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 219617 147134
rect 219853 146898 222881 147134
rect 223117 146898 226145 147134
rect 226381 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 270617 147134
rect 270853 146898 273881 147134
rect 274117 146898 277145 147134
rect 277381 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 69128 129454
rect 69364 129218 164192 129454
rect 164428 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 221249 129454
rect 221485 129218 224513 129454
rect 224749 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 272249 129454
rect 272485 129218 275513 129454
rect 275749 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 402586 129454
rect 402822 129218 405786 129454
rect 406022 129218 408986 129454
rect 409222 129218 412186 129454
rect 412422 129218 415386 129454
rect 415622 129218 418586 129454
rect 418822 129218 421786 129454
rect 422022 129218 424986 129454
rect 425222 129218 428186 129454
rect 428422 129218 431386 129454
rect 431622 129218 434586 129454
rect 434822 129218 437786 129454
rect 438022 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 69128 129134
rect 69364 128898 164192 129134
rect 164428 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 221249 129134
rect 221485 128898 224513 129134
rect 224749 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 272249 129134
rect 272485 128898 275513 129134
rect 275749 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 402586 129134
rect 402822 128898 405786 129134
rect 406022 128898 408986 129134
rect 409222 128898 412186 129134
rect 412422 128898 415386 129134
rect 415622 128898 418586 129134
rect 418822 128898 421786 129134
rect 422022 128898 424986 129134
rect 425222 128898 428186 129134
rect 428422 128898 431386 129134
rect 431622 128898 434586 129134
rect 434822 128898 437786 129134
rect 438022 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 219617 111454
rect 219853 111218 222881 111454
rect 223117 111218 226145 111454
rect 226381 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 270617 111454
rect 270853 111218 273881 111454
rect 274117 111218 277145 111454
rect 277381 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 404186 111454
rect 404422 111218 407386 111454
rect 407622 111218 410586 111454
rect 410822 111218 413786 111454
rect 414022 111218 416986 111454
rect 417222 111218 420186 111454
rect 420422 111218 423386 111454
rect 423622 111218 426586 111454
rect 426822 111218 429786 111454
rect 430022 111218 432986 111454
rect 433222 111218 436186 111454
rect 436422 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 219617 111134
rect 219853 110898 222881 111134
rect 223117 110898 226145 111134
rect 226381 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 270617 111134
rect 270853 110898 273881 111134
rect 274117 110898 277145 111134
rect 277381 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 404186 111134
rect 404422 110898 407386 111134
rect 407622 110898 410586 111134
rect 410822 110898 413786 111134
rect 414022 110898 416986 111134
rect 417222 110898 420186 111134
rect 420422 110898 423386 111134
rect 423622 110898 426586 111134
rect 426822 110898 429786 111134
rect 430022 110898 432986 111134
rect 433222 110898 436186 111134
rect 436422 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use wrapped_spell  wrapped_spell_1
timestamp 1640773853
transform 1 0 68770 0 1 241592
box 0 0 88000 88000
use wrapped_skullfet  wrapped_skullfet_5
timestamp 1640773853
transform 1 0 400000 0 1 100000
box -10 -52 40000 40000
use wrapped_silife  wrapped_silife_4
timestamp 1640773853
transform 1 0 200000 0 1 377600
box -10 0 156249 158393
use wrapped_ppm_decoder  wrapped_ppm_decoder_3
timestamp 1640773853
transform 1 0 68770 0 1 539166
box -10 0 20000 50000
use wrapped_ppm_coder  wrapped_ppm_coder_2
timestamp 1640773853
transform 1 0 68770 0 1 390356
box -10 0 51907 54051
use wrapped_function_generator  wrapped_function_generator_0
timestamp 1640773853
transform 1 0 200200 0 1 240182
box 0 0 44000 44000
use wb_openram_wrapper  wb_openram_wrapper
timestamp 1640773853
transform 1 0 217000 0 1 96000
box 0 144 12000 79688
use wb_bridge_2way  wb_bridge_2way
timestamp 1640773853
transform 1 0 268000 0 1 96000
box 0 0 12000 79688
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 1640773853
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 94000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 178000 218414 238182 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 176600 74414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 176600 110414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 176600 146414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 286182 218414 375600 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 375600 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 375600 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 375600 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 331592 74414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 331592 110414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 446407 74414 537166 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 591166 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 446407 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 331592 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 537993 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 537993 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 537993 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 537993 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 142000 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 142000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 94000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 178000 222134 238182 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 176600 78134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 176600 114134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 176600 150134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 286182 222134 375600 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 375600 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 375600 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 375600 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 331592 78134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 331592 114134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 446407 78134 537166 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 591166 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 446407 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 331592 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 537993 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 537993 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 537993 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 537993 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 142000 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 142000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 94000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 178000 225854 238182 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 176600 81854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 176600 117854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 176600 153854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 286182 225854 375600 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 375600 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 375600 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 375600 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 331592 81854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 331592 117854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 446407 81854 537166 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 591166 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 446407 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 331592 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 537993 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 537993 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 537993 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 537993 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 142000 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 142000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 94000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 178000 229574 238182 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 176600 85574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 176600 121574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 176600 157574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 286182 229574 375600 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 375600 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 375600 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 375600 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 331592 85574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 331592 121574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 446407 85574 537166 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 591166 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 446407 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 331592 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 537993 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 537993 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 537993 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 537993 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 142000 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 238182 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 238182 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 176600 99854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 176600 135854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 286182 207854 375600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 286182 243854 375600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 178000 279854 375600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 375600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 375600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 331592 99854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 446407 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 331592 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 537993 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 537993 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 537993 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 537993 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 537993 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 142000 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 238182 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 176600 67574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 176600 103574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 176600 139574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 286182 211574 375600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 375600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 375600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 375600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 375600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 331592 67574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 331592 103574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 446407 67574 537166 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 591166 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 446407 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 331592 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 537993 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 537993 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 537993 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 537993 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 537993 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 142000 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 238182 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 238182 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 176600 92414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 176600 128414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 286182 200414 375600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 286182 236414 375600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 178000 272414 375600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 375600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 375600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 331592 92414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 446407 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 331592 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 176600 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 537993 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 537993 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 537993 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 537993 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 537993 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 142000 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 238182 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 238182 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 176600 96134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 176600 132134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 286182 204134 375600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 286182 240134 375600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 178000 276134 375600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 375600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 375600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 331592 96134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 446407 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 331592 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 537993 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 537993 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 537993 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 537993 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 537993 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 142000 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
